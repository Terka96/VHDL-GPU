library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.definitions.all;

package texture is

constant TEX_SIZE_F : FLOAT16 := x"5400";
constant TEX_SIZE	: integer := 64;
type TEXTURE_MEM_LINE is array (0 to (TEX_SIZE-1)) of COLOR24;
type TEXTURE_MEM is array (0 to (TEX_SIZE-1)) of TEXTURE_MEM_LINE;

  constant texture_memory_const : TEXTURE_MEM := ( 
(x"5c5656",x"6f6764",x"504c4d",x"524e4d",x"5c5250",x"544e4e",x"5c5354",x"656160",x"584f50",x"615652",x"665c5a",x"69615e",x"8e817b",x"877c78",x"7f726c",x"81746c",x"7f7573",x"807674",x"8e8381",x"796c64",x"8c817b",x"948985",x"89807b",x"968c8b",x"8b807c",x"494544",x"8f8681",x"94857e",x"6f6b6a",x"7b7673",x"817670",x"746c69",x"5b5555",x"656364",x"696768",x"656366",x"62615f",x"5f5f5f",x"6b6a68",x"696768",x"66656a",x"5f5e63",x"626264",x"796e68",x"948a80",x"988b83",x"9a8d85",x"998a83",x"9e9590",x"998b82",x"9b8e86",x"988e85",x"968b85",x"988984",x"9c8e85",x"988e8c",x"907f77",x"9a8f89",x"928982",x"998c84",x"5c5250",x"615755",x"535250",x"57524f"),
(x"89807b",x"877e79",x"877c78",x"827771",x"827974",x"887b73",x"837872",x"7f726a",x"80736b",x"7e7169",x"8b7d7a",x"877a72",x"5f5a57",x"615957",x"565253",x"595051",x"625a57",x"655a58",x"544e4e",x"574f4d",x"655c57",x"545454",x"625c5c",x"625e5b",x"635f5e",x"6e6159",x"6a564f",x"595556",x"958b89",x"9e938d",x"9a8f89",x"9e948b",x"9c8e85",x"94877f",x"988b85",x"968d86",x"9c918b",x"998880",x"978e87",x"9a8f89",x"958882",x"92857f",x"a09591",x"9e948b",x"605c5d",x"68605d",x"625a58",x"675d5b",x"6c6260",x"645a58",x"5f5b5c",x"675d5b",x"655d5a",x"625a57",x"695e5c",x"605953",x"6f6661",x"594e4c",x"5f5959",x"695a53",x"928177",x"847a79",x"7e7472",x"837a75"),
(x"796c64",x"82736c",x"7b716f",x"837874",x"81776e",x"827771",x"7f7470",x"8a7972",x"907a6d",x"85746c",x"80736b",x"80736d",x"4a4647",x"5f5959",x"5b5253",x"554c47",x"5d585c",x"5e5654",x"5c5451",x"5a5250",x"54504d",x"5c5857",x"5a5859",x"626061",x"5e5956",x"72655d",x"685d59",x"686360",x"9d9088",x"988e85",x"968b85",x"978a82",x"92857d",x"90817a",x"95867f",x"6f6158",x"817068",x"96887f",x"988b85",x"a39892",x"8f827c",x"998c84",x"9e938f",x"a2988f",x"63595a",x"5e5c5d",x"665c5a",x"675c56",x"72685f",x"5c5754",x"6b6565",x"615c59",x"615755",x"5d5553",x"746963",x"62554f",x"695c56",x"6e6463",x"5e5452",x"685952",x"8c7f79",x"746761",x"776861",x"7d6c65"),
(x"7f7069",x"776c66",x"716660",x"796a63",x"82736c",x"7e716b",x"806c61",x"807269",x"85766f",x"86786f",x"786a61",x"7e6f68",x"4f4745",x"5c5452",x"665d58",x"584e4d",x"5e5956",x"645c5a",x"5d5553",x"4e4946",x"625856",x"5d564e",x"555354",x"5b595a",x"5b5754",x"575354",x"6c5f57",x"66615d",x"99908b",x"9a9087",x"9f958c",x"9f928a",x"978a82",x"988d87",x"938882",x"9a8c83",x"897871",x"978a82",x"978a84",x"9d948d",x"9a918a",x"9c938e",x"998c84",x"9c9289",x"6d6563",x"595353",x"635958",x"6e6560",x"685e5c",x"5e5654",x"645e5e",x"5e5a5b",x"625d5a",x"554b4c",x"5a4f4d",x"645a59",x"554c4d",x"4b403c",x"675c5a",x"5e5556",x"867b75",x"756862",x"776a64",x"7a6b64"),
(x"807269",x"796b68",x"87766e",x"8d7b71",x"8a7f7b",x"90817a",x"837268",x"817672",x"8e817b",x"8b7e78",x"83756c",x"8f8178",x"645a58",x"5f595b",x"5d5553",x"534f4c",x"665e5c",x"595353",x"665b57",x"605a5a",x"6d6361",x"615654",x"5a5657",x"5b595a",x"5d5855",x"595451",x"73665d",x"6b6263",x"a49993",x"9d938a",x"988982",x"a19690",x"a19997",x"988d87",x"9b8e86",x"978c86",x"93847d",x"9a8d85",x"968780",x"98918b",x"9b928b",x"978d84",x"8f8079",x"9d908a",x"726866",x"635b59",x"756c65",x"544f4c",x"4f4b4a",x"635e5b",x"5b5351",x"565050",x"5e5654",x"655b5a",x"5b5351",x"645655",x"52494a",x"62595a",x"645b5c",x"554d4b",x"7d726e",x"847771",x"726761",x"7d6e67"),
(x"776f6d",x"877c76",x"8b807a",x"837874",x"928785",x"907f75",x"857a74",x"7c7269",x"8e857e",x"8f827a",x"8f827c",x"8d7e77",x"6a6260",x"655c57",x"635a55",x"615654",x"605655",x"424242",x"5a5152",x"5f5754",x"534f50",x"574d4c",x"564e4b",x"4f4e4c",x"615650",x"4a4645",x"756663",x"7d6b5d",x"a39892",x"a49b94",x"94857e",x"9f9892",x"998a83",x"988a81",x"91847c",x"988f8a",x"948b84",x"574c46",x"948985",x"968983",x"968983",x"948983",x"97867f",x"988b83",x"5e5858",x"615755",x"605655",x"615b5b",x"635a5b",x"655d5b",x"625c5c",x"675d5c",x"655b5a",x"534d4f",x"5e5452",x"554f4f",x"5f5554",x"635854",x"615d5e",x"5c5859",x"817674",x"80716a",x"7c6b63",x"82736c"),
(x"766b67",x"655b5a",x"7d6f6c",x"918785",x"948b86",x"948781",x"8a817c",x"988780",x"8f817e",x"8f827c",x"897a75",x"8c7e75",x"6e605d",x"71645e",x"63595a",x"5c5452",x"4a4542",x"363231",x"3e3936",x"565251",x"686560",x"5c5656",x"635854",x"605654",x"5c5451",x"645d55",x"6f6460",x"6a5f5b",x"9f958c",x"a1978e",x"9d928c",x"9b9289",x"a49d97",x"9b928b",x"9e958e",x"988b83",x"9b948e",x"9e938d",x"9f928a",x"91827b",x"958882",x"897a73",x"90837b",x"91847e",x"6c6764",x"6b6361",x"5f5755",x"5b5555",x"736967",x"655b59",x"675c58",x"62595a",x"605655",x"645c5a",x"5e5654",x"615859",x"605a5a",x"5d595a",x"615d5e",x"5f5959",x"847975",x"857369",x"74655e",x"7f7069"),
(x"887d79",x"83766e",x"83756c",x"8b807c",x"8d827e",x"928783",x"94877f",x"938582",x"91847e",x"938882",x"857870",x"938b88",x"6a625f",x"6e6462",x"605655",x"5e5351",x"3e3936",x"393430",x"38302e",x"504c4d",x"514745",x"615956",x"565457",x"5b5350",x"595451",x"726761",x"5b5555",x"676161",x"a19891",x"958c85",x"978c86",x"a39690",x"8e847b",x"9a918a",x"9a8d87",x"998c84",x"a19690",x"948983",x"978e89",x"918682",x"8e817b",x"92837c",x"968981",x"90827f",x"675d5b",x"5f5755",x"6c6260",x"635958",x"5f5553",x"615756",x"6c6260",x"554d4b",x"625856",x"5e5452",x"605855",x"595353",x"6a605e",x"675c58",x"5c5859",x"5c5656",x"8b807c",x"81726b",x"81726b",x"786964"),
(x"7f746e",x"736967",x"7c716d",x"796e6c",x"918682",x"948985",x"958a86",x"938884",x"93867e",x"91847e",x"82756d",x"948983",x"695f5e",x"665e5c",x"5c5b59",x"605856",x"5a5152",x"6b6361",x"655b5a",x"484242",x"504a4a",x"5b5150",x"555354",x"5f5a56",x"685f58",x"504e4f",x"675e59",x"796a65",x"9a9188",x"9c8d86",x"9c938a",x"a0958f",x"9e948b",x"92857d",x"998c83",x"9a8d85",x"9a8b84",x"998b82",x"968981",x"9c8f87",x"948983",x"9c8a80",x"968480",x"948781",x"615755",x"675d5c",x"5f5657",x"605551",x"7d7573",x"84776f",x"615853",x"675d5c",x"665c5b",x"68635f",x"605654",x"685e5d",x"514f50",x"585252",x"615b5b",x"786d6b",x"786662",x"82756f",x"86786f",x"7a6f69"),
(x"897e7c",x"857872",x"867b77",x"90857f",x"918680",x"998e88",x"9b8e86",x"988b83",x"817068",x"887b73",x"9a8f8b",x"908279",x"646061",x"625c5c",x"5c5656",x"5c5857",x"695f5d",x"645a58",x"625857",x"5a5152",x"575256",x"554c4d",x"534e4b",x"4f4d4e",x"525053",x"665951",x"585453",x"5e5e60",x"9c938e",x"9a918a",x"978a84",x"9d928c",x"958a86",x"999089",x"989390",x"998c84",x"9a9087",x"94877f",x"998b82",x"90817a",x"968981",x"9b8e88",x"94857e",x"98918b",x"625d5a",x"685e5d",x"5d5553",x"5e5556",x"695f56",x"6a6057",x"6d625c",x"574f4d",x"5c5656",x"504846",x"5c5354",x"5e5a59",x"635a5b",x"695e5a",x"695a53",x"5b5758",x"918682",x"8e8179",x"91827b",x"857a76"),
(x"938882",x"8a7d74",x"847771",x"948983",x"978883",x"988f88",x"9b908c",x"897e7a",x"8a7b74",x"92857d",x"8a796f",x"9d908a",x"675e5f",x"675d5b",x"655c5d",x"5f5b5c",x"565253",x"645e5e",x"655b59",x"5e5858",x"615654",x"5f5755",x"5b5351",x"4c4849",x"4e4e50",x"58504e",x"655c57",x"61605e",x"9d9690",x"9e918b",x"988e85",x"9b908a",x"988d87",x"9e938d",x"9a8f89",x"9b8e85",x"9b8d84",x"998c84",x"8f8279",x"9d9087",x"968981",x"95877e",x"948983",x"998e8a",x"5a5250",x"5d5352",x"5d5457",x"695f5d",x"5e5452",x"605655",x"5c5754",x"665b59",x"615756",x"5a5250",x"584f50",x"5a5152",x"605a5a",x"625856",x"685e5d",x"635958",x"978a84",x"8a7f79",x"887b73",x"90817a"),
(x"8b807c",x"8d827e",x"92857d",x"968c8a",x"8f827c",x"9f9691",x"978c88",x"928982",x"8d7f76",x"988d87",x"786b62",x"887f78",x"646464",x"524e4f",x"534f50",x"4f4d4e",x"5f5554",x"5e5858",x"5b5150",x"605655",x"5e5654",x"504c4d",x"534e4b",x"5c534e",x"5e5654",x"534b49",x"635e5b",x"5a585d",x"8e8580",x"9f948e",x"93857c",x"a0968d",x"998f86",x"9c8f87",x"a0938b",x"9a8b84",x"9c938c",x"9a8a7d",x"9d8b81",x"998880",x"91827b",x"8e8179",x"968d88",x"907f77",x"625753",x"605856",x"4e4848",x"58504e",x"5e5453",x"655a58",x"625857",x"625a58",x"685e5d",x"655b5a",x"635957",x"655f5f",x"605a5c",x"5f5651",x"5e5452",x"564b47",x"897c74",x"978883",x"94867d",x"8b7d72"),
(x"83766e",x"8c7d76",x"9b908a",x"8e8482",x"998e8a",x"8b796d",x"92857f",x"988b83",x"95847a",x"8e837f",x"887a6f",x"8a7b74",x"6d625e",x"675d5c",x"635d5d",x"5d5553",x"4d4b4c",x"545253",x"5a524f",x"665e5c",x"605a5a",x"5c5754",x"5a504f",x"5a504f",x"605856",x"5d5553",x"59514e",x"5f5755",x"9f958c",x"978a82",x"8b807a",x"a69d96",x"9e948b",x"9c8f87",x"998c84",x"9b8e85",x"9b8d84",x"9f9289",x"9b8e86",x"968980",x"9b8e85",x"968780",x"998e8a",x"7e7473",x"615b5b",x"635d5d",x"625c5c",x"5f5554",x"645a59",x"685d59",x"5f5755",x"655b5a",x"615b5b",x"605654",x"695a53",x"5b514f",x"655b59",x"655b59",x"625755",x"655a58",x"867971",x"887f7a",x"756860",x"90837b"),
(x"958a84",x"8a7d77",x"99928c",x"908583",x"978e87",x"948b86",x"8a7f79",x"91827b",x"92837c",x"8e7f78",x"938680",x"8d8381",x"645a59",x"595556",x"5d5553",x"5a5657",x"615b5d",x"574f4c",x"504e4f",x"675f5c",x"615755",x"5a5152",x"645c5a",x"5e5654",x"635957",x"5d5958",x"4d4c4a",x"5a5655",x"a09790",x"9a918c",x"9f9490",x"9e948b",x"9c938c",x"988f88",x"9d948d",x"948b84",x"95887f",x"988b82",x"998b82",x"9c938c",x"988d87",x"958880",x"9e9189",x"9a9087",x"615957",x"656162",x"6b5f5f",x"675f5d",x"68605e",x"6b6361",x"665858",x"615652",x"716967",x"5d5958",x"655d5b",x"62534c",x"59514f",x"574c48",x"59514f",x"5a5454",x"877a71",x"95847d",x"837a75",x"968780"),
(x"7c6f67",x"948781",x"968983",x"8d8280",x"948a81",x"8c7d76",x"988984",x"8f8178",x"938980",x"8f8079",x"938884",x"877970",x"6b6162",x"5e5654",x"5d5757",x"585455",x"5d5553",x"58504e",x"615a54",x"645858",x"645a59",x"584e4c",x"5a4c4b",x"625856",x"5f5452",x"56514e",x"504f4d",x"5d5855",x"998f86",x"a09991",x"9b8e88",x"958a84",x"9e9590",x"9b9188",x"9c918b",x"9b9289",x"958d8a",x"998e8a",x"9e948a",x"968d86",x"988982",x"9e918b",x"9a8f89",x"9e9189",x"766c6d",x"626061",x"5c5050",x"6b605c",x"6b615f",x"625453",x"69615f",x"565050",x"5a5552",x"6c6260",x"625a58",x"5a5454",x"605856",x"665b55",x"5f5657",x"635554",x"938680",x"948781",x"8d7e77",x"988e84"),
(x"968b85",x"968981",x"9b908a",x"8b807a",x"8d7f7c",x"938a81",x"a29791",x"9e958c",x"988982",x"93847d",x"a19589",x"978d84",x"645a59",x"5b5555",x"595556",x"615756",x"5e5654",x"5a504f",x"615755",x"5c5452",x"685e5c",x"595556",x"5c5251",x"685b55",x"5f5554",x"575352",x"594f4d",x"5f5651",x"9b9188",x"9a8f89",x"978a82",x"a09694",x"9a918a",x"9c9290",x"958c85",x"9b928d",x"968c83",x"9d928c",x"978c86",x"958a84",x"998c86",x"968d86",x"9b8e86",x"9c9289",x"5e5c5f",x"67625f",x"696566",x"685c5c",x"645653",x"635a5b",x"5e5654",x"5f5755",x"6d645f",x"655b5a",x"605655",x"6a605f",x"5d5553",x"5a5657",x"756158",x"76635f",x"9d8f86",x"9d948d",x"a0938a",x"9c8b84"),
(x"9c8f87",x"9c8e85",x"8d7e77",x"998b82",x"9b8d84",x"a29795",x"9e8f88",x"968b85",x"908279",x"978a82",x"988b83",x"9c8f89",x"5d5354",x"554f4f",x"504a4a",x"665e5c",x"635856",x"665754",x"5d5455",x"584f50",x"585350",x"575352",x"5b5150",x"6c615f",x"5e5550",x"5b5351",x"605855",x"534e4b",x"a09287",x"a0938b",x"a3958c",x"9f9892",x"a69c9a",x"9d9088",x"a2958f",x"a19893",x"9c938e",x"9f958c",x"998e88",x"938886",x"8c837e",x"978a84",x"968885",x"9c938e",x"675c5a",x"736864",x"605758",x"6c6260",x"5b504e",x"5d5352",x"655c57",x"655b59",x"635958",x"625a58",x"625857",x"625a58",x"625857",x"5a585b",x"685e5d",x"5e5453",x"9a8b84",x"93847d",x"8e7d75",x"99887e"),
(x"75645c",x"877368",x"5e5654",x"6e6463",x"665c5b",x"726866",x"766b69",x"605856",x"645a58",x"615b5b",x"59514e",x"66615e",x"928781",x"9b9692",x"8c817d",x"9c958d",x"9b928b",x"95908d",x"938b88",x"999594",x"968f89",x"96918d",x"97908a",x"93867e",x"94877f",x"928781",x"958d8a",x"948a81",x"695b58",x"645e5e",x"6d6362",x"6d625e",x"665c5a",x"615b5b",x"675c5a",x"675f5d",x"7a6760",x"877873",x"665c5a",x"6b5c59",x"6a605e",x"594f4d",x"615957",x"695e5a",x"958a86",x"9d948f",x"9b908a",x"9a8f89",x"988a7f",x"95867f",x"9f928a",x"928781",x"998c83",x"9a8c83",x"9e938d",x"998c84",x"988d87",x"9b8d8a",x"8d847f",x"8f827c",x"6d6865",x"69615f",x"6b615f",x"625a58"),
(x"675c5a",x"544a48",x"615756",x"6a6663",x"6b625d",x"655b59",x"625a58",x"5b5557",x"6a625f",x"665c5a",x"6a5f5b",x"5d5757",x"8d827c",x"8c817d",x"968b87",x"a09790",x"948983",x"8d8078",x"8d8078",x"8f8480",x"908886",x"998e8a",x"948b86",x"8f867f",x"9b918f",x"968d88",x"8e8580",x"8e8381",x"6b6766",x"5b4f4f",x"615756",x"645c59",x"6a5e5e",x"675956",x"726763",x"635957",x"655a58",x"74635c",x"615957",x"5f5755",x"645b5c",x"5a5454",x"5d5855",x"665d58",x"9b8c85",x"a09695",x"a0958f",x"9e9188",x"9b908a",x"9b8e86",x"9a8d87",x"90837b",x"968981",x"968c83",x"988d87",x"9a8d87",x"968d88",x"9b8c85",x"958379",x"9a9087",x"57524f",x"635957",x"7e6c62",x"524847"),
(x"655d5b",x"6e6462",x"645c5a",x"6f625a",x"6d625c",x"5f5755",x"695f5d",x"645e5e",x"615859",x"665b57",x"645c59",x"635b59",x"91847c",x"9d938a",x"a09896",x"958a84",x"978e89",x"958b89",x"8f8681",x"97928f",x"99918e",x"9d948d",x"93867e",x"948983",x"938884",x"938b88",x"968d88",x"928783",x"6e6463",x"594f4d",x"645a58",x"6a605e",x"85726b",x"76655e",x"685952",x"645c5a",x"58504e",x"625857",x"625c5c",x"6f6564",x"5f5353",x"4f4949",x"62595a",x"595353",x"9b8e86",x"a09792",x"9e9087",x"90837d",x"928179",x"8e837d",x"9e938d",x"9a8d85",x"968981",x"978980",x"8e817b",x"958c85",x"93857c",x"968981",x"988e85",x"9a928f",x"52494a",x"584e4d",x"8e807f",x"675c5a"),
(x"736a65",x"605856",x"5d585c",x"545051",x"625c5c",x"6c6260",x"675f5d",x"615853",x"645c5a",x"6b615f",x"5e5a5b",x"685e5d",x"999491",x"9a8e82",x"9d928c",x"7f7979",x"9b918f",x"968c83",x"958c87",x"a69790",x"9a918a",x"999089",x"968b87",x"948985",x"978f8c",x"918a84",x"8d827e",x"958f8f",x"675e5f",x"5e5453",x"5e504f",x"6a6260",x"6e6262",x"6d6563",x"5f5755",x"675c58",x"575556",x"675f5d",x"5e5654",x"685d5b",x"5a5250",x"665c5a",x"605654",x"5a5250",x"9a8c83",x"9b9187",x"a0968c",x"837872",x"91837a",x"90817a",x"807061",x"9a908e",x"918174",x"9d9088",x"9b8f83",x"95867f",x"968980",x"978e87",x"95877e",x"9a8d85",x"605856",x"594f4e",x"85726b",x"605654"),
(x"635957",x"635b59",x"665c5b",x"5f5755",x"695f5e",x"726a67",x"675c58",x"564b47",x"655d5a",x"655653",x"686463",x"675d5b",x"938b88",x"94867d",x"998e88",x"8b8380",x"90837b",x"90837b",x"9c8e8d",x"988e85",x"968d86",x"938980",x"978f8c",x"968980",x"928783",x"968d88",x"948b84",x"948985",x"635957",x"655a58",x"685e5c",x"69615e",x"756a66",x"6f6563",x"6c6462",x"5c5452",x"524e4d",x"615b5b",x"665c5a",x"5e5653",x"58504e",x"625755",x"6b6160",x"5c5452",x"988e85",x"9a8d85",x"978c86",x"81746e",x"92837c",x"8f8079",x"99918f",x"5b504a",x"726159",x"92847b",x"9a8d85",x"968b85",x"918078",x"928781",x"948987",x"938884",x"615654",x"70655f",x"75665f",x"6c6260"),
(x"786a61",x"675d5b",x"635b59",x"635d5d",x"685f60",x"686360",x"655d5b",x"685e5c",x"565251",x"605758",x"5a5152",x"665e5c",x"9d9088",x"9a8f89",x"9a8d84",x"908279",x"988982",x"9a9592",x"8b807a",x"938882",x"9a908e",x"928781",x"968885",x"938a83",x"8b827d",x"8f827a",x"908c8b",x"908b88",x"6a6162",x"6d625e",x"80726f",x"756663",x"796e68",x"736562",x"6c5c5c",x"5a5250",x"56514e",x"5a5152",x"58504e",x"5b5555",x"5f5553",x"5e534f",x"635957",x"605654",x"a19996",x"9c9289",x"93867e",x"92857d",x"5b5148",x"948b86",x"988f8a",x"998c86",x"948983",x"9d9088",x"978e87",x"999089",x"9b908a",x"978a82",x"988b83",x"a89c9c",x"584e4c",x"665e5b",x"685e5c",x"5a5657"),
(x"645c59",x"6f6765",x"6a6162",x"5c5a5b",x"565455",x"585657",x"675d5b",x"595353",x"685e5c",x"625856",x"666263",x"625c5c",x"918d8a",x"8f827a",x"938a83",x"7f7979",x"968980",x"999491",x"8c8280",x"968b85",x"9e9590",x"999089",x"988f8a",x"9c938e",x"948b86",x"908684",x"918b8b",x"948f8b",x"847474",x"847570",x"857373",x"847570",x"7f706d",x"766865",x"594f4e",x"5f5755",x"494343",x"615555",x"615654",x"594f4d",x"595051",x"615755",x"615956",x"766865",x"988b82",x"94877f",x"94877f",x"9f928a",x"988d89",x"8f8480",x"9a918a",x"999089",x"988f88",x"978a81",x"948a81",x"9b8c85",x"988e85",x"978e89",x"978c86",x"918682",x"645955",x"685e5c",x"6a605e",x"72685f"),
(x"706561",x"6d625e",x"676362",x"6a6665",x"605a5a",x"59504b",x"605655",x"5a5250",x"605a5a",x"6d6361",x"6f615e",x"665b55",x"9b908c",x"98908d",x"9b908c",x"938e8a",x"948983",x"90837b",x"8d847f",x"978e87",x"9a938d",x"8e817b",x"99908b",x"8f8480",x"918883",x"9b9187",x"7b797c",x"8e837d",x"786d6b",x"7d6f6c",x"796f6d",x"685e5c",x"726b65",x"6c6260",x"615755",x"645655",x"5f5a57",x"5f5452",x"5c514d",x"625a58",x"645a58",x"5d5351",x"675d5b",x"625755",x"a0958f",x"9d948f",x"988b83",x"9d928c",x"9a8f89",x"948b86",x"998e88",x"988e8c",x"9c9491",x"9c8f86",x"948b86",x"928783",x"9b9391",x"948b84",x"9d9290",x"9f9794",x"5b5150",x"695f5e",x"615c59",x"7f6f62"),
(x"8d8078",x"685e5d",x"665b57",x"6e6868",x"6c615f",x"5d5757",x"665c5b",x"675c5a",x"5f5554",x"6b6361",x"646061",x"67625f",x"938882",x"918a84",x"958e86",x"938680",x"9f9289",x"8f857c",x"8f827a",x"91827d",x"a39e9b",x"92847b",x"8b807a",x"857d7a",x"8b7c77",x"8f8687",x"9a9697",x"92857f",x"655b5a",x"796e6c",x"766b67",x"726763",x"6a605e",x"665e5c",x"645a59",x"524a47",x"59514f",x"4e4a4b",x"736a65",x"615755",x"584e4d",x"5b514f",x"635856",x"665c5a",x"a1948c",x"9f928a",x"9f948e",x"958880",x"968b85",x"92857d",x"9d8f86",x"9b8e86",x"978e89",x"988f88",x"9b8e86",x"968d88",x"8f8180",x"9c9290",x"9b9188",x"988f88",x"635856",x"69625a",x"78665a",x"655b5a"),
(x"675d5c",x"746c6a",x"706762",x"655d5b",x"6b615f",x"7b706e",x"635f5e",x"635e5b",x"625a57",x"6b625d",x"635a55",x"5d5455",x"9a9693",x"9c9793",x"958c87",x"948c89",x"887e7c",x"8b7e78",x"90837b",x"8e8179",x"8d827c",x"938a83",x"948987",x"9a9290",x"91847c",x"998c84",x"948b84",x"847a79",x"6f6563",x"756b6a",x"666465",x"68605e",x"5e5654",x"6f6566",x"645e5e",x"58504e",x"605655",x"776a62",x"594f4e",x"695e5a",x"5d5553",x"5c5451",x"685d5b",x"5c5452",x"978980",x"94867d",x"958578",x"988a81",x"908071",x"988a81",x"998c86",x"807061",x"9d948f",x"9a918a",x"a09591",x"988b85",x"928886",x"978e87",x"9e9693",x"998e8a",x"625856",x"816f6b",x"7a7067",x"635b59"),
(x"716765",x"675e59",x"6b6361",x"746a68",x"645e5e",x"736d6d",x"716765",x"686262",x"635957",x"666060",x"675f5c",x"837977",x"918d8c",x"948b84",x"887d77",x"9d9391",x"94877f",x"928781",x"8c7e75",x"8f8079",x"958880",x"9b9693",x"938b89",x"968e8b",x"938a85",x"968c8a",x"918785",x"988f8a",x"6e6462",x"6a6464",x"6c6364",x"6a6260",x"5f5659",x"5d5151",x"5d5351",x"5e5452",x"685e5c",x"675d5b",x"786d69",x"6d625e",x"605654",x"685e5c",x"625857",x"625a58",x"9a9188",x"948983",x"9b908a",x"9b8f83",x"9c8e85",x"95877e",x"958880",x"9e948a",x"a0938b",x"978c86",x"978e87",x"9d928c",x"958784",x"968885",x"978e87",x"998f86",x"6b6160",x"7c6e65",x"84776f",x"716765"),
(x"6f6462",x"646061",x"665c5a",x"6f6563",x"696061",x"6a6260",x"6c6462",x"666060",x"665c5a",x"635f60",x"676161",x"716765",x"978c86",x"958a86",x"978881",x"8c7d76",x"8e8482",x"928781",x"6a5c53",x"9b908c",x"887f7a",x"988f88",x"8b807a",x"948b86",x"8b7e78",x"8f8583",x"948b86",x"9b908a",x"726867",x"726763",x"6a605e",x"665e5c",x"675c5a",x"665e5c",x"5b5351",x"605553",x"605655",x"706664",x"655c57",x"746761",x"6e635d",x"6f625c",x"6f655b",x"6a605e",x"998b82",x"9b8d84",x"a09289",x"9e9087",x"90765f",x"97897e",x"92847b",x"a1948e",x"9f9387",x"9e8d86",x"a39a95",x"9d9592",x"958b89",x"948e8e",x"938882",x"988f8a",x"6e6462",x"7e746b",x"685e5d",x"65605d"),
(x"676161",x"6a6260",x"605855",x"6c6764",x"656160",x"676163",x"6f6969",x"786e6d",x"685e5c",x"69615e",x"696363",x"5f5b5c",x"90857f",x"958880",x"988f8a",x"92857d",x"8e8077",x"837268",x"968b85",x"918a82",x"959192",x"988f8a",x"8f8785",x"8f8480",x"8e817b",x"90857f",x"90837b",x"91877e",x"6c6462",x"7a706f",x"64605f",x"635958",x"6d6361",x"5e5556",x"5b5150",x"473f3c",x"6c615f",x"675f5d",x"7d7067",x"635957",x"675c56",x"6f6661",x"776861",x"695b52",x"9d9088",x"a19184",x"a0968d",x"a4958e",x"9b8d84",x"a1948b",x"978b7f",x"9d8f86",x"998b7e",x"a19690",x"968981",x"9a8b84",x"9e958e",x"978e87",x"9b908c",x"9b928b",x"6a605f",x"716360",x"615957",x"615d5e"),
(x"726761",x"6c615f",x"625e5d",x"7c7472",x"686262",x"666060",x"655d5b",x"685e5d",x"605856",x"726866",x"5c5250",x"69615f",x"8c817b",x"92857f",x"968885",x"998e8a",x"928785",x"897f76",x"8d8381",x"948b86",x"92857f",x"86817e",x"948a8b",x"8f8480",x"89807b",x"817775",x"9a918c",x"938680",x"686262",x"6c6364",x"686465",x"696564",x"665e5c",x"665b59",x"6a605f",x"635a5b",x"5e5452",x"675d5b",x"726765",x"5e5556",x"554a46",x"726765",x"726765",x"665e5c",x"9d9087",x"998c84",x"958a84",x"a1948c",x"978c86",x"9f9691",x"918680",x"91827b",x"99887e",x"93847d",x"9f9691",x"9c9491",x"9d8f86",x"9d9087",x"9f9593",x"9e958e",x"635b59",x"786d6b",x"786b65",x"645a59"),
(x"6c6461",x"726866",x"645e5e",x"686360",x"635e5b",x"635e5b",x"776c68",x"68605e",x"6b6663",x"6d6260",x"5d5455",x"62595a",x"988b83",x"9b948c",x"978c88",x"988b85",x"978e89",x"75685f",x"8f8784",x"8c8481",x"877e7f",x"8f8482",x"847c7a",x"888282",x"8a7f79",x"93847d",x"8f8583",x"7e7168",x"6a6667",x"666263",x"7f7a7e",x"796f6e",x"6e6462",x"696564",x"6c6764",x"706866",x"776f6d",x"6d6361",x"7c7374",x"6b6360",x"766b69",x"6a605f",x"6e615b",x"5b504c",x"9f9490",x"9d9088",x"988f88",x"9d9087",x"a1938a",x"a19690",x"91837a",x"8e7c70",x"9c8f86",x"9f928c",x"8f8079",x"9a897f",x"988b83",x"988b85",x"958a86",x"9c938c",x"665d5e",x"736866",x"6a6162",x"68605d"),
(x"695b58",x"766b67",x"786f70",x"696061",x"726a68",x"766c6b",x"6a6162",x"665b59",x"6b6263",x"695f5e",x"665855",x"686264",x"9f8e84",x"887972",x"92857c",x"928781",x"9f9089",x"9c9897",x"8d827c",x"978e89",x"948781",x"968c83",x"8b8180",x"978d84",x"8e7f78",x"928984",x"918889",x"8b807c",x"6a605e",x"6c6261",x"766b69",x"74706f",x"706866",x"736b68",x"776f6d",x"6c615f",x"736967",x"756b69",x"716360",x"736967",x"746965",x"69615f",x"6f6563",x"645a58",x"a19690",x"aba19f",x"958c85",x"8e8179",x"998c84",x"948b86",x"897c73",x"968d84",x"a09591",x"9c9491",x"978c88",x"91847e",x"938987",x"97928f",x"928d8a",x"9a8f8b",x"786d69",x"706961",x"534f4e",x"686262"),
(x"84776f",x"7f766f",x"786d69",x"8d807a",x"8e817b",x"8e837f",x"7d746f",x"8b7e76",x"7f726a",x"847b76",x"847b72",x"817775",x"554c4d",x"72645b",x"5c5354",x"554f4f",x"534e4a",x"514d4c",x"4f4b4a",x"564e4c",x"605553",x"645953",x"5c5859",x"8e755f",x"67625f",x"6c6970",x"5c5354",x"514947",x"958c87",x"988e85",x"998c86",x"958d8b",x"8c7d76",x"9a9290",x"9b948e",x"998b82",x"938884",x"8a7f79",x"958a84",x"8e8482",x"968e8b",x"8b827d",x"8a7f7b",x"968e8b",x"625856",x"605553",x"4f4744",x"534b49",x"5d5351",x"5e5452",x"615957",x"5c5251",x"6d645f",x"534f50",x"625753",x"544c49",x"6c5f59",x"494748",x"4c4a4d",x"535355",x"8e8179",x"867971",x"887d77",x"7c6f67"),
(x"877871",x"897b72",x"877a72",x"8f847e",x"8c837e",x"8e837f",x"8c817b",x"897e78",x"8a7d75",x"867971",x"897e78",x"817670",x"605b58",x"696661",x"5b5350",x"625954",x"62554d",x"5c5250",x"6c5f59",x"6d6058",x"4e4c4d",x"514e49",x"4a4849",x"4e4a47",x"56514e",x"504e4f",x"5b5350",x"4d4948",x"8e837d",x"90817a",x"92837c",x"897e7a",x"978e85",x"8c8885",x"99928a",x"9a918c",x"998c83",x"95928d",x"908885",x"908782",x"9d9592",x"958d8b",x"938b88",x"978980",x"6c6461",x"6a5d57",x"584e4f",x"534b49",x"61544e",x"605654",x"6e6055",x"72655d",x"675f5c",x"645b56",x"685d59",x"5c5a5b",x"625e5d",x"56555a",x"535257",x"515055",x"8d7f76",x"8c7e75",x"897c74",x"8a8077"),
(x"8a7d75",x"8f827a",x"84776f",x"8d827c",x"887d77",x"827771",x"817672",x"85766f",x"877a72",x"867971",x"84756e",x"7e7371",x"5e534d",x"625d5a",x"565455",x"675c56",x"796c64",x"635a55",x"574c48",x"554b49",x"65615e",x"5c5452",x"4c4849",x"59514f",x"4b4748",x"615c59",x"585657",x"5e5956",x"8c7f77",x"96887f",x"998c84",x"9b928d",x"988e85",x"958a86",x"9b8a82",x"93867e",x"9b8b7e",x"938680",x"9e9993",x"958a84",x"928a88",x"857a74",x"8d827c",x"8b807a",x"5c5d5f",x"706865",x"635958",x"594f4d",x"605551",x"6a605e",x"685b55",x"71635a",x"7f6d5f",x"665b57",x"83756a",x"686360",x"5b5b5d",x"5a5b5f",x"5c5d61",x"545358",x"92857d",x"877871",x"93847d",x"8a7d75"),
(x"756860",x"867973",x"887770",x"8e8179",x"7d726c",x"847973",x"7f726c",x"847973",x"847975",x"837874",x"7a6d65",x"827974",x"524c4c",x"504846",x"5a5454",x"5f5b58",x"5c5250",x"60564d",x"574e49",x"5c5249",x"514c49",x"4b4341",x"594f4d",x"4b4642",x"504c49",x"575352",x"514f50",x"4a4647",x"9a918a",x"9c8f87",x"96887f",x"9f9188",x"94857e",x"968e8b",x"99928c",x"978a82",x"918076",x"9e958e",x"9f948e",x"a69f99",x"8e837f",x"9b9693",x"8d827e",x"867770",x"555356",x"5d5b5c",x"625e5d",x"5f5b5a",x"5c5250",x"625753",x"635854",x"695e5a",x"67594e",x"5d5c5a",x"83746d",x"7f7168",x"4b494a",x"484848",x"4f4f51",x"545456",x"91847c",x"837970",x"887972",x"92857d"),
(x"887b73",x"8b7c75",x"817670",x"8c7f77",x"8e8179",x"887d79",x"887b73",x"877c76",x"847975",x"877c76",x"7d726c",x"827773",x"4e4946",x"5c514b",x"645d57",x"656160",x"645f5b",x"6a5f59",x"4c4847",x"564b49",x"443c3a",x"48403d",x"524d4a",x"545255",x"5e5654",x"575757",x"514d4e",x"534f4e",x"9a9087",x"93908b",x"9b9188",x"998c84",x"958880",x"9a8f8b",x"9b8d84",x"92887f",x"989390",x"9c9491",x"93867e",x"8d827c",x"867770",x"95908c",x"9b908c",x"7b706a",x"525358",x"5d5c61",x"5e5c5d",x"5f5f5d",x"5c5250",x"5c5250",x"5f5452",x"605553",x"625954",x"847a71",x"776758",x"75675c",x"525254",x"5f5452",x"58504d",x"62554f",x"968782",x"867b75",x"8c7e75",x"897c74"),
(x"857870",x"887972",x"8a7d75",x"92857d",x"867971",x"92857d",x"877a72",x"847977",x"887f7a",x"837874",x"847973",x"817672",x"595353",x"716059",x"636260",x"6a5f5b",x"5b5b5b",x"4f4b4a",x"4c4849",x"584e4c",x"5a4f4b",x"5f524c",x"574d4b",x"635e5b",x"5b5555",x"565455",x"555150",x"5b5653",x"958880",x"9f958c",x"a29992",x"a2958c",x"9a918a",x"9a9592",x"9f9a97",x"a29791",x"998e8a",x"a0968d",x"93867e",x"91827b",x"8f8079",x"968e8b",x"92887c",x"968277",x"4f5055",x"57565b",x"555459",x"595959",x"5c5250",x"584e4c",x"514946",x"74635c",x"71645c",x"7a6c5f",x"7a6d65",x"5f5b5a",x"635a55",x"7b6859",x"6b625d",x"695b4e",x"998c86",x"8b7a72",x"8d8078",x"8e7f78"),
(x"83766e",x"83746d",x"877a72",x"897b72",x"897c74",x"8d807a",x"857a74",x"837876",x"897e7a",x"8c8280",x"887d79",x"7f7573",x"554b49",x"605b58",x"524e4d",x"534e4a",x"6b5c55",x"5f5754",x"5f5651",x"645a58",x"5c5451",x"554d4b",x"333335",x"655852",x"69554a",x"564e4c",x"545253",x"5d5250",x"9e8f88",x"9d948d",x"9e9590",x"92887e",x"a19388",x"a49993",x"9b8e86",x"a69790",x"9b908a",x"998c84",x"9e9189",x"9e948b",x"978c86",x"9f9892",x"928d8a",x"92857c",x"56575b",x"5c575b",x"504e4f",x"655852",x"595051",x"584f4a",x"5b504a",x"756359",x"7b6d62",x"615b5d",x"726459",x"675c56",x"605752",x"665f59",x"574c46",x"6f625a",x"95877e",x"908279",x"8f8079",x"8e8077"),
(x"897a73",x"8e8077",x"91827d",x"8a7b74",x"8d7e79",x"8f827a",x"8b7e76",x"8b817f",x"857a74",x"837874",x"7c7270",x"857b7a",x"5c534e",x"544f4c",x"5b5351",x"5f5651",x"554b49",x"645f5c",x"665e5b",x"675d5b",x"594f4d",x"5d5757",x"554f4f",x"544c4a",x"6b5e58",x"5e514b",x"5b504e",x"4d494a",x"9b8e88",x"a19690",x"978e89",x"918682",x"988d87",x"a29992",x"a89992",x"a39592",x"a39a95",x"988f8a",x"9c938c",x"9d9088",x"928d8a",x"968d88",x"938d8d",x"897a73",x"4f4d4e",x"545253",x"504e4f",x"57524f",x"6d5f54",x"635a55",x"5b5351",x"857464",x"62554f",x"5c514f",x"7b6a60",x"655c57",x"6e5f5a",x"6b5d54",x"695c56",x"5c5859",x"978c86",x"91837a",x"8b7e78",x"8a7b74"),
(x"877871",x"7c7676",x"8b7d72",x"837872",x"8d8078",x"86786f",x"8c7f77",x"7d6f64",x"7d726e",x"857774",x"7f746e",x"827773",x"565251",x"71645c",x"615853",x"695851",x"615957",x"5b595a",x"655c57",x"585453",x"574f4c",x"4e4a4b",x"5b5653",x"5d5352",x"5c514d",x"574f4c",x"695a53",x"554b49",x"8b827d",x"9a9087",x"918078",x"9e958e",x"a4a09f",x"a59c97",x"ab9e96",x"a69991",x"a69d98",x"9a9087",x"9c918b",x"9c938e",x"988e8c",x"907f75",x"8f8079",x"928783",x"655d5a",x"565455",x"555150",x"645955",x"655b59",x"635957",x"5f554c",x"635854",x"574d4b",x"6d5e57",x"645a51",x"6a625f",x"6a6057",x"5c4e4e",x"63564e",x"6b5e56",x"988b85",x"8a7c71",x"8d827c",x"94877f"),
(x"90857f",x"8b7c75",x"92847b",x"847973",x"807571",x"80756f",x"827775",x"837a75",x"8b827d",x"89807b",x"766961",x"827773",x"685d59",x"615652",x"675956",x"5d5455",x"665d5e",x"59575c",x"605856",x"675f5c",x"5e5556",x"5d5351",x"5f5450",x"695b52",x"605752",x"796860",x"665b55",x"554c45",x"968d86",x"96887d",x"9a8b84",x"9e9590",x"a89d97",x"9b948e",x"a49993",x"9b928b",x"9e938d",x"a09790",x"989189",x"938a85",x"988f88",x"84776f",x"897c73",x"8b796d",x"7f7166",x"665e5b",x"514946",x"625857",x"71645e",x"73655c",x"807269",x"705f57",x"665951",x"7a6c61",x"434240",x"5c5451",x"534b49",x"534d4d",x"574e49",x"534844",x"908279",x"8f8079",x"857872",x"968b87"),
(x"82756d",x"8f8079",x"8f8178",x"867971",x"80736b",x"82756f",x"847771",x"827771",x"837872",x"827773",x"81746e",x"786d69",x"554a48",x"585350",x"5c5754",x"575350",x"59514f",x"605654",x"615756",x"55504d",x"5d5855",x"524a47",x"544c4a",x"575151",x"5f524c",x"5e534f",x"66554d",x"5e534f",x"9d9392",x"96857d",x"8a8077",x"a09993",x"9a9086",x"9a9591",x"938a85",x"a0958f",x"9d948d",x"9c918b",x"968f87",x"9b9188",x"94867d",x"918682",x"8b7a70",x"978e89",x"514f50",x"635d5d",x"6b6158",x"5d5351",x"736258",x"5e534f",x"7b6859",x"766659",x"776a61",x"74635b",x"584a49",x"58504d",x"58504d",x"584e4c",x"5e5452",x"5e5351",x"91837a",x"8e7f78",x"877970",x"8e7d73"),
(x"90837b",x"887b75",x"8c7e75",x"90817a",x"817672",x"8c7d76",x"887b75",x"837874",x"807571",x"83766e",x"82756f",x"89807b",x"46423f",x"444243",x"6d625c",x"6e5f58",x"5a514a",x"5b5557",x"615c59",x"5e5550",x"5c5250",x"5e5452",x"544b4c",x"564e4c",x"64554e",x"554d4a",x"554d4b",x"524a47",x"9a8e82",x"8b7c75",x"938b88",x"928783",x"948983",x"a09b97",x"958d8a",x"9d948f",x"918883",x"998e88",x"928984",x"9d948d",x"928179",x"99908b",x"887f7a",x"9b9693",x"7a6c63",x"6c635c",x"483e32",x"524846",x"604d3f",x"7d746f",x"67564f",x"625856",x"77665c",x"837061",x"61524b",x"534947",x"4e4443",x"70625f",x"5b5350",x"836d5f",x"9b8e86",x"8a7c73",x"897c74",x"8b7e76"),
(x"81746e",x"8d7e77",x"8c7d76",x"8c8279",x"85766f",x"877a72",x"897f76",x"93867e",x"786d67",x"7b706c",x"7b706a",x"81746e",x"59514f",x"4c4847",x"635856",x"5d5553",x"73655a",x"615654",x"615859",x"6f6158",x"685e5c",x"534a4b",x"5e534f",x"59504b",x"685a51",x"625656",x"5b5351",x"514745",x"908684",x"92857c",x"8c817d",x"8e857e",x"8e8580",x"8c8783",x"8e8683",x"99918e",x"999089",x"97928f",x"918986",x"91847c",x"867770",x"84776f",x"8d7f7c",x"8f8583",x"595451",x"74655e",x"635c56",x"635a55",x"7f6860",x"817162",x"5c5250",x"484647",x"4f4b4c",x"7c6a5e",x"635950",x"72635c",x"504845",x"6c5f59",x"675851",x"675e55",x"9c8e85",x"8e8077",x"897c74",x"897f76"),
(x"8d8078",x"83766e",x"83746d",x"7e7169",x"8b7d74",x"837670",x"8c7f77",x"8e8179",x"7e736d",x"857872",x"80766d",x"837977",x"625954",x"5b524d",x"635a55",x"68574f",x"635957",x"68605e",x"6b6768",x"62534e",x"655b59",x"655a58",x"635d5d",x"5c5857",x"615756",x"635a5b",x"5c514d",x"6f6661",x"9f968d",x"999089",x"958c85",x"92837e",x"978f8c",x"958a84",x"807772",x"918682",x"938582",x"857872",x"8c7d76",x"91847e",x"8f847e",x"8d7e79",x"938376",x"8f827c",x"6c6260",x"6a615a",x"5e5550",x"7a685c",x"736258",x"856f62",x"5e574f",x"76685d",x"826f61",x"5e5550",x"5d5352",x"564b49",x"584d4b",x"655a54",x"504a4a",x"685a51",x"94867d",x"96857b",x"857671",x"8b807a"),
(x"8a7f79",x"877c78",x"81746c",x"897c76",x"857a76",x"796e68",x"8d807a",x"857870",x"7e7371",x"8d827c",x"7e7371",x"7a706e",x"514745",x"615652",x"6a5b54",x"756253",x"6b6263",x"5f5554",x"645858",x"645b54",x"675d5c",x"58504d",x"585453",x"615755",x"565457",x"615b5b",x"4c4a4d",x"706963",x"978a82",x"8d8280",x"7a6d65",x"948781",x"91837a",x"827167",x"897b70",x"81726b",x"8a7972",x"83746d",x"81746e",x"928481",x"928783",x"887b73",x"8e857e",x"867973",x"6b6263",x"7c6b61",x"88786b",x"867160",x"685954",x"88766a",x"6b5a53",x"716056",x"594f46",x"615956",x"6d6968",x"574e49",x"6d5e57",x"615c59",x"645953",x"524d4a",x"9e9188",x"92837c",x"7e736d",x"867d78"),
(x"7e7371",x"82756d",x"84776f",x"8c7f79",x"74655e",x"8c817b",x"8b807c",x"8f847e",x"8d827e",x"81776e",x"6c635e",x"867c7b",x"84736b",x"665d58",x"806e64",x"675a54",x"705d56",x"555150",x"5f5554",x"59514f",x"6b5957",x"695e5a",x"5d5552",x"56514e",x"5c5452",x"67605a",x"5f5d5e",x"6e6158",x"908b88",x"938b88",x"8d827c",x"837872",x"908684",x"8e837d",x"91847e",x"92837c",x"90837b",x"94877f",x"90857f",x"90837d",x"978f8d",x"8a7f7b",x"90837b",x"8c7b71",x"60554f",x"796861",x"746152",x"645957",x"614f43",x"7f685a",x"73645d",x"5d5855",x"615652",x"6a5f59",x"584942",x"6c615b",x"655a56",x"64574f",x"615853",x"575757",x"948983",x"8e7f7a",x"877c78",x"857a78"),
(x"4d4747",x"6e5c58",x"6a5f5d",x"655a56",x"5f5554",x"645c59",x"625857",x"585453",x"5f5b5a",x"5b5555",x"5b5351",x"625857",x"7e756e",x"837977",x"8e817b",x"8e8179",x"90817a",x"897a73",x"8e8179",x"908782",x"94877f",x"8b7e76",x"897f7d",x"8c8784",x"978c86",x"958d8a",x"8a7f7b",x"8d8078",x"6c6462",x"615755",x"655b5c",x"62584f",x"5e5452",x"5e5956",x"5e5956",x"635856",x"635a55",x"7a6d64",x"888687",x"74675f",x"73615d",x"7e6c5e",x"79695c",x"6e5f5a",x"94857e",x"8c7e75",x"91827b",x"938278",x"988b82",x"8c7d76",x"94867b",x"8f827a",x"8b7d7a",x"8f8279",x"8e837d",x"8f827a",x"8c7f76",x"877c78",x"877c78",x"8b827d",x"695f5d",x"615755",x"655f5f",x"5a5657"),
(x"675c58",x"695753",x"6b6160",x"6c5e5b",x"60554f",x"726964",x"605856",x"544b4c",x"544e50",x"565251",x"5f5b5a",x"5b5557",x"80736d",x"887f7a",x"8f8681",x"84756e",x"8f827a",x"988e85",x"90837d",x"958784",x"8f847e",x"867e7b",x"928781",x"877c78",x"92857f",x"948985",x"7c7270",x"80726f",x"4b494a",x"484443",x"514d4c",x"5c5451",x"5d5855",x"4b494a",x"5b5350",x"70635a",x"675f5d",x"645957",x"5d5553",x"4d4946",x"55504d",x"4e4c4f",x"545454",x"6d625e",x"998b82",x"8f847e",x"938278",x"968780",x"968c8b",x"91837a",x"93847d",x"8c7f79",x"8f8079",x"8f8178",x"8f827a",x"867971",x"877c76",x"918378",x"958882",x"8e7f78",x"695f5e",x"584e4c",x"564d50",x"5a5552"),
(x"675d5b",x"67524d",x"6d5e57",x"675555",x"726866",x"5d5958",x"494748",x"635957",x"54504f",x"5f5959",x"5a5152",x"5e585a",x"8b7d74",x"898481",x"807875",x"897c74",x"958880",x"8f827a",x"847268",x"877a74",x"887e7c",x"7d7371",x"8d827c",x"8e847b",x"877c76",x"887b75",x"887d79",x"7b7168",x"5c5859",x"555658",x"5d5352",x"595556",x"504c4b",x"665d58",x"74675f",x"675f5d",x"605655",x"6e5f58",x"5b595a",x"59575a",x"59575a",x"5c5c5e",x"6a5d57",x"746359",x"90837b",x"8d8077",x"8b7c77",x"93867e",x"948379",x"9a908e",x"90817a",x"948983",x"877c78",x"88776d",x"887b73",x"857870",x"867971",x"7e7570",x"7f726c",x"81726b",x"625656",x"59514f",x"554c4d",x"5a5454"),
(x"6c6060",x"75625b",x"6c5c5c",x"5f5553",x"5e5453",x"504846",x"635957",x"5d5351",x"5f5b5a",x"4e4946",x"5c5452",x"5e5453",x"796c64",x"8b7e76",x"897a73",x"8f8583",x"958880",x"7d726e",x"857c77",x"827974",x"938f90",x"918680",x"7e736d",x"90837b",x"92857d",x"837670",x"7b706a",x"8c817d",x"4f4f4d",x"514e49",x"64605f",x"535154",x"585657",x"625a58",x"807063",x"796a63",x"635e5b",x"514b4b",x"5b5a58",x"565553",x"675c56",x"78645b",x"70635b",x"595355",x"9c9290",x"908581",x"92857d",x"8f827a",x"91827d",x"9a8981",x"8d7e77",x"988e8c",x"8e847b",x"97867e",x"958b82",x"84776f",x"897b70",x"8a7f7b",x"8c7f77",x"8f7e76",x"5e5654",x"574f4d",x"645b56",x"675d5c"),
(x"665c5a",x"726360",x"6e605d",x"5c5250",x"5c5251",x"615b5b",x"675d5b",x"635e5b",x"635f5c",x"685d5b",x"605c5d",x"5b504e",x"7a6d67",x"867973",x"8d807a",x"867d78",x"918680",x"928781",x"948781",x"8c7d76",x"8b817f",x"958880",x"877c76",x"867b77",x"90867c",x"7e736d",x"877a72",x"948b86",x"6f625c",x"7e7067",x"6c6261",x"6c6260",x"7a716c",x"635b58",x"6a5d57",x"7e7266",x"5e5858",x"6e6463",x"535152",x"554f51",x"595353",x"615b5b",x"645a58",x"57524f",x"9d8f86",x"988e84",x"93867e",x"8f847e",x"8e8077",x"8e7d73",x"928177",x"8c8481",x"8f8279",x"978980",x"978a84",x"8c7e75",x"857369",x"8c7f77",x"897e78",x"8e8179",x"574d4e",x"60524f",x"5e5a5b",x"5f5554"),
(x"695b58",x"615957",x"635854",x"665c5a",x"615756",x"5e5654",x"595556",x"645f63",x"575556",x"585453",x"5d595a",x"5f5b5a",x"7b6e66",x"8e8179",x"8c7d76",x"90857f",x"817670",x"94877f",x"8a7d77",x"8e837d",x"887b73",x"8d8078",x"8d827c",x"93847d",x"8e837d",x"7f7470",x"898079",x"938a85",x"7c6861",x"5b595c",x"616163",x"504e51",x"65605c",x"5d5855",x"6e635d",x"615650",x"4d4b4c",x"565457",x"6a6260",x"575759",x"595451",x"6b5e58",x"726056",x"585254",x"9b8d84",x"97867e",x"958a86",x"8c817d",x"93857c",x"8e7f78",x"8c7e75",x"958b89",x"908277",x"887d77",x"8f857c",x"96887f",x"97897e",x"867770",x"6f6661",x"92817a",x"5e5654",x"635a5b",x"584e4d",x"6c6462"),
(x"565455",x"635f5e",x"595554",x"6e635d",x"655b59",x"69615f",x"5a5657",x"746b66",x"645c5a",x"5f5b5a",x"5a5657",x"5a5454",x"83766e",x"92887f",x"928781",x"92837c",x"93867e",x"887d7b",x"8b7e76",x"8b7d74",x"8e8179",x"857a74",x"897e78",x"877a71",x"857870",x"84756e",x"877c76",x"8c837e",x"5c5c5e",x"6f6a67",x"5f5d60",x"5d5b5e",x"524c4c",x"545358",x"57585c",x"736660",x"535152",x"4a494e",x"535152",x"605454",x"685f5a",x"655d5b",x"443f43",x"584a49",x"9a908e",x"948983",x"877970",x"95847c",x"978a82",x"998f86",x"8f7e74",x"918076",x"8e7f78",x"8e8381",x"8f8178",x"918078",x"8c7e7b",x"91837a",x"91847c",x"897c76",x"615957",x"5d5757",x"655b59",x"635958"),
(x"4e4a4b",x"524e4d",x"595556",x"58504e",x"665c5a",x"665c5a",x"565050",x"615853",x"746967",x"5a5454",x"655b59",x"65524b",x"8f8178",x"91827b",x"897e7a",x"867971",x"90837d",x"8f8079",x"89807b",x"8c7f76",x"958a84",x"867973",x"867b77",x"7a6d65",x"887b73",x"8a7d75",x"8c7f77",x"8a7d75",x"595554",x"616163",x"696564",x"57565b",x"5b595c",x"726a67",x"514f50",x"655b5a",x"545255",x"585350",x"605856",x"534e4a",x"535250",x"685d5b",x"565455",x"605b58",x"95867f",x"978a82",x"918378",x"8b7871",x"86786f",x"938987",x"897c76",x"746153",x"948278",x"968780",x"968b87",x"908279",x"8d8078",x"9c938e",x"938b89",x"8d847f",x"585252",x"675c5a",x"4a4444",x"5f5657"),
(x"585453",x"555150",x"555152",x"5c5754",x"605758",x"645b5c",x"605758",x"675c5a",x"5f5755",x"7d6c62",x"645b5c",x"6b6263",x"877871",x"81746e",x"92887f",x"92857f",x"93857c",x"91837a",x"92847b",x"93847d",x"90817a",x"8c817d",x"8b7e76",x"8a7d77",x"887b73",x"887b73",x"877a72",x"8c817d",x"585453",x"6f6765",x"86786d",x"6d6562",x"615a54",x"515153",x"585657",x"504e51",x"56514e",x"545351",x"555150",x"675e57",x"595554",x"535355",x"5a5a5c",x"535355",x"998c83",x"9a8c81",x"9c8e85",x"90837a",x"8f8079",x"93857c",x"907e72",x"8a796f",x"837366",x"95877e",x"90837b",x"948781",x"8d8077",x"94857e",x"90827f",x"827771",x"5c5656",x"5f5959",x"695f5d",x"5b5351"),
(x"5d5757",x"544f4c",x"5c5656",x"666263",x"60575a",x"605856",x"5b5756",x"5d5352",x"564c4a",x"605654",x"5c5859",x"6a605e",x"8d807a",x"928785",x"887d77",x"857a74",x"8f827c",x"867973",x"867970",x"8a7d75",x"92857f",x"938b88",x"92837c",x"8f8784",x"857b72",x"7d746f",x"877a74",x"887d77",x"525252",x"6f5e56",x"5e5a59",x"655c55",x"4c4a4f",x"675e5f",x"72685f",x"555354",x"555354",x"616163",x"66676c",x"585453",x"66615e",x"5d5e60",x"535152",x"504e51",x"9e9087",x"95877e",x"948278",x"9b8c85",x"988b83",x"97908a",x"94857e",x"938980",x"887a71",x"8c7e75",x"978c88",x"8c7b73",x"93867d",x"8e7f78",x"978a82",x"968b85",x"605758",x"5a5655",x"655d5b",x"565457"),
(x"665b57",x"635856",x"645955",x"5c5857",x"625a57",x"504c4d",x"5e5956",x"5b5653",x"696363",x"574d4c",x"695e5c",x"635957",x"978a82",x"8a7f79",x"958b89",x"9b918f",x"8d807a",x"90817a",x"8f827a",x"8c8482",x"978c88",x"8b7d74",x"887b73",x"8e8179",x"7b706c",x"817873",x"776a64",x"81746e",x"716966",x"555557",x"655d5a",x"635957",x"4d4c51",x"5b595a",x"626264",x"68635d",x"7b695d",x"5c5a5d",x"5a5a5c",x"715f55",x"5b595a",x"555658",x"665b55",x"6a635d",x"96887f",x"95847a",x"93827a",x"958880",x"91827b",x"8e8077",x"8d8078",x"90837d",x"90857f",x"887e75",x"8e817b",x"978881",x"958a84",x"91847e",x"9b8e86",x"978881",x"534d4d",x"585453",x"635b58",x"6a6562"),
(x"685d59",x"534f4e",x"595353",x"585252",x"5e5556",x"5b5253",x"55504d",x"5c4f49",x"5b5350",x"5b5351",x"5f5755",x"5c5250",x"908581",x"9d9088",x"9a938d",x"948985",x"89786e",x"91827b",x"90837d",x"7c7471",x"867970",x"887b75",x"827771",x"877c76",x"7e736d",x"887d77",x"877a72",x"7f726c",x"6d6d6f",x"64605d",x"676566",x"68686a",x"545456",x"635e5b",x"68615b",x"7d6f66",x"6b696c",x"6c6461",x"867970",x"565553",x"595758",x"5f5a57",x"5f5a57",x"7f6d63",x"9e9188",x"988b82",x"93867e",x"998e88",x"988b83",x"978881",x"877871",x"93847d",x"91827d",x"958a84",x"8b7d74",x"9c9289",x"958882",x"8e8179",x"988b83",x"978a81",x"5e5654",x"655d5b",x"625a58",x"554c4d"),
(x"655b5a",x"514947",x"6b6361",x"655b59",x"5e5556",x"605856",x"5b5351",x"726964",x"635e5b",x"635957",x"665d58",x"665c5b",x"968983",x"8b8178",x"93847f",x"a09790",x"998e88",x"94877e",x"82736c",x"928781",x"8c817b",x"8d827c",x"7f7470",x"7c6f69",x"7c716b",x"877a72",x"81746e",x"8e837d",x"696562",x"6c6b69",x"6f6d70",x"645e5e",x"575556",x"443a38",x"817069",x"5a5859",x"56555a",x"5f5e63",x"5e5e60",x"656162",x"6b6360",x"565658",x"5c5a5b",x"83726a",x"897e78",x"95867f",x"90817a",x"968980",x"998c84",x"9b918f",x"90827f",x"8f827a",x"8f817e",x"8b7e76",x"837874",x"877c76",x"988b83",x"93867e",x"9b8e86",x"91847c",x"504c4d",x"615956",x"685e5c",x"5e5654"),
(x"524c4c",x"504c4b",x"54504f",x"534f50",x"5e5654",x"5a5250",x"5f5959",x"59514e",x"796b62",x"625856",x"695f56",x"4f4b4c",x"92837c",x"8f827a",x"877c78",x"8e8a8b",x"938987",x"999089",x"938988",x"948a88",x"948781",x"7f7470",x"7f7470",x"867b75",x"92857d",x"8c817d",x"90857f",x"857872",x"6f6969",x"5f5a57",x"746c69",x"615f62",x"736862",x"646061",x"606060",x"696564",x"636164",x"5e5c61",x"615f60",x"616065",x"6e6159",x"646263",x"5e5c5d",x"7d6b61",x"9d9088",x"958b82",x"9b8e86",x"908279",x"897c74",x"8f8079",x"9a8c81",x"94877f",x"94867b",x"998c84",x"93857c",x"92847b",x"9b9289",x"9c938e",x"9c8f89",x"9a887e",x"555150",x"5f5755",x"5b5756",x"5c5656"),
(x"585453",x"555150",x"565253",x"5e5858",x"645a59",x"615b5b",x"544c49",x"786b65",x"565251",x"564e4c",x"645955",x"6a605f",x"8d7f7c",x"92857d",x"908b85",x"8b7e76",x"948781",x"958b89",x"7e7472",x"908684",x"8d8381",x"8f8583",x"857d7a",x"8d8582",x"91847e",x"90857f",x"91877e",x"998e8a",x"6e6d6b",x"6c6869",x"676566",x"81746e",x"817672",x"686765",x"5e5c5d",x"676568",x"69696b",x"686669",x"5f5e63",x"5c5b60",x"706a6a",x"605e61",x"616163",x"625e5d",x"92857f",x"948580",x"998a83",x"93867d",x"978d84",x"988b82",x"9c8e85",x"99877d",x"817674",x"8f8480",x"968b87",x"7e6f68",x"93877b",x"95847c",x"92887f",x"91847e",x"5a5454",x"6a6260",x"605a5a",x"595451")
);

end texture;

package body texture is


end texture;
