----------------------------------------------------------------------------------
-- Copyright 2020 Piotr Terczyński
--
-- Permission is hereby granted, free of charge, to any person
-- obtaining a copy of this software and associated           
-- documentation files (the "Software"), to deal in the       
-- Software without restriction, including without limitation 
-- the rights to use, copy, modify, merge, publish,           
-- distribute, sublicense, and/or sell copies of the Software,
-- and to permit persons to whom the Software is furnished to
-- do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice 
-- shall be included in all copies or substantial portions of
-- the Software.
--
-- 		THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF 
-- ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO 
-- THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR
-- PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS 
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR   
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR 
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE 
-- SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;
use work.definitions.all;

package model_presets is

constant light_norm_X_const : FLOAT16 := x"3565";
constant light_norm_Y_const : FLOAT16 := x"34c3";
constant light_norm_Z_const : FLOAT16 := x"3b24";

constant matrix_pp_const : TRANSFORM_MATRIX := (
(x"c30e",x"0000",x"c175",x"0000"),
(x"0000",x"4538",x"0000",x"c5be"),
(x"3918",x"0000",x"ba96",x"3e68"),
(x"40fe",x"0000",x"c274",x"491a")
);

subtype MM_ADDRESS is integer range 0 to 12171;
type MODEL_MEM is array (0 to 12171) of MOD_TRIANGLE;
constant AVAILABLE_TRIANGLES : integer := 12170;

constant model_const : MODEL_MEM :=(
empty_m_tri,
(x"b944",x"349b",x"3649",x"0000",x"8000",x"bc00",x"38ba",x"3b5b",x"b944",x"31a5",x"3649",x"0000",x"8000",x"bc00",x"38f2",x"3b5b",x"3a1c",x"349b",x"3649",x"0000",x"8000",x"bc00",x"38ba",x"39e5"),
(x"b944",x"345f",x"3745",x"0000",x"ba15",x"3932",x"3929",x"3b5b",x"b944",x"3468",x"3748",x"0000",x"ae16",x"3bf6",x"3933",x"3b5b",x"3a1c",x"345f",x"3745",x"8000",x"b970",x"39dd",x"3929",x"3a40"),
(x"b944",x"31a5",x"3727",x"0000",x"0000",x"3c00",x"38f2",x"3b5b",x"b944",x"3449",x"3727",x"0000",x"0000",x"3c00",x"3920",x"3b5b",x"3a1c",x"31a5",x"3727",x"0000",x"0000",x"3c00",x"38f2",x"39e5"),
(x"b944",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3b5b",x"b944",x"34b9",x"3649",x"0000",x"3c00",x"1a59",x"395b",x"3b5b",x"3a1c",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3a40"),
(x"b944",x"3468",x"3748",x"0000",x"ae16",x"3bf6",x"3933",x"3b5b",x"b944",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3b5b",x"3a1c",x"3468",x"3748",x"0000",x"a67a",x"3bff",x"3933",x"3a40"),
(x"b944",x"31a5",x"3649",x"0000",x"bc00",x"0000",x"395b",x"3b5b",x"b944",x"31a5",x"3727",x"0000",x"bc00",x"0000",x"3976",x"3b5b",x"3a1c",x"31a5",x"3649",x"0000",x"bc00",x"0000",x"395b",x"39e5"),
(x"b9bc",x"3d46",x"3653",x"0000",x"3c00",x"8000",x"2d82",x"3ab8",x"b9bc",x"3d46",x"b64b",x"0000",x"3c00",x"8000",x"1d3c",x"3ab8",x"3a8c",x"3d46",x"3653",x"0000",x"3c00",x"8000",x"2d82",x"3bfb"),
(x"b9c0",x"3d1e",x"3657",x"0000",x"bc00",x"0000",x"3b46",x"368f",x"3a88",x"3d1e",x"3657",x"0000",x"bc00",x"0000",x"3b46",x"37ad",x"b9c0",x"3d1e",x"b64b",x"0000",x"bc00",x"0000",x"3b90",x"368f"),
(x"3a8c",x"3d46",x"3653",x"0000",x"2631",x"3bff",x"399e",x"39c7",x"3a88",x"3d1e",x"3657",x"0000",x"2631",x"3bff",x"398a",x"39c7",x"b9bc",x"3d46",x"3653",x"0000",x"2631",x"3bff",x"399e",x"3b5b"),
(x"ba29",x"40b3",x"377b",x"b9af",x"39a0",x"8000",x"3728",x"3abe",x"ba29",x"40b3",x"b74a",x"ba61",x"38d2",x"0000",x"3726",x"3911",x"ba1e",x"40b8",x"376a",x"bb44",x"36ae",x"0000",x"3719",x"3abb"),
(x"ba22",x"4094",x"b74a",x"bba9",x"b498",x"8000",x"382d",x"39ad",x"ba27",x"4096",x"b74a",x"ba2e",x"b913",x"0000",x"3828",x"39ad",x"ba22",x"4094",x"3767",x"bb41",x"b6be",x"8000",x"382d",x"3ac9"),
(x"ba73",x"40a2",x"b74a",x"b892",x"ba90",x"0000",x"3775",x"3911",x"ba77",x"40a4",x"b74a",x"bb97",x"b50b",x"0000",x"3767",x"3911",x"ba73",x"40a2",x"3807",x"b8f8",x"ba45",x"0000",x"3775",x"3acc"),
(x"ba27",x"4096",x"b74a",x"ba2e",x"b913",x"0000",x"3828",x"39ad",x"ba30",x"4098",x"b74a",x"b91e",x"ba25",x"0000",x"3824",x"39ad",x"ba27",x"4096",x"3773",x"b9a4",x"b9ac",x"0000",x"3828",x"3acd"),
(x"ba12",x"408e",x"b751",x"0000",x"bc00",x"0000",x"3824",x"39ce",x"ba1f",x"408e",x"b74a",x"b1b5",x"bbdf",x"0000",x"3820",x"39cf",x"ba12",x"408e",x"3753",x"0000",x"bc00",x"0000",x"3824",x"3aca"),
(x"ba77",x"40a4",x"380c",x"bb97",x"b50c",x"0000",x"3767",x"3ad1",x"ba77",x"40a4",x"b74a",x"bb97",x"b50b",x"0000",x"3767",x"3911",x"ba77",x"40a6",x"380b",x"bbc1",x"33d8",x"8000",x"3759",x"3ad0"),
(x"ba30",x"4098",x"b74a",x"a918",x"bbfe",x"0000",x"37eb",x"3872",x"ba47",x"4098",x"b74a",x"adde",x"bbf7",x"0000",x"37e4",x"3872",x"ba30",x"4098",x"3785",x"a918",x"bbfe",x"0000",x"37eb",x"3967"),
(x"ba1f",x"408e",x"b74a",x"b1b5",x"bbdf",x"0000",x"3820",x"39cf",x"ba27",x"408f",x"b74a",x"b99f",x"b9b0",x"0000",x"381b",x"39cf",x"ba1f",x"408e",x"3769",x"b61a",x"bb65",x"8000",x"381f",x"3acd"),
(x"ba77",x"40a6",x"380b",x"bbc1",x"33d8",x"8000",x"3759",x"3ad0",x"ba77",x"40a6",x"b74a",x"baf6",x"37df",x"868d",x"3759",x"3911",x"ba72",x"40a7",x"3805",x"b7c0",x"3aff",x"0000",x"374b",x"3acc"),
(x"ba47",x"4098",x"b74a",x"adde",x"bbf7",x"0000",x"37e4",x"3872",x"ba4a",x"4099",x"b74a",x"baa8",x"b86e",x"0000",x"37dc",x"3872",x"ba47",x"4098",x"37b7",x"b2b5",x"bbd2",x"0000",x"37e4",x"396c"),
(x"ba27",x"408f",x"b74a",x"b99f",x"b9b0",x"0000",x"381b",x"39cf",x"ba29",x"4091",x"b74a",x"bbdb",x"31fa",x"0000",x"3817",x"39cf",x"ba27",x"408f",x"3777",x"bac3",x"b845",x"0000",x"381b",x"3ad0"),
(x"ba72",x"40a7",x"3805",x"b7c0",x"3aff",x"0000",x"374b",x"3acc",x"ba72",x"40a7",x"b74a",x"b671",x"3b52",x"868d",x"374b",x"3911",x"ba4d",x"40ab",x"37c7",x"b79e",x"3b08",x"0000",x"373b",x"3ac5"),
(x"ba4a",x"4099",x"b74a",x"baa8",x"b86e",x"0000",x"37dc",x"3872",x"ba4b",x"409a",x"b74a",x"bbfc",x"abd5",x"0000",x"37d3",x"3872",x"ba4a",x"4099",x"37bf",x"bb8d",x"b548",x"8000",x"37db",x"3970"),
(x"ba29",x"4091",x"3778",x"bbdb",x"31fb",x"0000",x"3817",x"3ad1",x"ba29",x"4091",x"b74a",x"bbdb",x"31fa",x"0000",x"3817",x"39cf",x"ba26",x"4092",x"3775",x"b8a6",x"3a82",x"0000",x"3813",x"3acf"),
(x"ba4d",x"40ab",x"37c7",x"b79e",x"3b08",x"0000",x"373b",x"3ac5",x"ba4d",x"40ab",x"b74a",x"b890",x"3a91",x"0000",x"373a",x"3911",x"ba29",x"40b3",x"377b",x"b9af",x"39a0",x"8000",x"3728",x"3abe"),
(x"ba4b",x"409a",x"37c0",x"bbfc",x"abd5",x"0000",x"37d3",x"3971",x"ba4b",x"409a",x"b74a",x"bbfc",x"abd5",x"0000",x"37d3",x"3872",x"ba4b",x"409b",x"37bd",x"bbb8",x"3431",x"8000",x"37cb",x"396e"),
(x"ba26",x"4092",x"3775",x"b8a6",x"3a82",x"0000",x"3813",x"3acf",x"ba26",x"4092",x"b74a",x"b5d6",x"3b72",x"8000",x"3813",x"39cf",x"ba21",x"4092",x"3766",x"b033",x"3bee",x"0000",x"380f",x"3aca"),
(x"ba4b",x"409b",x"37bd",x"bbb8",x"3431",x"8000",x"37cb",x"396e",x"ba4b",x"409b",x"b74a",x"bb4e",x"3681",x"068d",x"37cb",x"3872",x"ba49",x"409b",x"37ba",x"bad7",x"3825",x"0000",x"37c3",x"396c"),
(x"ba21",x"4092",x"b74a",x"bbe9",x"b0c1",x"0000",x"3831",x"39ad",x"ba22",x"4094",x"b74a",x"bba9",x"b498",x"8000",x"382d",x"39ad",x"ba21",x"4092",x"3766",x"bbe9",x"b0c2",x"0000",x"3832",x"3ac9"),
(x"ba49",x"409b",x"b74a",x"b863",x"bab0",x"0000",x"378a",x"3911",x"ba73",x"40a2",x"b74a",x"b892",x"ba90",x"0000",x"3775",x"3911",x"ba49",x"409b",x"37ba",x"b863",x"bab0",x"0000",x"378a",x"3ac3"),
(x"ba12",x"3d46",x"b578",x"b9e8",x"3889",x"35d4",x"2dfc",x"2140",x"ba05",x"3d46",x"b544",x"ba14",x"38d9",x"337c",x"2dd6",x"20e8",x"ba12",x"3d41",x"b55a",x"b9cc",x"38ee",x"34e9",x"2de7",x"218f"),
(x"ba12",x"3d41",x"b55a",x"b9cc",x"38ee",x"34e9",x"2de7",x"218f",x"ba05",x"3d46",x"b544",x"ba14",x"38d9",x"337c",x"2dd6",x"20e8",x"ba12",x"3d3b",x"b522",x"ba50",x"38e8",x"2604",x"2dbf",x"21f1"),
(x"ba12",x"3d3b",x"b522",x"ba50",x"38e8",x"2604",x"2dbf",x"21f1",x"ba02",x"3d46",x"b515",x"ba7c",x"38ae",x"1c81",x"2db6",x"20d0",x"ba12",x"3d3a",x"b07b",x"ba7d",x"38ad",x"9e59",x"2b8b",x"21f1"),
(x"ba12",x"3d46",x"af74",x"ba37",x"3832",x"b58f",x"2b03",x"211f",x"ba12",x"3d3f",x"b00e",x"ba6d",x"3864",x"b364",x"2b40",x"219c",x"ba09",x"3d45",x"b010",x"ba60",x"3855",x"b446",x"2b42",x"20ee"),
(x"ba12",x"3d3a",x"b07b",x"ba7d",x"38ad",x"9e59",x"2b8b",x"21f1",x"ba03",x"3d45",x"b075",x"baa1",x"3878",x"a594",x"2b88",x"20ca",x"ba12",x"3d3f",x"b00e",x"ba6d",x"3864",x"b364",x"2b40",x"219c"),
(x"b9dc",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"b9dc",x"3d46",x"aca4",x"9d38",x"3c00",x"8cea",x"2392",x"2238",x"ba02",x"3d46",x"b515",x"9f10",x"3c00",x"1018",x"2b3f",x"23cc"),
(x"b9dc",x"3d46",x"aca4",x"9d38",x"3c00",x"8cea",x"2392",x"2238",x"ba12",x"3d46",x"af74",x"1f79",x"3c00",x"9c81",x"25b4",x"243e",x"ba09",x"3d45",x"b010",x"20d0",x"3bff",x"a081",x"262a",x"240d"),
(x"ba12",x"4070",x"af8a",x"0000",x"bc00",x"0000",x"2d06",x"2458",x"b9dc",x"4070",x"aca4",x"0e8d",x"bc00",x"8000",x"2c87",x"257b",x"ba09",x"4070",x"b010",x"0000",x"bc00",x"0000",x"2d20",x"248a"),
(x"b9dc",x"4070",x"b64e",x"11bc",x"bc00",x"8000",x"3005",x"257b",x"ba02",x"4070",x"b515",x"128d",x"bc00",x"868d",x"2f35",x"24b1",x"b9dc",x"4070",x"aca4",x"0e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"b9f4",x"4047",x"b504",x"ba04",x"8000",x"b945",x"31d7",x"35aa",x"b9f4",x"3d94",x"b504",x"ba04",x"8000",x"b945",x"31d8",x"3356",x"b9dc",x"404e",x"b53c",x"ba04",x"8000",x"b945",x"31be",x"35b4"),
(x"b9f4",x"3d94",x"b504",x"ba28",x"b91a",x"0000",x"31e3",x"290c",x"b9f4",x"3d94",x"b0a7",x"ba28",x"b91a",x"0000",x"30f8",x"290c",x"b9dc",x"3d85",x"b53c",x"ba28",x"b91a",x"0000",x"31f6",x"2973"),
(x"b9dc",x"3d85",x"b032",x"ba1b",x"0000",x"392a",x"317f",x"3342",x"b9f4",x"3d94",x"b0a7",x"ba1b",x"0000",x"392a",x"3165",x"3356",x"b9dc",x"404e",x"b032",x"ba1b",x"0000",x"392a",x"317f",x"35b4"),
(x"ba12",x"4076",x"b07b",x"ba77",x"b8b5",x"9fc8",x"310a",x"2c8f",x"ba12",x"4073",x"b00e",x"ba59",x"b87c",x"b388",x"30f7",x"2c99",x"ba03",x"4070",x"b075",x"ba96",x"b888",x"a5cf",x"3109",x"2cb3"),
(x"ba12",x"4073",x"b00e",x"ba59",x"b87c",x"b388",x"30f7",x"2c99",x"ba12",x"4070",x"af8a",x"ba0f",x"b848",x"b5fa",x"30ea",x"2ca7",x"ba09",x"4070",x"b010",x"ba44",x"b877",x"b45c",x"30f8",x"2cae"),
(x"b9f4",x"4047",x"b0a7",x"bc00",x"0000",x"0000",x"301e",x"3185",x"b9f4",x"3d94",x"b0a7",x"bc00",x"0000",x"0000",x"301e",x"2c2f",x"b9f4",x"4047",x"b504",x"bc00",x"0000",x"0000",x"2ea8",x"3185"),
(x"b9dc",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"31dc",x"b9dc",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"2b18",x"b9dc",x"404e",x"b032",x"bc00",x"0000",x"0000",x"302e",x"318f"),
(x"ba12",x"4076",x"b522",x"ba50",x"b8e8",x"25a1",x"3207",x"2c8f",x"ba12",x"4076",x"b07b",x"ba77",x"b8b5",x"9fc8",x"310a",x"2c8f",x"ba02",x"4070",x"b515",x"ba76",x"b8b6",x"1ac2",x"3203",x"2cb3"),
(x"b9dc",x"3d85",x"b032",x"bc00",x"0000",x"0000",x"302e",x"2c1c",x"b9dc",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"2b18",x"b9dc",x"3d85",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"2c1c"),
(x"b9dc",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2def",x"31dc",x"b9dc",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"31dc",x"b9dc",x"404e",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"318f"),
(x"b9dc",x"3d85",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"2c1c",x"b9dc",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2def",x"2b18",x"b9dc",x"404e",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"318f"),
(x"ba12",x"4073",x"b55a",x"b9cc",x"b8ee",x"34e9",x"321b",x"2c9b",x"ba12",x"4076",x"b522",x"ba50",x"b8e8",x"25a1",x"3207",x"2c8f",x"ba05",x"4070",x"b544",x"ba14",x"b8d9",x"337c",x"3212",x"2cb0"),
(x"ba05",x"4070",x"b544",x"ba14",x"b8d9",x"337c",x"3212",x"2cb0",x"ba12",x"4070",x"b578",x"b9e8",x"b889",x"35d4",x"3226",x"2ca5",x"ba12",x"4073",x"b55a",x"b9cc",x"b8ee",x"34e9",x"321b",x"2c9b"),
(x"b9dc",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"3350",x"b9dc",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"2cf5",x"ba12",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"3350"),
(x"b9dc",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"ba05",x"3d46",x"b544",x"0000",x"3c00",x"8000",x"2b7e",x"23f3",x"ba12",x"3d46",x"b578",x"0000",x"3c00",x"8000",x"2bc6",x"243e"),
(x"b9dc",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"ba07",x"3d83",x"aca4",x"0000",x"8000",x"bc00",x"312d",x"2d9a",x"ba12",x"3d7a",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2d80"),
(x"b9dc",x"404e",x"b032",x"ba28",x"391a",x"0000",x"30e4",x"297b",x"b9f4",x"4047",x"b0a7",x"ba28",x"391a",x"0000",x"30f8",x"29e2",x"b9dc",x"404e",x"b53c",x"ba28",x"391a",x"0000",x"31f6",x"297b"),
(x"ba12",x"4070",x"b578",x"0e8d",x"bc00",x"868d",x"2f78",x"2458",x"ba05",x"4070",x"b544",x"0cea",x"bc00",x"8a8d",x"2f54",x"249e",x"b9dc",x"4070",x"b64e",x"11bc",x"bc00",x"8000",x"3005",x"257b"),
(x"ba12",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"31e6",x"ba12",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"2af0",x"ba12",x"3cb5",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"31f0"),
(x"ba07",x"3d83",x"aca4",x"b9a1",x"3488",x"b935",x"31de",x"3350",x"ba12",x"3d84",x"ac3b",x"b9ce",x"340f",x"b91d",x"31ea",x"3351",x"ba12",x"3d7a",x"aca4",x"b950",x"3666",x"b90d",x"31e3",x"3342"),
(x"b9dc",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"b9dc",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"b9ff",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe"),
(x"b9dc",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"ba12",x"4057",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"330c",x"ba02",x"404f",x"aca4",x"0000",x"8000",x"bc00",x"312a",x"32f6"),
(x"ba12",x"3d92",x"abd9",x"ba32",x"17c8",x"b90f",x"31ef",x"3364",x"ba12",x"3d84",x"ac3b",x"b9ce",x"340f",x"b91d",x"31ea",x"3351",x"b9ff",x"3d91",x"aca4",x"ba3a",x"1e3f",x"b904",x"31db",x"3363"),
(x"ba12",x"404b",x"abe1",x"ba2a",x"96f6",x"b918",x"31ef",x"35b8",x"ba12",x"3d92",x"abd9",x"ba32",x"17c8",x"b90f",x"31ef",x"3364",x"b9ff",x"404b",x"aca4",x"ba32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"ba02",x"404f",x"aca4",x"b9d3",x"b46b",x"b903",x"31dc",x"35bd",x"ba12",x"404f",x"ac0f",x"b9ea",x"b3b0",x"b908",x"31ed",x"35bd",x"b9ff",x"404b",x"aca4",x"ba32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"ba12",x"4057",x"aca4",x"b9ad",x"b59c",x"b8e3",x"31e3",x"35c9",x"ba12",x"404f",x"ac0f",x"b9ea",x"b3b0",x"b908",x"31ed",x"35bd",x"ba02",x"404f",x"aca4",x"b9d3",x"b46b",x"b903",x"31dc",x"35bd"),
(x"ba07",x"3d45",x"3551",x"ba36",x"38b3",x"b345",x"2477",x"1cd0",x"ba12",x"3d46",x"3587",x"ba16",x"3888",x"b50c",x"23b9",x"1d50",x"ba12",x"3d3e",x"3554",x"ba2c",x"38a8",x"b41a",x"246e",x"1e40"),
(x"ba12",x"3d3e",x"3554",x"ba2c",x"38a8",x"b41a",x"246e",x"1e40",x"ba12",x"3d3a",x"3523",x"ba4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"ba07",x"3d45",x"3551",x"ba36",x"38b3",x"b345",x"2477",x"1cd0"),
(x"ba12",x"3d3a",x"3523",x"ba4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"ba12",x"3d3a",x"3099",x"ba5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"ba01",x"3d45",x"351f",x"ba5d",x"38d8",x"9f93",x"2503",x"1c77"),
(x"ba12",x"3d3e",x"3026",x"ba1b",x"38d7",x"3338",x"2aab",x"1e54",x"ba12",x"3d46",x"2f74",x"b9ff",x"3898",x"3541",x"2af9",x"1d4d",x"ba06",x"3d45",x"302e",x"ba14",x"38b9",x"3455",x"2aa5",x"1cb4"),
(x"ba12",x"3d3a",x"3099",x"ba5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"ba12",x"3d3e",x"3026",x"ba1b",x"38d7",x"3338",x"2aab",x"1e54",x"ba01",x"3d45",x"307d",x"ba66",x"38cb",x"2460",x"2a6e",x"1c77"),
(x"b9dc",x"3d46",x"364e",x"9e0a",x"3c00",x"91bc",x"2392",x"257f",x"ba01",x"3d45",x"351f",x"a259",x"3bff",x"068d",x"2705",x"2646",x"b9dc",x"3d46",x"2ce6",x"a067",x"3c00",x"1018",x"2c69",x"257f"),
(x"ba12",x"3d46",x"2f74",x"1ea7",x"3c00",x"1c67",x"2bf4",x"26a1",x"b9dc",x"3d46",x"2ce6",x"a067",x"3c00",x"1018",x"2c69",x"257f",x"ba06",x"3d45",x"302e",x"2025",x"3bff",x"2025",x"2ba5",x"265f"),
(x"b9dc",x"4070",x"2ce6",x"0e8d",x"bc00",x"8000",x"2c74",x"27d3",x"ba12",x"4070",x"2f82",x"0000",x"bc00",x"0000",x"2c02",x"26b0",x"ba09",x"4070",x"300c",x"0000",x"bc00",x"0000",x"2bd2",x"26e2"),
(x"b9dc",x"4070",x"364e",x"11bc",x"bc00",x"8000",x"23e8",x"27d3",x"b9dc",x"4070",x"2ce6",x"0e8d",x"bc00",x"8000",x"2c74",x"27d3",x"ba02",x"4070",x"3524",x"128d",x"bc00",x"068d",x"2720",x"2709"),
(x"b9dc",x"3d85",x"354b",x"ba04",x"0000",x"3945",x"31ba",x"3342",x"b9f4",x"3d94",x"3513",x"ba04",x"0000",x"3945",x"31a1",x"3356",x"b9dc",x"404e",x"354b",x"ba04",x"0000",x"3945",x"31ba",x"35b4"),
(x"b9dc",x"3d85",x"3069",x"ba28",x"b91a",x"0000",x"31f8",x"2b0f",x"b9f4",x"3d94",x"30dd",x"ba28",x"b91a",x"0000",x"31e4",x"2aa8",x"b9dc",x"3d85",x"354b",x"ba28",x"b91a",x"0000",x"30ea",x"2b0f"),
(x"b9dc",x"3d85",x"3069",x"ba15",x"8000",x"b931",x"3183",x"3342",x"b9dc",x"404e",x"3069",x"ba15",x"8000",x"b931",x"3183",x"35b4",x"b9f4",x"3d94",x"30dd",x"ba15",x"8000",x"b931",x"319d",x"3356"),
(x"ba12",x"4076",x"3076",x"ba76",x"b8b6",x"1fc8",x"2a73",x"1f14",x"ba03",x"4070",x"3071",x"ba97",x"b888",x"25b5",x"2a77",x"20ad",x"ba12",x"4073",x"300a",x"ba59",x"b87c",x"3388",x"2abf",x"1fbf"),
(x"ba12",x"4070",x"2f82",x"ba0f",x"b848",x"35fa",x"2af4",x"2050",x"ba12",x"4073",x"300a",x"ba59",x"b87c",x"3388",x"2abf",x"1fbf",x"ba09",x"4070",x"300c",x"ba44",x"b877",x"345b",x"2abd",x"2088"),
(x"b9f4",x"4047",x"30dd",x"bc00",x"0000",x"0000",x"272f",x"317f",x"b9f4",x"4047",x"3513",x"bc00",x"0000",x"0000",x"2aa7",x"317f",x"b9f4",x"3d94",x"30dd",x"bc00",x"0000",x"0000",x"272f",x"2c38"),
(x"b9dc",x"3d85",x"3069",x"bc00",x"0000",x"0000",x"26a2",x"2c24",x"b9dc",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"2b2a",x"b9dc",x"404e",x"3069",x"bc00",x"0000",x"0000",x"26a2",x"318a"),
(x"ba12",x"4076",x"3532",x"ba50",x"b8e8",x"a587",x"24d1",x"1f14",x"ba02",x"4070",x"3524",x"ba76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"ba12",x"4076",x"3076",x"ba76",x"b8b6",x"1fc8",x"2a73",x"1f14"),
(x"b9dc",x"3d85",x"3069",x"bc00",x"0000",x"0000",x"26a2",x"2c24",x"b9dc",x"3d85",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"2c24",x"b9dc",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"2b2a"),
(x"b9dc",x"404e",x"3069",x"bc00",x"0000",x"0000",x"26a2",x"318a",x"b9dc",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"31d6",x"b9dc",x"404e",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"318a"),
(x"b9dc",x"3d85",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"2c24",x"b9dc",x"404e",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"318a",x"b9dc",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"2c00",x"2b2a"),
(x"ba12",x"4073",x"3569",x"b9cc",x"b8ee",x"b4e9",x"2433",x"1fda",x"ba05",x"4070",x"3553",x"ba14",x"b8d9",x"b37c",x"2475",x"2093",x"ba12",x"4076",x"3532",x"ba50",x"b8e8",x"a587",x"24d1",x"1f14"),
(x"ba12",x"4070",x"3587",x"b9e8",x"b889",x"b5d4",x"23b9",x"203c",x"ba05",x"4070",x"3553",x"ba14",x"b8d9",x"b37c",x"2475",x"2093",x"ba12",x"4073",x"3569",x"b9cc",x"b8ee",x"b4e9",x"2433",x"1fda"),
(x"ba12",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"315d",x"2cf5",x"b9dc",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"3138",x"2cf5",x"ba12",x"4070",x"364e",x"0000",x"8000",x"bc00",x"315d",x"3350"),
(x"ba12",x"3d46",x"3587",x"204d",x"3c00",x"9cb5",x"25e8",x"26a2",x"ba07",x"3d45",x"3551",x"14ea",x"3c00",x"9dd6",x"267b",x"2668",x"b9dc",x"3d46",x"364e",x"9e0a",x"3c00",x"91bc",x"2392",x"257f"),
(x"ba12",x"3d7a",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2d50",x"ba08",x"3d84",x"2ce6",x"0000",x"0000",x"3c00",x"3169",x"2d69",x"b9dc",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"b9dc",x"404e",x"3069",x"ba28",x"391a",x"0000",x"31f8",x"2b16",x"b9dc",x"404e",x"354b",x"ba28",x"391a",x"0000",x"30ea",x"2b16",x"b9f4",x"4047",x"30dd",x"ba28",x"391a",x"0000",x"31e4",x"2b7e"),
(x"b9dc",x"4070",x"364e",x"11bc",x"bc00",x"8000",x"23e8",x"27d3",x"ba05",x"4070",x"3553",x"10ea",x"bc00",x"068d",x"26a2",x"26f5",x"ba12",x"4070",x"3587",x"0e8d",x"bc00",x"0a8d",x"2613",x"26b0"),
(x"ba12",x"404f",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"355a",x"ba12",x"4057",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3564",x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583"),
(x"ba12",x"3d85",x"2c89",x"b9d0",x"342d",x"3915",x"31f9",x"3351",x"ba08",x"3d84",x"2ce6",x"b9a5",x"3468",x"3938",x"3203",x"3350",x"ba12",x"3d7a",x"2ce6",x"b96d",x"35b1",x"3924",x"31ff",x"3342"),
(x"ba01",x"3d90",x"2ce6",x"0000",x"0000",x"3c00",x"316e",x"2d8c",x"b9ff",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1",x"b9dc",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"ba12",x"4056",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"32f1",x"b9dc",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"ba03",x"404f",x"2ce6",x"0000",x"0000",x"3c00",x"316c",x"32dd"),
(x"ba08",x"3d84",x"2ce6",x"b9a5",x"3468",x"3938",x"3203",x"3350",x"ba12",x"3d85",x"2c89",x"b9d0",x"342d",x"3915",x"31f9",x"3351",x"ba01",x"3d90",x"2ce6",x"ba49",x"1ec2",x"38f2",x"3206",x"3362"),
(x"ba01",x"3d90",x"2ce6",x"ba49",x"1ec2",x"38f2",x"3206",x"3362",x"ba12",x"3d92",x"2c35",x"ba20",x"184d",x"3924",x"31f3",x"3363",x"b9ff",x"404a",x"2ce6",x"ba20",x"935f",x"3925",x"3206",x"35b6"),
(x"b9ff",x"404a",x"2ce6",x"ba20",x"935f",x"3925",x"3206",x"35b6",x"ba12",x"404b",x"2c40",x"b9f4",x"9af6",x"3957",x"31f3",x"35b7",x"ba03",x"404f",x"2ce6",x"b9e5",x"b3cc",x"390b",x"3204",x"35bc"),
(x"ba12",x"404e",x"2c57",x"b9db",x"b485",x"38f4",x"31f4",x"35bc",x"ba12",x"4056",x"2ce6",x"b9b2",x"b5ad",x"38d8",x"31fe",x"35c7",x"ba03",x"404f",x"2ce6",x"b9e5",x"b3cc",x"390b",x"3204",x"35bc"),
(x"ba12",x"3507",x"b578",x"b9e8",x"3889",x"35d4",x"3227",x"2c75",x"ba05",x"3507",x"b544",x"ba14",x"38d9",x"337c",x"3214",x"2c6a",x"ba12",x"34f4",x"b55a",x"b9cc",x"38ee",x"34e9",x"321c",x"2c7f"),
(x"ba12",x"34f4",x"b55a",x"b9cc",x"38ee",x"34e9",x"321c",x"2c7f",x"ba05",x"3507",x"b544",x"ba14",x"38d9",x"337c",x"3214",x"2c6a",x"ba12",x"34dc",x"b522",x"ba50",x"38e8",x"2604",x"3209",x"2c8b"),
(x"ba12",x"34dc",x"b522",x"ba50",x"38e8",x"2604",x"3209",x"2c8b",x"ba02",x"3507",x"b515",x"ba7c",x"38ae",x"1c81",x"3204",x"2c67",x"ba12",x"34d8",x"b07b",x"ba7d",x"38ad",x"9e59",x"310c",x"2c8b"),
(x"ba12",x"3507",x"af74",x"ba37",x"3832",x"b58f",x"30ea",x"2c71",x"ba12",x"34eb",x"b00e",x"ba6d",x"3864",x"b364",x"30f9",x"2c80",x"ba09",x"3506",x"b010",x"ba5f",x"3855",x"b446",x"30f9",x"2c6a"),
(x"ba12",x"34d8",x"b07b",x"ba7d",x"38ad",x"9e59",x"310c",x"2c8b",x"ba03",x"3506",x"b075",x"baa1",x"3878",x"a594",x"310b",x"2c66",x"ba12",x"34eb",x"b00e",x"ba6d",x"3864",x"b364",x"30f9",x"2c80"),
(x"b9dc",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"b9dc",x"3507",x"aca4",x"9d38",x"3c00",x"8cea",x"2c87",x"224e",x"ba02",x"3507",x"b515",x"9f10",x"3c00",x"1018",x"2f35",x"23e3"),
(x"b9dc",x"3507",x"aca4",x"9d38",x"3c00",x"8cea",x"2c87",x"224e",x"ba12",x"3507",x"af74",x"1f79",x"3c00",x"9c81",x"2d02",x"244a",x"ba09",x"3506",x"b010",x"20d0",x"3bff",x"a081",x"2d20",x"2418"),
(x"ba12",x"3cac",x"af8a",x"0000",x"bc00",x"0000",x"25c3",x"244d",x"b9dc",x"3cac",x"aca4",x"0e8d",x"bc00",x"8000",x"2392",x"2570",x"ba09",x"3cac",x"b010",x"0000",x"bc00",x"0000",x"262a",x"247f"),
(x"b9dc",x"3cac",x"b64e",x"11bc",x"bc00",x"8000",x"2c74",x"2570",x"ba02",x"3cac",x"b515",x"128d",x"bc00",x"868d",x"2b3f",x"24a6",x"b9dc",x"3cac",x"aca4",x"0e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"b9dc",x"3c69",x"b53c",x"ba04",x"8000",x"b945",x"3127",x"35a2",x"b9f4",x"3c5a",x"b504",x"ba04",x"8000",x"b945",x"3140",x"3598",x"b9dc",x"35ff",x"b53c",x"ba04",x"8000",x"b945",x"3127",x"335c"),
(x"b9f4",x"3638",x"b504",x"ba0b",x"b93d",x"0000",x"31e9",x"2bf4",x"b9f4",x"3638",x"b0a7",x"ba0b",x"b93d",x"0000",x"30fe",x"2bf4",x"b9dc",x"35ff",x"b53c",x"ba0b",x"b93d",x"0000",x"31fc",x"2c2c"),
(x"b9f4",x"3638",x"b0a7",x"ba1b",x"0000",x"392a",x"30ec",x"336f",x"b9f4",x"3c5a",x"b0a7",x"ba1b",x"0000",x"392a",x"30ec",x"3598",x"b9dc",x"35ff",x"b032",x"ba1b",x"0000",x"392a",x"3106",x"335c"),
(x"ba12",x"3cb8",x"b07b",x"ba77",x"b8b5",x"9fc8",x"24df",x"20ca",x"ba12",x"3cb3",x"b00e",x"ba59",x"b87c",x"b388",x"2447",x"2120",x"ba03",x"3cac",x"b075",x"ba96",x"b888",x"a5cf",x"24d8",x"21ed"),
(x"ba12",x"3cb3",x"b00e",x"ba59",x"b87c",x"b388",x"2447",x"2120",x"ba12",x"3cac",x"af8a",x"ba0f",x"b848",x"b5fa",x"23b9",x"2190",x"ba09",x"3cac",x"b010",x"ba44",x"b877",x"b45c",x"244b",x"21c8"),
(x"b9f4",x"3c5a",x"b0a7",x"bc00",x"0000",x"0000",x"2ac8",x"3545",x"b9f4",x"3638",x"b0a7",x"bc00",x"0000",x"0000",x"2ac8",x"330c",x"b9f4",x"3c5a",x"b504",x"bc00",x"0000",x"0000",x"26b9",x"3545"),
(x"b9dc",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"3575",x"b9dc",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"32d0",x"b9dc",x"3c69",x"b032",x"bc00",x"0000",x"0000",x"3036",x"354d"),
(x"ba12",x"3cb7",x"b522",x"ba50",x"b8e8",x"25a8",x"2a63",x"20cc",x"ba12",x"3cb8",x"b07b",x"ba77",x"b8b5",x"9fc8",x"24df",x"20ca",x"ba02",x"3cac",x"b515",x"ba76",x"b8b6",x"1ac2",x"2a51",x"21ed"),
(x"b9dc",x"35ff",x"b032",x"bc00",x"0000",x"0000",x"3036",x"331b",x"b9dc",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"32d0",x"b9dc",x"35ff",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"331b"),
(x"b9dc",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2ddb",x"3575",x"b9dc",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"3575",x"b9dc",x"3c69",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"354d"),
(x"b9dc",x"35ff",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"331b",x"b9dc",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2ddb",x"32d0",x"b9dc",x"3c69",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"354d"),
(x"ba12",x"3cb1",x"b55a",x"b9cc",x"b8ee",x"34e9",x"2ab1",x"212f",x"ba12",x"3cb7",x"b522",x"ba50",x"b8e8",x"25a8",x"2a63",x"20cc",x"ba05",x"3cac",x"b544",x"ba14",x"b8d9",x"337c",x"2a90",x"21d6"),
(x"ba05",x"3cac",x"b544",x"ba14",x"b8d9",x"337c",x"2a90",x"21d6",x"ba12",x"3cac",x"b578",x"b9e8",x"b889",x"35d4",x"2add",x"217f",x"ba12",x"3cb1",x"b55a",x"b9cc",x"b8ee",x"34e9",x"2ab1",x"212f"),
(x"b9dc",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"333a",x"b9dc",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"2d4a",x"ba12",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"333a"),
(x"b9dc",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"ba05",x"3507",x"b544",x"0000",x"3c00",x"8000",x"2f54",x"2404",x"ba12",x"3507",x"b578",x"0000",x"3c00",x"8000",x"2f78",x"244a"),
(x"b9dc",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a",x"ba07",x"35fb",x"aca4",x"0000",x"8000",x"bc00",x"31fc",x"2dee",x"ba12",x"35d5",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2dd4"),
(x"b9dc",x"3c69",x"b032",x"ba28",x"391a",x"0000",x"30ea",x"2a0f",x"b9f4",x"3c5a",x"b0a7",x"ba28",x"391a",x"0000",x"30fe",x"2a76",x"b9dc",x"3c69",x"b53c",x"ba28",x"391a",x"0000",x"31fc",x"2a0f"),
(x"ba12",x"3cac",x"b578",x"0e8d",x"bc00",x"8a8d",x"2bc6",x"244d",x"ba05",x"3cac",x"b544",x"10ea",x"bc00",x"868d",x"2b7e",x"2492",x"b9dc",x"3cac",x"b64e",x"11bc",x"bc00",x"8000",x"2c74",x"2570"),
(x"ba07",x"35fb",x"aca4",x"b9a1",x"3488",x"b935",x"320d",x"3350",x"ba12",x"35fe",x"ac3b",x"b9ce",x"340f",x"b91d",x"3219",x"3351",x"ba12",x"35d5",x"aca4",x"b950",x"3666",x"b90d",x"3212",x"3342"),
(x"b9dc",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"b9ff",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"b9dc",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"b9dc",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"ba12",x"3c7a",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"32f6",x"ba02",x"3c6a",x"aca4",x"0000",x"8000",x"bc00",x"31f9",x"32e0"),
(x"ba12",x"3635",x"abd9",x"ba32",x"1818",x"b90f",x"321e",x"3364",x"ba12",x"35fe",x"ac3b",x"b9ce",x"340f",x"b91d",x"3219",x"3351",x"b9ff",x"3631",x"aca4",x"ba3a",x"1e8d",x"b905",x"320a",x"3363"),
(x"ba12",x"3c61",x"abe1",x"ba2a",x"97c8",x"b918",x"321e",x"3597",x"ba12",x"3635",x"abd9",x"ba32",x"1818",x"b90f",x"321e",x"3364",x"b9ff",x"3c61",x"aca4",x"ba32",x"9624",x"b90f",x"320a",x"3597"),
(x"ba02",x"3c6a",x"aca4",x"b9d3",x"b46b",x"b903",x"320b",x"359d",x"ba12",x"3c6a",x"ac0f",x"b9ea",x"b3b0",x"b908",x"321c",x"359d",x"b9ff",x"3c61",x"aca4",x"ba32",x"9624",x"b90f",x"320a",x"3597"),
(x"ba12",x"3c7a",x"aca4",x"b9ad",x"b59c",x"b8e3",x"3212",x"35a9",x"ba12",x"3c6a",x"ac0f",x"b9ea",x"b3b0",x"b908",x"321c",x"359d",x"ba02",x"3c6a",x"aca4",x"b9d3",x"b46b",x"b903",x"320b",x"359d"),
(x"ba07",x"3505",x"3551",x"ba36",x"38b3",x"b345",x"2b55",x"1cd0",x"ba12",x"3507",x"3587",x"ba16",x"3888",x"b50c",x"2b07",x"1d50",x"ba12",x"34ea",x"3554",x"ba2c",x"38a8",x"b41a",x"2b50",x"1e40"),
(x"ba12",x"34ea",x"3554",x"ba2c",x"38a8",x"b41a",x"2b50",x"1e40",x"ba12",x"34db",x"3523",x"ba4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"ba07",x"3505",x"3551",x"ba36",x"38b3",x"b345",x"2b55",x"1cd0"),
(x"ba12",x"34db",x"3523",x"ba4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"ba12",x"34d8",x"3099",x"ba5b",x"38da",x"1d38",x"2dba",x"1ed9",x"ba01",x"3506",x"351f",x"ba5d",x"38d8",x"9f93",x"2b9a",x"1c77"),
(x"ba12",x"34e8",x"3026",x"ba1b",x"38d7",x"3338",x"2de2",x"1e54",x"ba12",x"3507",x"2f74",x"b9ff",x"3898",x"3541",x"2e09",x"1d4d",x"ba06",x"3506",x"302e",x"ba14",x"38b9",x"3455",x"2ddf",x"1cb4"),
(x"ba12",x"34d8",x"3099",x"ba5b",x"38da",x"1d38",x"2dba",x"1ed9",x"ba12",x"34e8",x"3026",x"ba1b",x"38d7",x"3338",x"2de2",x"1e54",x"ba01",x"3506",x"307d",x"ba66",x"38cb",x"2460",x"2dc4",x"1c77"),
(x"b9dc",x"3507",x"364e",x"9e0a",x"3c00",x"91bc",x"2c87",x"258a",x"ba01",x"3506",x"351f",x"a259",x"3bff",x"868d",x"2d56",x"2651",x"b9dc",x"3507",x"2ce6",x"a067",x"3c00",x"1018",x"2fff",x"258a"),
(x"ba12",x"3507",x"2f74",x"1ea7",x"3c00",x"1c67",x"2f8f",x"26ad",x"b9dc",x"3507",x"2ce6",x"a067",x"3c00",x"1018",x"2fff",x"258a",x"ba06",x"3506",x"302e",x"2032",x"3bff",x"2025",x"2f68",x"266a"),
(x"b9dc",x"3cac",x"2ce6",x"0e8d",x"bc00",x"8000",x"2fff",x"27de",x"ba12",x"3cac",x"2f82",x"0000",x"bc00",x"0000",x"2f8d",x"26bb",x"ba09",x"3cac",x"300c",x"0000",x"bc00",x"0000",x"2f73",x"26ed"),
(x"b9dc",x"3cac",x"364e",x"11bc",x"bc00",x"8000",x"2c87",x"27de",x"b9dc",x"3cac",x"2ce6",x"0e8d",x"bc00",x"8000",x"2fff",x"27de",x"ba02",x"3cac",x"3524",x"128d",x"bc00",x"068d",x"2d52",x"2714"),
(x"b9dc",x"3c69",x"354b",x"ba04",x"0000",x"3945",x"315d",x"35a1",x"b9dc",x"3600",x"354b",x"ba04",x"0000",x"3945",x"315d",x"335c",x"b9f4",x"3c5a",x"3513",x"ba04",x"0000",x"3945",x"3144",x"3597"),
(x"b9dc",x"3600",x"3069",x"ba0f",x"b938",x"0000",x"31f8",x"2c62",x"b9f4",x"3639",x"30dd",x"ba0f",x"b938",x"0000",x"31e4",x"2c30",x"b9dc",x"3600",x"354b",x"ba0f",x"b938",x"0000",x"30ea",x"2c62"),
(x"b9dc",x"3c69",x"3069",x"ba15",x"8000",x"b931",x"3109",x"35a1",x"b9f4",x"3c5a",x"30dd",x"ba15",x"8000",x"b931",x"3123",x"3597",x"b9dc",x"3600",x"3069",x"ba15",x"8000",x"b931",x"3109",x"335c"),
(x"ba12",x"3cb8",x"3076",x"ba76",x"b8b6",x"1fc8",x"2dc6",x"1f14",x"ba03",x"3cac",x"3071",x"ba97",x"b888",x"25b5",x"2dc8",x"20ad",x"ba12",x"3cb3",x"300a",x"ba59",x"b87c",x"3388",x"2dec",x"1fbf"),
(x"ba12",x"3cac",x"2f82",x"ba0f",x"b848",x"35fa",x"2e07",x"2050",x"ba12",x"3cb3",x"300a",x"ba59",x"b87c",x"3388",x"2dec",x"1fbf",x"ba09",x"3cac",x"300c",x"ba44",x"b877",x"345c",x"2deb",x"2088"),
(x"b9f4",x"3c5a",x"30dd",x"bc00",x"0000",x"0000",x"2eaa",x"3547",x"b9f4",x"3c5a",x"3513",x"bc00",x"0000",x"0000",x"3028",x"3547",x"b9f4",x"3639",x"30dd",x"bc00",x"0000",x"0000",x"2eaa",x"3323"),
(x"b9dc",x"3600",x"3069",x"bc00",x"0000",x"0000",x"2658",x"3304",x"b9dc",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"32b8",x"b9dc",x"3c69",x"3069",x"bc00",x"0000",x"0000",x"2658",x"354a"),
(x"ba12",x"3cb7",x"3532",x"ba50",x"b8e8",x"a587",x"2b82",x"1f14",x"ba02",x"3cac",x"3524",x"ba76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"ba12",x"3cb8",x"3076",x"ba76",x"b8b6",x"1fc8",x"2dc6",x"1f14"),
(x"b9dc",x"3600",x"3069",x"bc00",x"0000",x"0000",x"2658",x"3304",x"b9dc",x"3600",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"3304",x"b9dc",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"32b8"),
(x"b9dc",x"3c69",x"3069",x"bc00",x"0000",x"0000",x"2658",x"354a",x"b9dc",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"3573",x"b9dc",x"3c69",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"354a"),
(x"b9dc",x"3600",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"3304",x"b9dc",x"3c69",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"354a",x"b9dc",x"3507",x"364e",x"bc00",x"0000",x"0000",x"2c23",x"32b8"),
(x"ba12",x"3cb1",x"3569",x"b9cc",x"b8ee",x"b4e9",x"2b33",x"1fda",x"ba05",x"3cac",x"3553",x"ba14",x"b8d9",x"b37c",x"2b54",x"2093",x"ba12",x"3cb7",x"3532",x"ba50",x"b8e8",x"a587",x"2b82",x"1f14"),
(x"ba12",x"3cac",x"3587",x"b9e8",x"b889",x"b5d4",x"2b07",x"203c",x"ba05",x"3cac",x"3553",x"ba14",x"b8d9",x"b37c",x"2b54",x"2093",x"ba12",x"3cb1",x"3569",x"b9cc",x"b8ee",x"b4e9",x"2b33",x"1fda"),
(x"ba12",x"3507",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"2d4a",x"b9dc",x"3507",x"364e",x"0000",x"8000",x"bc00",x"318d",x"2d4a",x"ba12",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"333a"),
(x"ba12",x"3507",x"3587",x"204d",x"3c00",x"9cb5",x"2d0f",x"26ad",x"ba07",x"3505",x"3551",x"14ea",x"3c00",x"9dd6",x"2d34",x"2673",x"b9dc",x"3507",x"364e",x"9e0a",x"3c00",x"91bc",x"2c87",x"258a"),
(x"ba12",x"35d7",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2dd5",x"ba08",x"35fd",x"2ce6",x"0000",x"0000",x"3c00",x"31bd",x"2def",x"b9dc",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"b9dc",x"3c69",x"3069",x"ba28",x"391a",x"0000",x"31f8",x"2b85",x"b9dc",x"3c69",x"354b",x"ba28",x"391a",x"0000",x"30ea",x"2b85",x"b9f4",x"3c5a",x"30dd",x"ba28",x"391a",x"0000",x"31e4",x"2bed"),
(x"b9dc",x"3cac",x"364e",x"11bc",x"bc00",x"8000",x"2c87",x"27de",x"ba05",x"3cac",x"3553",x"10ea",x"bc00",x"068d",x"2d33",x"2701",x"ba12",x"3cac",x"3587",x"0e8d",x"bc00",x"0a8d",x"2d0f",x"26bb"),
(x"ba12",x"3c6a",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"3195",x"ba12",x"3c7a",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31a9",x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6"),
(x"ba12",x"3601",x"2c89",x"b9d0",x"342d",x"3915",x"3227",x"3351",x"ba08",x"35fd",x"2ce6",x"b9a5",x"3468",x"3938",x"3231",x"3350",x"ba12",x"35d7",x"2ce6",x"b96d",x"35b1",x"3924",x"322d",x"3342"),
(x"ba01",x"3630",x"2ce6",x"0000",x"0000",x"3c00",x"31c2",x"2e11",x"b9ff",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4",x"b9dc",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"ba12",x"3c78",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"32f4",x"b9dc",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"ba03",x"3c69",x"2ce6",x"0000",x"0000",x"3c00",x"31c0",x"32e0"),
(x"ba08",x"35fd",x"2ce6",x"b9a5",x"3468",x"3938",x"3231",x"3350",x"ba12",x"3601",x"2c89",x"b9d0",x"342d",x"3915",x"3227",x"3351",x"ba01",x"3630",x"2ce6",x"ba49",x"1f45",x"38f2",x"3235",x"3362"),
(x"ba01",x"3630",x"2ce6",x"ba49",x"1f45",x"38f2",x"3235",x"3362",x"ba12",x"3635",x"2c35",x"ba20",x"1881",x"3924",x"3221",x"3363",x"b9ff",x"3c60",x"2ce6",x"ba20",x"9418",x"3925",x"3234",x"3596"),
(x"b9ff",x"3c60",x"2ce6",x"ba20",x"9418",x"3925",x"3234",x"3596",x"ba12",x"3c61",x"2c40",x"b9f4",x"9b5f",x"3957",x"3221",x"3597",x"ba03",x"3c69",x"2ce6",x"b9e5",x"b3cd",x"390b",x"3233",x"359c"),
(x"ba12",x"3c69",x"2c57",x"b9db",x"b485",x"38f4",x"3223",x"359c",x"ba12",x"3c78",x"2ce6",x"b9b2",x"b5ad",x"38d8",x"322c",x"35a7",x"ba03",x"3c69",x"2ce6",x"b9e5",x"b3cd",x"390b",x"3233",x"359c"),
(x"ba12",x"34d8",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"2ab8",x"ba12",x"34db",x"3523",x"bc00",x"0000",x"0000",x"3029",x"2abb",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"4062",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"3947",x"ba12",x"408e",x"3753",x"10ea",x"a1e3",x"3bff",x"39a1",x"3966",x"b940",x"4062",x"374f",x"1e73",x"9cb5",x"3c00",x"39c7",x"3946"),
(x"b940",x"0000",x"374f",x"2138",x"0000",x"3bff",x"39c7",x"3436",x"ba12",x"3227",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"34c4",x"b940",x"4062",x"374f",x"1e73",x"9cb5",x"3c00",x"39c7",x"3946"),
(x"ba12",x"3227",x"3753",x"bc00",x"0000",x"0000",x"30de",x"2890",x"ba12",x"0000",x"3753",x"bc00",x"0000",x"0000",x"30de",x"1e82",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"3cb1",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"31ec",x"ba12",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"31e6",x"ba12",x"3d41",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"329b"),
(x"ba12",x"8000",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"1e82",x"ba12",x"8000",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"1e82",x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c"),
(x"ba12",x"3154",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"280f",x"ba12",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"2af0",x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c"),
(x"ba12",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3583",x"ba12",x"4056",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3563",x"ba12",x"404e",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"355a"),
(x"ba12",x"0000",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"3436",x"ba12",x"3227",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"34c4",x"b940",x"0000",x"374f",x"2138",x"0000",x"3bff",x"39c7",x"3436"),
(x"b9b6",x"3154",x"364d",x"0000",x"bc00",x"15bc",x"38db",x"39de",x"b9b7",x"314b",x"b64f",x"9e3f",x"bc00",x"1418",x"38da",x"3917",x"ba12",x"3154",x"364d",x"9e3f",x"bc00",x"1418",x"38be",x"39de"),
(x"ba12",x"314f",x"b64f",x"0000",x"0000",x"3c00",x"395b",x"3403",x"b9b7",x"314b",x"b64f",x"0000",x"0000",x"3c00",x"396a",x"3402",x"ba12",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"395b",x"3342"),
(x"b941",x"3161",x"b694",x"3c00",x"0000",x"0000",x"38a5",x"3980",x"b941",x"8000",x"b64f",x"3c00",x"8000",x"868d",x"3899",x"3914",x"b941",x"3161",x"b64f",x"3c00",x"0000",x"0000",x"389d",x"3981"),
(x"b941",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404",x"b941",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"397d",x"3342",x"b9b7",x"314b",x"b64f",x"0000",x"868d",x"3c00",x"396a",x"3402"),
(x"b941",x"8000",x"b751",x"0000",x"0cea",x"bc00",x"3ba1",x"34f7",x"b941",x"3161",x"b751",x"0cea",x"8000",x"bc00",x"3ba1",x"355c",x"ba12",x"8000",x"b751",x"11bc",x"868d",x"bc00",x"3bbf",x"34f7"),
(x"3a12",x"3d3f",x"b6b0",x"0000",x"8a8d",x"bc00",x"3aed",x"3929",x"3a12",x"4092",x"b6b0",x"0000",x"8a8d",x"bc00",x"3aed",x"3881",x"b941",x"3d3f",x"b6b0",x"0000",x"8a8d",x"bc00",x"39fa",x"3929"),
(x"b941",x"34e4",x"b751",x"0e8d",x"8000",x"bc00",x"3ba1",x"35af",x"ba12",x"8000",x"b751",x"1018",x"8000",x"bc00",x"3bbf",x"34f7",x"b941",x"3161",x"b751",x"0cea",x"8000",x"bc00",x"3ba1",x"355c"),
(x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7",x"ba12",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"3583",x"ba12",x"3d42",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"329d"),
(x"b941",x"34e4",x"b751",x"0e8d",x"8000",x"bc00",x"3ba1",x"35af",x"b941",x"3cb4",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"37bb",x"ba12",x"3cb5",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"37bc"),
(x"b941",x"4092",x"b751",x"0000",x"23e2",x"bbff",x"3ba1",x"392c",x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929",x"b941",x"3d3f",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"3807"),
(x"b941",x"3cb4",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"37bb",x"b941",x"3d3f",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"3807",x"ba12",x"3cb5",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"37bc"),
(x"ba12",x"3d42",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"329d",x"ba12",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"32a1",x"ba12",x"3cb5",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"31f0"),
(x"3a12",x"3161",x"b751",x"0000",x"8000",x"bc00",x"39f6",x"355c",x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af",x"b941",x"3161",x"b751",x"0cea",x"8000",x"bc00",x"3ba1",x"355c"),
(x"b941",x"34e4",x"b751",x"3c00",x"0000",x"0000",x"3b80",x"380d",x"b941",x"34e4",x"b6b0",x"3c00",x"0000",x"0000",x"3b75",x"380d",x"b941",x"3cb4",x"b751",x"3c00",x"0000",x"0000",x"3b80",x"3926"),
(x"b941",x"3d3f",x"b6b0",x"3c00",x"0000",x"0000",x"3b84",x"3813",x"b941",x"4092",x"b6b0",x"3c00",x"0000",x"0000",x"3b84",x"391f",x"b941",x"3d3f",x"b751",x"3c00",x"0000",x"0000",x"3b8e",x"3813"),
(x"ba72",x"40a7",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3938",x"ba77",x"40a6",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3938",x"ba73",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3935"),
(x"ba49",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba4d",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"393b",x"ba73",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3935"),
(x"ba47",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc7",x"392f",x"ba4b",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba4a",x"4099",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3930"),
(x"ba30",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc4",x"392f",x"ba49",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba47",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc7",x"392f"),
(x"ba29",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"393f",x"ba4d",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"393b",x"ba30",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc4",x"392f"),
(x"ba1e",x"40b8",x"b74a",x"9418",x"257a",x"bbff",x"3bc1",x"3942",x"ba29",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"393f",x"ba27",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392e"),
(x"ba1f",x"408e",x"b74a",x"b075",x"a386",x"bbeb",x"3bc1",x"3929",x"ba26",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"3bc2",x"392c",x"ba27",x"408f",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392a"),
(x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929",x"ba21",x"4092",x"b74a",x"b299",x"a65f",x"bbd3",x"3bc2",x"392c",x"ba1f",x"408e",x"b74a",x"b075",x"a386",x"bbeb",x"3bc1",x"3929"),
(x"ba22",x"4094",x"b74a",x"b0ee",x"1881",x"bbe7",x"3bc2",x"392d",x"ba1e",x"40b8",x"b74a",x"9418",x"257a",x"bbff",x"3bc1",x"3942",x"ba27",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392e"),
(x"b941",x"4092",x"b751",x"0000",x"23e2",x"bbff",x"3ba1",x"392c",x"ba1e",x"40b8",x"b74a",x"9418",x"257a",x"bbff",x"3bc1",x"3942",x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929"),
(x"ba21",x"4092",x"b74a",x"b299",x"a65f",x"bbd3",x"3bc2",x"392c",x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929",x"ba22",x"4094",x"b74a",x"b0ee",x"1881",x"bbe7",x"3bc2",x"392d"),
(x"b940",x"4062",x"374f",x"3c00",x"0000",x"0000",x"394f",x"346c",x"b940",x"4062",x"364d",x"3c00",x"0000",x"0000",x"393e",x"346c",x"b940",x"0000",x"374f",x"3c00",x"0000",x"0000",x"394f",x"3888"),
(x"b9b7",x"40b6",x"364d",x"068d",x"0000",x"bc00",x"393a",x"3867",x"b940",x"4062",x"364d",x"0a8d",x"068d",x"bc00",x"3928",x"383c",x"b940",x"40b6",x"364d",x"0000",x"8000",x"bc00",x"3928",x"3867"),
(x"b9b6",x"3154",x"364d",x"1818",x"8000",x"bc00",x"393a",x"3464",x"ba12",x"0000",x"364d",x"1624",x"8e8d",x"bc00",x"3948",x"340e",x"b940",x"0000",x"364d",x"1a8d",x"8000",x"bc00",x"3929",x"340e"),
(x"b9b7",x"40b6",x"364d",x"3c00",x"0cea",x"0000",x"2d77",x"38e0",x"b9b7",x"40b6",x"b64d",x"3c00",x"0cea",x"8a8d",x"1ca6",x"38e0",x"b9b6",x"3154",x"364d",x"3c00",x"0a8d",x"8e8d",x"2d77",x"3aac"),
(x"b9b7",x"314b",x"b64f",x"0000",x"868d",x"3c00",x"396a",x"3402",x"b9b7",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"396a",x"3887",x"b941",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404"),
(x"b941",x"40b6",x"b64d",x"3c00",x"0000",x"0000",x"38b2",x"3bef",x"b941",x"40b6",x"b694",x"3c00",x"0000",x"0000",x"38b9",x"3bef",x"b941",x"3161",x"b64f",x"3c00",x"0000",x"0000",x"389d",x"3981"),
(x"b941",x"3161",x"b751",x"3c00",x"0000",x"0000",x"38b9",x"397f",x"b941",x"8000",x"b751",x"3c00",x"0000",x"0000",x"38b5",x"3912",x"b941",x"3161",x"b694",x"3c00",x"0000",x"0000",x"38a5",x"3980"),
(x"b9c7",x"3527",x"364c",x"0000",x"3c00",x"8000",x"3199",x"3ab7",x"b9c7",x"3527",x"b696",x"0000",x"3c00",x"8000",x"2de7",x"3ab7",x"3a98",x"3527",x"364c",x"0000",x"3c00",x"8000",x"3199",x"3bfc"),
(x"b9cb",x"3488",x"3650",x"0000",x"bc00",x"0000",x"3af7",x"3689",x"3a94",x"3488",x"3650",x"0000",x"bc00",x"0000",x"3af7",x"37a8",x"b9cb",x"3488",x"b696",x"0000",x"bc00",x"0000",x"3b42",x"3689"),
(x"3a98",x"3527",x"364c",x"0000",x"2631",x"3bff",x"398a",x"39c4",x"3a94",x"3488",x"3650",x"0000",x"2631",x"3bff",x"3976",x"39c4",x"b9c7",x"3527",x"364c",x"0000",x"2631",x"3bff",x"398a",x"3b5b"),
(x"3a1c",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3a40",x"b944",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3b5b",x"3a1c",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3a40"),
(x"b944",x"3449",x"3727",x"0000",x"ba5c",x"38da",x"3920",x"3b5b",x"b944",x"345f",x"3745",x"0000",x"ba15",x"3932",x"3929",x"3b5b",x"3a1c",x"3449",x"3727",x"0000",x"ba5c",x"38da",x"3920",x"3a40"),
(x"3af9",x"40b3",x"377b",x"39af",x"39a0",x"8000",x"370a",x"3aba",x"3aef",x"40b8",x"376a",x"3b44",x"36ae",x"0000",x"3718",x"3ab8",x"3af9",x"40b3",x"b74a",x"3a61",x"38d2",x"0000",x"370a",x"3910"),
(x"ba29",x"40b3",x"377b",x"8000",x"39b1",x"399e",x"3692",x"3ab6",x"ba1e",x"40b8",x"376a",x"0000",x"3587",x"3b81",x"36a6",x"3ab2",x"3af9",x"40b3",x"377b",x"8000",x"38b6",x"3a76",x"3692",x"3863"),
(x"3af9",x"40b3",x"377b",x"8000",x"38b6",x"3a76",x"3692",x"3863",x"3b1e",x"40ab",x"37c7",x"8000",x"3a96",x"388a",x"367e",x"385b",x"ba29",x"40b3",x"377b",x"8000",x"39b1",x"399e",x"3692",x"3ab6"),
(x"3b1e",x"40ab",x"37c7",x"8000",x"3a96",x"388a",x"367e",x"385b",x"3b43",x"40a7",x"3805",x"0000",x"3b38",x"36e2",x"366b",x"3852",x"ba4d",x"40ab",x"37c7",x"0000",x"3af8",x"37d8",x"367f",x"3abe"),
(x"3b43",x"40a7",x"3805",x"0000",x"3b38",x"36e2",x"366b",x"3852",x"3b48",x"40a6",x"380b",x"0000",x"3824",x"3ad7",x"3656",x"384c",x"ba72",x"40a7",x"3805",x"8000",x"3ae3",x"3811",x"366b",x"3ac9"),
(x"3b48",x"40a6",x"380b",x"0000",x"3824",x"3ad7",x"3656",x"384c",x"3b48",x"40a4",x"380c",x"0000",x"b0b3",x"3be9",x"3642",x"384c",x"ba77",x"40a6",x"380b",x"0000",x"34ea",x"3b9c",x"3656",x"3ad1"),
(x"3b48",x"40a4",x"380c",x"0000",x"b0b3",x"3be9",x"3642",x"384c",x"3b44",x"40a2",x"3807",x"8000",x"ba4c",x"38ee",x"362d",x"3853",x"ba77",x"40a4",x"380c",x"0000",x"b607",x"3b69",x"3641",x"3ad1"),
(x"3b44",x"40a2",x"3807",x"8000",x"ba4c",x"38ee",x"362d",x"3853",x"3b1a",x"409b",x"37ba",x"0000",x"baba",x"3854",x"3619",x"385c",x"ba73",x"40a2",x"3807",x"0000",x"ba9a",x"3884",x"362d",x"3acb"),
(x"3b1a",x"409b",x"37ba",x"0000",x"3897",x"3a8d",x"37c2",x"3974",x"3b1c",x"409b",x"37bd",x"8000",x"3873",x"3aa5",x"37b7",x"3971",x"ba49",x"409b",x"37ba",x"0000",x"3897",x"3a8d",x"37c2",x"3ace"),
(x"3b1c",x"409b",x"37bd",x"8000",x"3873",x"3aa5",x"37b7",x"3971",x"3b1c",x"409a",x"37c0",x"0000",x"32ec",x"3bcf",x"37ac",x"3971",x"ba4b",x"409b",x"37bd",x"0000",x"384b",x"3abf",x"37b7",x"3ad1"),
(x"3b1c",x"409a",x"37c0",x"0000",x"32ec",x"3bcf",x"37ac",x"3971",x"3b1b",x"4099",x"37bf",x"0000",x"b654",x"3b58",x"37a1",x"3972",x"ba4b",x"409a",x"37c0",x"8000",x"8cea",x"3c00",x"37ac",x"3ad1"),
(x"3b1b",x"4099",x"37bf",x"0000",x"b654",x"3b58",x"37a1",x"3972",x"3b18",x"4098",x"37b7",x"0000",x"bbda",x"3211",x"3795",x"3976",x"ba4a",x"4099",x"37bf",x"8000",x"b927",x"3a1e",x"37a1",x"3ad1"),
(x"3b18",x"4098",x"37b7",x"0000",x"bbda",x"3211",x"3795",x"3976",x"3b01",x"4098",x"3785",x"0000",x"bbfe",x"28cc",x"378a",x"397c",x"ba47",x"4098",x"37b7",x"8000",x"bbf8",x"2d73",x"3795",x"3acd"),
(x"3b01",x"4098",x"3785",x"0000",x"ba3a",x"3905",x"380f",x"3947",x"3af8",x"4096",x"3773",x"0000",x"b9da",x"3973",x"3809",x"394c",x"ba30",x"4098",x"3785",x"0000",x"ba3a",x"3905",x"380f",x"3ad7"),
(x"3af8",x"4096",x"3773",x"0000",x"b9da",x"3973",x"3809",x"394c",x"3af3",x"4094",x"3767",x"8000",x"b745",x"3b20",x"3802",x"3950",x"ba27",x"4096",x"3773",x"8000",x"b967",x"39e6",x"3809",x"3ad2"),
(x"3af3",x"4094",x"3767",x"8000",x"b745",x"3b20",x"3802",x"3950",x"3af1",x"4092",x"3766",x"0000",x"ac55",x"3bfb",x"37f9",x"3951",x"ba22",x"4094",x"3767",x"8000",x"b449",x"3bb5",x"3802",x"3acf"),
(x"3af1",x"4092",x"3766",x"0000",x"3bf8",x"2da0",x"37f8",x"3986",x"3af6",x"4092",x"3775",x"0000",x"3ba1",x"34ce",x"37ee",x"3983",x"ba21",x"4092",x"3766",x"0000",x"3bf8",x"2d9e",x"37f8",x"3ac8"),
(x"3af6",x"4092",x"3775",x"0000",x"3ba1",x"34ce",x"37ee",x"3983",x"3afa",x"4091",x"3778",x"0000",x"326d",x"3bd6",x"37e3",x"397e",x"ba26",x"4092",x"3775",x"8000",x"3a53",x"38e6",x"37ee",x"3acc"),
(x"3afa",x"4091",x"3778",x"0000",x"326d",x"3bd6",x"37e3",x"397e",x"3af8",x"408f",x"3777",x"8000",x"b682",x"3b4e",x"37d8",x"3980",x"ba29",x"4091",x"3778",x"0000",x"26d5",x"3bff",x"37e3",x"3ad1"),
(x"3af8",x"408f",x"3777",x"8000",x"b682",x"3b4e",x"37d8",x"3980",x"3af0",x"408e",x"3769",x"8000",x"bb26",x"372c",x"37cd",x"3985",x"ba27",x"408f",x"3777",x"0000",x"b8ed",x"3a4d",x"37d8",x"3acf"),
(x"3af8",x"4096",x"3773",x"39a4",x"b9ac",x"0000",x"382d",x"39a9",x"3af8",x"4096",x"b74a",x"3a2e",x"b913",x"0000",x"382d",x"3888",x"3af3",x"4094",x"3767",x"3b41",x"b6be",x"8000",x"3829",x"39a6"),
(x"3b48",x"40a4",x"380c",x"3b97",x"b50c",x"0000",x"36c9",x"3ad1",x"3b48",x"40a4",x"b74a",x"3b97",x"b50b",x"8000",x"36c9",x"3910",x"3b44",x"40a2",x"3807",x"38f8",x"ba45",x"0000",x"36ba",x"3acd"),
(x"3b01",x"4098",x"3785",x"391e",x"ba25",x"0000",x"3832",x"39ac",x"3b01",x"4098",x"b74a",x"391e",x"ba25",x"0000",x"3832",x"3888",x"3af8",x"4096",x"3773",x"39a4",x"b9ac",x"0000",x"382d",x"39a9"),
(x"3af0",x"408e",x"3769",x"361a",x"bb65",x"8000",x"3813",x"39ca",x"3af0",x"408e",x"b74a",x"31b5",x"bbdf",x"0000",x"3813",x"38cb",x"3ae3",x"408e",x"3753",x"0000",x"bc00",x"0000",x"380f",x"39c7"),
(x"3b48",x"40a4",x"380c",x"3b97",x"b50c",x"0000",x"36c9",x"3ad1",x"3b48",x"40a6",x"380b",x"3bc1",x"33d8",x"8000",x"36d8",x"3ad0",x"3b48",x"40a4",x"b74a",x"3b97",x"b50b",x"8000",x"36c9",x"3910"),
(x"3b18",x"4098",x"37b7",x"32b5",x"bbd2",x"0000",x"3793",x"396c",x"3b18",x"4098",x"b74a",x"2dde",x"bbf7",x"8000",x"3793",x"3872",x"3b01",x"4098",x"3785",x"2918",x"bbfe",x"0000",x"378b",x"3968"),
(x"3af8",x"408f",x"3777",x"3ac3",x"b845",x"0000",x"3817",x"39cd",x"3af8",x"408f",x"b74a",x"399f",x"b9b0",x"068d",x"3817",x"38cc",x"3af0",x"408e",x"3769",x"361a",x"bb65",x"8000",x"3813",x"39ca"),
(x"3b48",x"40a6",x"380b",x"3bc1",x"33d8",x"8000",x"36d8",x"3ad0",x"3b43",x"40a7",x"3805",x"37c0",x"3aff",x"8000",x"36e6",x"3acb",x"3b48",x"40a6",x"b74a",x"3af6",x"37df",x"0000",x"36d8",x"3910"),
(x"3b1b",x"4099",x"37bf",x"3b8d",x"b548",x"8000",x"379b",x"3970",x"3b1b",x"4099",x"b74a",x"3aa8",x"b86e",x"0000",x"379b",x"3872",x"3b18",x"4098",x"37b7",x"32b5",x"bbd2",x"0000",x"3793",x"396c"),
(x"3afa",x"4091",x"3778",x"3bdb",x"31fa",x"8000",x"381b",x"39cd",x"3afa",x"4091",x"b74a",x"3bdb",x"31fa",x"8000",x"381b",x"38cc",x"3af8",x"408f",x"3777",x"3ac3",x"b845",x"0000",x"3817",x"39cd"),
(x"3b43",x"40a7",x"3805",x"37c0",x"3aff",x"8000",x"36e6",x"3acb",x"3b1e",x"40ab",x"37c7",x"379e",x"3b08",x"0000",x"36f6",x"3ac3",x"3b43",x"40a7",x"b74a",x"3671",x"3b52",x"0000",x"36e6",x"3910"),
(x"3b1c",x"409a",x"37c0",x"3bfc",x"abd5",x"8000",x"37a3",x"3971",x"3b1c",x"409a",x"b74a",x"3bfc",x"abd5",x"8000",x"37a3",x"3873",x"3b1b",x"4099",x"37bf",x"3b8d",x"b548",x"8000",x"379b",x"3970"),
(x"3afa",x"4091",x"3778",x"3bdb",x"31fa",x"8000",x"381b",x"39cd",x"3af6",x"4092",x"3775",x"38a6",x"3a82",x"0000",x"381f",x"39cc",x"3afa",x"4091",x"b74a",x"3bdb",x"31fa",x"8000",x"381b",x"38cc"),
(x"3b1e",x"40ab",x"37c7",x"379e",x"3b08",x"0000",x"36f6",x"3ac3",x"3af9",x"40b3",x"377b",x"39af",x"39a0",x"8000",x"370a",x"3aba",x"3b1e",x"40ab",x"b74a",x"3890",x"3a91",x"8000",x"36f6",x"3910"),
(x"3b1c",x"409a",x"37c0",x"3bfc",x"abd5",x"8000",x"37a3",x"3971",x"3b1c",x"409b",x"37bd",x"3bb8",x"3431",x"8000",x"37ab",x"396e",x"3b1c",x"409a",x"b74a",x"3bfc",x"abd5",x"8000",x"37a3",x"3873"),
(x"3af6",x"4092",x"3775",x"38a6",x"3a82",x"0000",x"381f",x"39cc",x"3af1",x"4092",x"3766",x"3033",x"3bee",x"0000",x"3824",x"39c5",x"3af6",x"4092",x"b74a",x"35d6",x"3b72",x"0000",x"3820",x"38cc"),
(x"3b1c",x"409b",x"37bd",x"3bb8",x"3431",x"8000",x"37ab",x"396e",x"3b1a",x"409b",x"37ba",x"3ad7",x"3825",x"0000",x"37b3",x"396b",x"3b1c",x"409b",x"b74a",x"3b4e",x"3681",x"0000",x"37ab",x"3873"),
(x"3af3",x"4094",x"3767",x"3b41",x"b6be",x"8000",x"3829",x"39a6",x"3af3",x"4094",x"b74a",x"3ba9",x"b498",x"0000",x"3829",x"3888",x"3af1",x"4092",x"3766",x"3be9",x"b0c2",x"0000",x"3824",x"39a5"),
(x"3b44",x"40a2",x"3807",x"38f8",x"ba45",x"0000",x"36ba",x"3acd",x"3b44",x"40a2",x"b74a",x"3892",x"ba90",x"068d",x"36bb",x"3910",x"3b1a",x"409b",x"37ba",x"3863",x"bab0",x"0000",x"36a6",x"3ac4"),
(x"3af0",x"408e",x"3769",x"8000",x"bb26",x"372c",x"37cd",x"3985",x"3ae3",x"408e",x"3753",x"0000",x"bc00",x"0000",x"37c3",x"398c",x"ba1f",x"408e",x"3769",x"0000",x"bbd1",x"32c7",x"37cd",x"3aca"),
(x"3ae3",x"408e",x"3753",x"8cea",x"a1fd",x"3bff",x"3bf9",x"3966",x"3ae3",x"4062",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"3947",x"3a11",x"4062",x"374f",x"a018",x"9953",x"3c00",x"3bd3",x"3946"),
(x"3ae3",x"4062",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"3947",x"3ae3",x"3227",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"34c4",x"3a11",x"4062",x"374f",x"a018",x"9953",x"3c00",x"3bd3",x"3946"),
(x"3ae3",x"3227",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"34c4",x"3ae3",x"0000",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"3436",x"3a11",x"0000",x"374f",x"a138",x"0000",x"3bff",x"3bd3",x"3436"),
(x"3ae3",x"314f",x"b64f",x"224c",x"bbff",x"11bc",x"38f7",x"3917",x"3a88",x"314b",x"b64f",x"1e3f",x"bc00",x"1418",x"38db",x"3917",x"3ae3",x"3154",x"364d",x"1e3f",x"bc00",x"1418",x"38f7",x"39de"),
(x"3ae3",x"314f",x"b64f",x"0000",x"0000",x"3c00",x"399f",x"3403",x"3ae3",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"399f",x"3342",x"3a88",x"314b",x"b64f",x"0000",x"0000",x"3c00",x"3990",x"3402"),
(x"3a12",x"8000",x"b64f",x"bc00",x"0000",x"0000",x"3899",x"3914",x"3a12",x"3161",x"b694",x"bc00",x"0000",x"0000",x"388e",x"3980",x"3a12",x"3161",x"b64f",x"bc00",x"0000",x"0000",x"3895",x"3981"),
(x"3a12",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"397d",x"3342",x"3a12",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404",x"3a88",x"314b",x"b64f",x"0000",x"868d",x"3c00",x"3990",x"3402"),
(x"3a12",x"3161",x"b751",x"0000",x"8000",x"bc00",x"39f6",x"355c",x"3a12",x"8000",x"b751",x"0000",x"0cea",x"bc00",x"39f6",x"34f7",x"3ae3",x"8000",x"b751",x"8a8d",x"0a8d",x"bc00",x"39d8",x"34f7"),
(x"b941",x"3cb4",x"b751",x"0000",x"bc00",x"0000",x"39d2",x"3494",x"b941",x"3cb4",x"b6af",x"0000",x"bc00",x"0000",x"39d2",x"34a6",x"3a12",x"3cb4",x"b751",x"0000",x"bc00",x"0000",x"3bc8",x"3494"),
(x"3ae3",x"8000",x"b751",x"8a8d",x"0a8d",x"bc00",x"39d8",x"34f7",x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af",x"3a12",x"3161",x"b751",x"0000",x"8000",x"bc00",x"39f6",x"355c"),
(x"3a12",x"3cb4",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"37bb",x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807",x"b941",x"3cb4",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"37bb"),
(x"3ae3",x"3154",x"b751",x"9018",x"8000",x"bc00",x"39d8",x"355b",x"3ae3",x"3cb5",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"37bc",x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af"),
(x"3ae3",x"3d42",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"3807",x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807"),
(x"3a12",x"3cb4",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"37bb",x"3ae3",x"3cb5",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"37bc",x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807"),
(x"3a12",x"34e4",x"b751",x"0000",x"3c00",x"8000",x"3bc8",x"34b8",x"3a12",x"34e4",x"b6b0",x"0000",x"3c00",x"8000",x"3bc8",x"34a6",x"b941",x"34e4",x"b751",x"0000",x"3c00",x"8000",x"39d2",x"34b8"),
(x"3a12",x"34e4",x"b751",x"bc00",x"0000",x"0000",x"3b69",x"380d",x"3a12",x"3cb4",x"b751",x"bc00",x"0000",x"0000",x"3b69",x"3926",x"3a12",x"34e4",x"b6b0",x"bc00",x"0000",x"0000",x"3b75",x"380d"),
(x"3a12",x"4092",x"b751",x"bc00",x"0000",x"0000",x"3b90",x"3922",x"3a12",x"4092",x"b6b0",x"bc00",x"0000",x"0000",x"3b9e",x"3922",x"3a12",x"3d3f",x"b751",x"bc00",x"0000",x"0000",x"3b90",x"3814"),
(x"b941",x"4092",x"b6b0",x"0000",x"bc00",x"0000",x"39ce",x"3475",x"3a12",x"4092",x"b6b0",x"0000",x"bc00",x"0000",x"3bcd",x"3475",x"b941",x"4092",x"b751",x"0000",x"bc00",x"0000",x"39ce",x"345e"),
(x"3a11",x"4062",x"374f",x"a018",x"9953",x"3c00",x"3bd3",x"3946",x"b940",x"4062",x"374f",x"1e73",x"9cb5",x"3c00",x"39c7",x"3946",x"3ae3",x"408e",x"3753",x"8cea",x"a1fd",x"3bff",x"3bf9",x"3966"),
(x"3b48",x"40a4",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3936",x"3b48",x"40a6",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3938",x"3b44",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3935"),
(x"3b1a",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3931",x"3b44",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3935",x"3b1e",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"393b"),
(x"3b18",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d0",x"392f",x"3b1b",x"4099",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3930",x"3b1c",x"409b",x"b74a",x"068d",x"0000",x"bc00",x"39cf",x"3931"),
(x"3b01",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d3",x"392f",x"3b18",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d0",x"392f",x"3b1a",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3931"),
(x"3af9",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"393f",x"3b01",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d3",x"392f",x"3b1e",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"393b"),
(x"3b01",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d3",x"392f",x"3af9",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"393f",x"3af8",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392e"),
(x"3af0",x"408e",x"b74a",x"3075",x"a386",x"bbeb",x"39d6",x"3929",x"3af8",x"408f",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392a",x"3af6",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"39d5",x"392c"),
(x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3af0",x"408e",x"b74a",x"3075",x"a386",x"bbeb",x"39d6",x"3929",x"3af1",x"4092",x"b74a",x"3299",x"a666",x"bbd3",x"39d5",x"392c"),
(x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942",x"3af3",x"4094",x"b74a",x"30ed",x"1881",x"bbe7",x"39d5",x"392d",x"3af8",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392e"),
(x"3a12",x"4092",x"b751",x"068d",x"21e3",x"bbff",x"39f6",x"392c",x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942"),
(x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3af1",x"4092",x"b74a",x"3299",x"a666",x"bbd3",x"39d5",x"392c",x"3af3",x"4094",x"b74a",x"30ed",x"1881",x"bbe7",x"39d5",x"392d"),
(x"3aef",x"40b8",x"b74a",x"0000",x"3c00",x"8000",x"346a",x"38f0",x"3aef",x"40b8",x"376a",x"0000",x"3c00",x"8000",x"316c",x"38f0",x"ba1e",x"40b8",x"b74a",x"0000",x"3c00",x"8000",x"346a",x"3a98"),
(x"3a12",x"4092",x"b751",x"068d",x"21e3",x"bbff",x"39f6",x"392c",x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942",x"b941",x"4092",x"b751",x"0000",x"23e2",x"bbff",x"3ba1",x"392c"),
(x"b941",x"34e4",x"b6b0",x"0000",x"0cea",x"bc00",x"39fa",x"37b1",x"3a12",x"34e4",x"b6b0",x"0000",x"0cea",x"bc00",x"3aed",x"37b1",x"b941",x"3cb4",x"b6af",x"0000",x"0cea",x"bc00",x"39fa",x"3687"),
(x"3a11",x"4062",x"374f",x"0000",x"bc00",x"0000",x"3166",x"38dd",x"3a11",x"4062",x"364d",x"0000",x"bc00",x"0000",x"3166",x"38eb",x"b940",x"4062",x"374f",x"0000",x"bc00",x"0000",x"3592",x"38dd"),
(x"3a11",x"4062",x"364d",x"9018",x"8000",x"bc00",x"36e3",x"383c",x"3a11",x"40b6",x"364d",x"0000",x"8000",x"bc00",x"36e3",x"3866",x"b940",x"4062",x"364d",x"0a8d",x"068d",x"bc00",x"3928",x"383c"),
(x"3a11",x"4062",x"374f",x"bc00",x"0000",x"0000",x"3953",x"341e",x"3a11",x"0000",x"374f",x"bc00",x"0000",x"0000",x"3953",x"3861",x"3a11",x"4062",x"364d",x"bc00",x"0000",x"0000",x"3964",x"341e"),
(x"b941",x"40b6",x"b694",x"0000",x"068d",x"3c00",x"2da6",x"375f",x"3a12",x"40b6",x"b694",x"0000",x"068d",x"3c00",x"2da6",x"38d9",x"b941",x"3161",x"b694",x"0000",x"068d",x"3c00",x"3501",x"375f"),
(x"3a11",x"4062",x"364d",x"9018",x"8000",x"bc00",x"36e3",x"383c",x"3a88",x"40b6",x"364d",x"8e8d",x"068d",x"bc00",x"36bf",x"3866",x"3a11",x"40b6",x"364d",x"0000",x"8000",x"bc00",x"36e3",x"3866"),
(x"3a11",x"0000",x"364d",x"9ac2",x"8000",x"bc00",x"36e3",x"340e",x"3ae3",x"0000",x"364d",x"968d",x"8e8d",x"bc00",x"36a4",x"340e",x"3a87",x"3154",x"364d",x"96f6",x"0000",x"bc00",x"36c0",x"3464"),
(x"3a88",x"40b6",x"364d",x"bc00",x"0cea",x"0000",x"315f",x"3aac",x"3a87",x"3154",x"364d",x"bc00",x"0a8d",x"8e8d",x"315f",x"38e0",x"3a88",x"40b6",x"b64d",x"bc00",x"0cea",x"8a8d",x"2d91",x"3aac"),
(x"3a12",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"397d",x"3887",x"3a88",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"3990",x"3887",x"3a12",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404"),
(x"3a11",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"374a",x"3a12",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"374a",x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd"),
(x"3a12",x"3161",x"b694",x"0000",x"bc00",x"0000",x"3bc8",x"3494",x"3a12",x"3161",x"b751",x"0000",x"bc00",x"0000",x"3bc8",x"347e",x"b941",x"3161",x"b694",x"0000",x"bc00",x"0000",x"39d2",x"3494"),
(x"3a87",x"3154",x"364d",x"96f6",x"0000",x"bc00",x"36c0",x"3464",x"3ae3",x"0000",x"364d",x"968d",x"8e8d",x"bc00",x"36a4",x"340e",x"3ae3",x"3154",x"364d",x"0000",x"8000",x"bc00",x"36a4",x"3464"),
(x"3a12",x"3161",x"b694",x"bc00",x"0000",x"0000",x"388e",x"3980",x"3a12",x"40b6",x"b694",x"bc00",x"0000",x"0000",x"3879",x"3bef",x"3a12",x"3161",x"b64f",x"bc00",x"0000",x"0000",x"3895",x"3981"),
(x"3a12",x"8000",x"b64f",x"bc00",x"8000",x"868d",x"3899",x"3914",x"3a12",x"8000",x"b751",x"bc00",x"8000",x"868d",x"387d",x"3912",x"3a12",x"3161",x"b694",x"bc00",x"0000",x"0000",x"388e",x"3980"),
(x"b941",x"3d3f",x"b6b0",x"0000",x"3c00",x"8000",x"39ce",x"3447",x"b941",x"3d3f",x"b751",x"0000",x"3c00",x"8000",x"39ce",x"345e",x"3a12",x"3d3f",x"b6b0",x"0000",x"3c00",x"8000",x"3bcd",x"3447"),
(x"b944",x"31a5",x"3649",x"0000",x"8000",x"bc00",x"38f2",x"3b5b",x"3a1c",x"31a5",x"3649",x"0000",x"8000",x"bc00",x"38f2",x"39e5",x"3a1c",x"349b",x"3649",x"0000",x"8000",x"bc00",x"38ba",x"39e5"),
(x"b944",x"3468",x"3748",x"0000",x"ae16",x"3bf6",x"3933",x"3b5b",x"3a1c",x"3468",x"3748",x"0000",x"a67a",x"3bff",x"3933",x"3a40",x"3a1c",x"345f",x"3745",x"8000",x"b970",x"39dd",x"3929",x"3a40"),
(x"b944",x"3449",x"3727",x"0000",x"0000",x"3c00",x"3920",x"3b5b",x"3a1c",x"3449",x"3727",x"0000",x"0000",x"3c00",x"3920",x"39e5",x"3a1c",x"31a5",x"3727",x"0000",x"0000",x"3c00",x"38f2",x"39e5"),
(x"b944",x"34b9",x"3649",x"0000",x"3c00",x"1a59",x"395b",x"3b5b",x"3a1c",x"34b9",x"3649",x"0000",x"3c00",x"1a59",x"395b",x"3a40",x"3a1c",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3a40"),
(x"b944",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3b5b",x"3a1c",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3a40",x"3a1c",x"3468",x"3748",x"0000",x"a67a",x"3bff",x"3933",x"3a40"),
(x"b944",x"31a5",x"3727",x"0000",x"bc00",x"0000",x"3976",x"3b5b",x"3a1c",x"31a5",x"3727",x"0000",x"bc00",x"0000",x"3976",x"39e5",x"3a1c",x"31a5",x"3649",x"0000",x"bc00",x"0000",x"395b",x"39e5"),
(x"b9bc",x"3d46",x"b64b",x"0000",x"3c00",x"8000",x"1d3c",x"3ab8",x"3a8c",x"3d46",x"b64b",x"0000",x"3c00",x"8000",x"1d3c",x"3bfb",x"3a8c",x"3d46",x"3653",x"0000",x"3c00",x"8000",x"2d82",x"3bfb"),
(x"3a88",x"3d1e",x"3657",x"0000",x"bc00",x"0000",x"3b46",x"37ad",x"3a88",x"3d1e",x"b64b",x"0000",x"bc00",x"0000",x"3b90",x"37ad",x"b9c0",x"3d1e",x"b64b",x"0000",x"bc00",x"0000",x"3b90",x"368f"),
(x"3a88",x"3d1e",x"3657",x"0000",x"2631",x"3bff",x"398a",x"39c7",x"b9c0",x"3d1e",x"3657",x"0000",x"2631",x"3bff",x"398a",x"3b5b",x"b9bc",x"3d46",x"3653",x"0000",x"2631",x"3bff",x"399e",x"3b5b"),
(x"ba29",x"40b3",x"b74a",x"ba61",x"38d2",x"0000",x"3726",x"3911",x"ba1e",x"40b8",x"b74a",x"bb44",x"36ae",x"0000",x"3718",x"3911",x"ba1e",x"40b8",x"376a",x"bb44",x"36ae",x"0000",x"3719",x"3abb"),
(x"ba27",x"4096",x"b74a",x"ba2e",x"b913",x"0000",x"3828",x"39ad",x"ba27",x"4096",x"3773",x"b9a4",x"b9ac",x"0000",x"3828",x"3acd",x"ba22",x"4094",x"3767",x"bb41",x"b6be",x"8000",x"382d",x"3ac9"),
(x"ba77",x"40a4",x"b74a",x"bb97",x"b50b",x"0000",x"3767",x"3911",x"ba77",x"40a4",x"380c",x"bb97",x"b50c",x"0000",x"3767",x"3ad1",x"ba73",x"40a2",x"3807",x"b8f8",x"ba45",x"0000",x"3775",x"3acc"),
(x"ba30",x"4098",x"b74a",x"b91e",x"ba25",x"0000",x"3824",x"39ad",x"ba30",x"4098",x"3785",x"b91e",x"ba25",x"0000",x"3824",x"3ad1",x"ba27",x"4096",x"3773",x"b9a4",x"b9ac",x"0000",x"3828",x"3acd"),
(x"ba1f",x"408e",x"b74a",x"b1b5",x"bbdf",x"0000",x"3820",x"39cf",x"ba1f",x"408e",x"3769",x"b61a",x"bb65",x"8000",x"381f",x"3acd",x"ba12",x"408e",x"3753",x"0000",x"bc00",x"0000",x"3824",x"3aca"),
(x"ba77",x"40a4",x"b74a",x"bb97",x"b50b",x"0000",x"3767",x"3911",x"ba77",x"40a6",x"b74a",x"baf6",x"37df",x"868d",x"3759",x"3911",x"ba77",x"40a6",x"380b",x"bbc1",x"33d8",x"8000",x"3759",x"3ad0"),
(x"ba47",x"4098",x"b74a",x"adde",x"bbf7",x"0000",x"37e4",x"3872",x"ba47",x"4098",x"37b7",x"b2b5",x"bbd2",x"0000",x"37e4",x"396c",x"ba30",x"4098",x"3785",x"a918",x"bbfe",x"0000",x"37eb",x"3967"),
(x"ba27",x"408f",x"b74a",x"b99f",x"b9b0",x"0000",x"381b",x"39cf",x"ba27",x"408f",x"3777",x"bac3",x"b845",x"0000",x"381b",x"3ad0",x"ba1f",x"408e",x"3769",x"b61a",x"bb65",x"8000",x"381f",x"3acd"),
(x"ba77",x"40a6",x"b74a",x"baf6",x"37df",x"868d",x"3759",x"3911",x"ba72",x"40a7",x"b74a",x"b671",x"3b52",x"868d",x"374b",x"3911",x"ba72",x"40a7",x"3805",x"b7c0",x"3aff",x"0000",x"374b",x"3acc"),
(x"ba4a",x"4099",x"b74a",x"baa8",x"b86e",x"0000",x"37dc",x"3872",x"ba4a",x"4099",x"37bf",x"bb8d",x"b548",x"8000",x"37db",x"3970",x"ba47",x"4098",x"37b7",x"b2b5",x"bbd2",x"0000",x"37e4",x"396c"),
(x"ba29",x"4091",x"b74a",x"bbdb",x"31fa",x"0000",x"3817",x"39cf",x"ba29",x"4091",x"3778",x"bbdb",x"31fb",x"0000",x"3817",x"3ad1",x"ba27",x"408f",x"3777",x"bac3",x"b845",x"0000",x"381b",x"3ad0"),
(x"ba72",x"40a7",x"b74a",x"b671",x"3b52",x"868d",x"374b",x"3911",x"ba4d",x"40ab",x"b74a",x"b890",x"3a91",x"0000",x"373a",x"3911",x"ba4d",x"40ab",x"37c7",x"b79e",x"3b08",x"0000",x"373b",x"3ac5"),
(x"ba4b",x"409a",x"b74a",x"bbfc",x"abd5",x"0000",x"37d3",x"3872",x"ba4b",x"409a",x"37c0",x"bbfc",x"abd5",x"0000",x"37d3",x"3971",x"ba4a",x"4099",x"37bf",x"bb8d",x"b548",x"8000",x"37db",x"3970"),
(x"ba29",x"4091",x"b74a",x"bbdb",x"31fa",x"0000",x"3817",x"39cf",x"ba26",x"4092",x"b74a",x"b5d6",x"3b72",x"8000",x"3813",x"39cf",x"ba26",x"4092",x"3775",x"b8a6",x"3a82",x"0000",x"3813",x"3acf"),
(x"ba4d",x"40ab",x"b74a",x"b890",x"3a91",x"0000",x"373a",x"3911",x"ba29",x"40b3",x"b74a",x"ba61",x"38d2",x"0000",x"3726",x"3911",x"ba29",x"40b3",x"377b",x"b9af",x"39a0",x"8000",x"3728",x"3abe"),
(x"ba4b",x"409a",x"b74a",x"bbfc",x"abd5",x"0000",x"37d3",x"3872",x"ba4b",x"409b",x"b74a",x"bb4e",x"3681",x"068d",x"37cb",x"3872",x"ba4b",x"409b",x"37bd",x"bbb8",x"3431",x"8000",x"37cb",x"396e"),
(x"ba26",x"4092",x"b74a",x"b5d6",x"3b72",x"8000",x"3813",x"39cf",x"ba21",x"4092",x"b74a",x"b033",x"3bee",x"0000",x"380f",x"39cf",x"ba21",x"4092",x"3766",x"b033",x"3bee",x"0000",x"380f",x"3aca"),
(x"ba4b",x"409b",x"b74a",x"bb4e",x"3681",x"068d",x"37cb",x"3872",x"ba49",x"409b",x"b74a",x"bad7",x"3825",x"0000",x"37c3",x"3872",x"ba49",x"409b",x"37ba",x"bad7",x"3825",x"0000",x"37c3",x"396c"),
(x"ba22",x"4094",x"b74a",x"bba9",x"b498",x"8000",x"382d",x"39ad",x"ba22",x"4094",x"3767",x"bb41",x"b6be",x"8000",x"382d",x"3ac9",x"ba21",x"4092",x"3766",x"bbe9",x"b0c2",x"0000",x"3832",x"3ac9"),
(x"ba73",x"40a2",x"b74a",x"b892",x"ba90",x"0000",x"3775",x"3911",x"ba73",x"40a2",x"3807",x"b8f8",x"ba45",x"0000",x"3775",x"3acc",x"ba49",x"409b",x"37ba",x"b863",x"bab0",x"0000",x"378a",x"3ac3"),
(x"ba05",x"3d46",x"b544",x"ba14",x"38d9",x"337c",x"2dd6",x"20e8",x"ba02",x"3d46",x"b515",x"ba7c",x"38ae",x"1c81",x"2db6",x"20d0",x"ba12",x"3d3b",x"b522",x"ba50",x"38e8",x"2604",x"2dbf",x"21f1"),
(x"ba02",x"3d46",x"b515",x"ba7c",x"38ae",x"1c81",x"2db6",x"20d0",x"ba03",x"3d45",x"b075",x"baa1",x"3878",x"a594",x"2b88",x"20ca",x"ba12",x"3d3a",x"b07b",x"ba7d",x"38ad",x"9e59",x"2b8b",x"21f1"),
(x"ba03",x"3d45",x"b075",x"baa1",x"3878",x"a594",x"2b88",x"20ca",x"ba09",x"3d45",x"b010",x"ba60",x"3855",x"b446",x"2b42",x"20ee",x"ba12",x"3d3f",x"b00e",x"ba6d",x"3864",x"b364",x"2b40",x"219c"),
(x"b9dc",x"3d46",x"aca4",x"9d38",x"3c00",x"8cea",x"2392",x"2238",x"ba03",x"3d45",x"b075",x"a49b",x"3bff",x"1418",x"26b4",x"23d9",x"ba02",x"3d46",x"b515",x"9f10",x"3c00",x"1018",x"2b3f",x"23cc"),
(x"ba12",x"3d46",x"af74",x"1f79",x"3c00",x"9c81",x"25b4",x"243e",x"b9dc",x"3d46",x"aca4",x"9d38",x"3c00",x"8cea",x"2392",x"2238",x"ba12",x"3d46",x"aca4",x"0000",x"3c00",x"8000",x"2392",x"243e"),
(x"ba09",x"3d45",x"b010",x"20d0",x"3bff",x"a081",x"262a",x"240d",x"ba03",x"3d45",x"b075",x"a49b",x"3bff",x"1418",x"26b4",x"23d9",x"b9dc",x"3d46",x"aca4",x"9d38",x"3c00",x"8cea",x"2392",x"2238"),
(x"ba09",x"4070",x"b010",x"0000",x"bc00",x"0000",x"2d20",x"248a",x"b9dc",x"4070",x"aca4",x"0e8d",x"bc00",x"8000",x"2c87",x"257b",x"ba03",x"4070",x"b075",x"0000",x"bc00",x"0000",x"2d42",x"24ab"),
(x"ba12",x"4070",x"af8a",x"0000",x"bc00",x"0000",x"2d06",x"2458",x"ba12",x"4070",x"aca4",x"0000",x"bc00",x"0000",x"2c87",x"2458",x"b9dc",x"4070",x"aca4",x"0e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"ba02",x"4070",x"b515",x"128d",x"bc00",x"868d",x"2f35",x"24b1",x"ba03",x"4070",x"b075",x"0000",x"bc00",x"0000",x"2d42",x"24ab",x"b9dc",x"4070",x"aca4",x"0e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"b9f4",x"3d94",x"b504",x"ba04",x"8000",x"b945",x"31d8",x"3356",x"b9dc",x"3d85",x"b53c",x"ba04",x"8000",x"b945",x"31be",x"3342",x"b9dc",x"404e",x"b53c",x"ba04",x"8000",x"b945",x"31be",x"35b4"),
(x"b9f4",x"3d94",x"b0a7",x"ba28",x"b91a",x"0000",x"30f8",x"290c",x"b9dc",x"3d85",x"b032",x"ba28",x"b91a",x"0000",x"30e4",x"2973",x"b9dc",x"3d85",x"b53c",x"ba28",x"b91a",x"0000",x"31f6",x"2973"),
(x"b9f4",x"3d94",x"b0a7",x"ba1b",x"0000",x"392a",x"3165",x"3356",x"b9f4",x"4047",x"b0a7",x"ba1b",x"0000",x"392a",x"3165",x"35aa",x"b9dc",x"404e",x"b032",x"ba1b",x"0000",x"392a",x"317f",x"35b4"),
(x"ba12",x"4073",x"b00e",x"ba59",x"b87c",x"b388",x"30f7",x"2c99",x"ba09",x"4070",x"b010",x"ba44",x"b877",x"b45c",x"30f8",x"2cae",x"ba03",x"4070",x"b075",x"ba96",x"b888",x"a5cf",x"3109",x"2cb3"),
(x"b9f4",x"3d94",x"b0a7",x"bc00",x"0000",x"0000",x"301e",x"2c2f",x"b9f4",x"3d94",x"b504",x"bc00",x"0000",x"0000",x"2ea9",x"2c2f",x"b9f4",x"4047",x"b504",x"bc00",x"0000",x"0000",x"2ea8",x"3185"),
(x"b9dc",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"2b18",x"b9dc",x"3d85",x"b032",x"bc00",x"0000",x"0000",x"302e",x"2c1c",x"b9dc",x"404e",x"b032",x"bc00",x"0000",x"0000",x"302e",x"318f"),
(x"ba12",x"4076",x"b07b",x"ba77",x"b8b5",x"9fc8",x"310a",x"2c8f",x"ba03",x"4070",x"b075",x"ba96",x"b888",x"a5cf",x"3109",x"2cb3",x"ba02",x"4070",x"b515",x"ba76",x"b8b6",x"1ac2",x"3203",x"2cb3"),
(x"b9dc",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"2b18",x"b9dc",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2def",x"2b18",x"b9dc",x"3d85",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"2c1c"),
(x"b9dc",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"3073",x"31dc",x"b9dc",x"404e",x"b032",x"bc00",x"0000",x"0000",x"302e",x"318f",x"b9dc",x"404e",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"318f"),
(x"b9dc",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2def",x"2b18",x"b9dc",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2def",x"31dc",x"b9dc",x"404e",x"b53c",x"bc00",x"0000",x"0000",x"2e8c",x"318f"),
(x"ba12",x"4076",x"b522",x"ba50",x"b8e8",x"25a1",x"3207",x"2c8f",x"ba02",x"4070",x"b515",x"ba76",x"b8b6",x"1ac2",x"3203",x"2cb3",x"ba05",x"4070",x"b544",x"ba14",x"b8d9",x"337c",x"3212",x"2cb0"),
(x"b9dc",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"2cf5",x"ba12",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"2cf5",x"ba12",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"3350"),
(x"ba12",x"3d46",x"b578",x"0000",x"3c00",x"8000",x"2bc6",x"243e",x"ba12",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"243e",x"b9dc",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238"),
(x"b9dc",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"ba02",x"3d46",x"b515",x"9f10",x"3c00",x"1018",x"2b3f",x"23cc",x"ba05",x"3d46",x"b544",x"0000",x"3c00",x"8000",x"2b7e",x"23f3"),
(x"ba12",x"3d7a",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2d80",x"ba12",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2cf5",x"b9dc",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5"),
(x"b9dc",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"b9ff",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe",x"ba07",x"3d83",x"aca4",x"0000",x"8000",x"bc00",x"312d",x"2d9a"),
(x"b9f4",x"4047",x"b0a7",x"ba28",x"391a",x"0000",x"30f8",x"29e2",x"b9f4",x"4047",x"b504",x"ba28",x"391a",x"0000",x"31e3",x"29e2",x"b9dc",x"404e",x"b53c",x"ba28",x"391a",x"0000",x"31f6",x"297b"),
(x"b9dc",x"4070",x"b64e",x"11bc",x"bc00",x"8000",x"3005",x"257b",x"ba12",x"4070",x"b64e",x"11bc",x"bc00",x"8000",x"3005",x"2458",x"ba12",x"4070",x"b578",x"0e8d",x"bc00",x"868d",x"2f78",x"2458"),
(x"ba05",x"4070",x"b544",x"0cea",x"bc00",x"8a8d",x"2f54",x"249e",x"ba02",x"4070",x"b515",x"128d",x"bc00",x"868d",x"2f35",x"24b1",x"b9dc",x"4070",x"b64e",x"11bc",x"bc00",x"8000",x"3005",x"257b"),
(x"ba12",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"2af0",x"ba12",x"3154",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"280f",x"ba12",x"3cb5",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"31f0"),
(x"b9dc",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"b9ff",x"404b",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"32eb",x"b9ff",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe"),
(x"ba12",x"4057",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"330c",x"b9dc",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"ba12",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"3350"),
(x"ba02",x"404f",x"aca4",x"0000",x"8000",x"bc00",x"312a",x"32f6",x"b9ff",x"404b",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"32eb",x"b9dc",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350"),
(x"ba12",x"3d84",x"ac3b",x"b9ce",x"340f",x"b91d",x"31ea",x"3351",x"ba07",x"3d83",x"aca4",x"b9a1",x"3488",x"b935",x"31de",x"3350",x"b9ff",x"3d91",x"aca4",x"ba3a",x"1e3f",x"b904",x"31db",x"3363"),
(x"ba12",x"3d92",x"abd9",x"ba32",x"17c8",x"b90f",x"31ef",x"3364",x"b9ff",x"3d91",x"aca4",x"ba3a",x"1e3f",x"b904",x"31db",x"3363",x"b9ff",x"404b",x"aca4",x"ba32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"ba12",x"404f",x"ac0f",x"b9ea",x"b3b0",x"b908",x"31ed",x"35bd",x"ba12",x"404b",x"abe1",x"ba2a",x"96f6",x"b918",x"31ef",x"35b8",x"b9ff",x"404b",x"aca4",x"ba32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"ba12",x"3d3a",x"3523",x"ba4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"ba01",x"3d45",x"351f",x"ba5d",x"38d8",x"9f93",x"2503",x"1c77",x"ba07",x"3d45",x"3551",x"ba36",x"38b3",x"b345",x"2477",x"1cd0"),
(x"ba12",x"3d3a",x"3099",x"ba5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"ba01",x"3d45",x"307d",x"ba66",x"38cb",x"2460",x"2a6e",x"1c77",x"ba01",x"3d45",x"351f",x"ba5d",x"38d8",x"9f93",x"2503",x"1c77"),
(x"ba12",x"3d3e",x"3026",x"ba1b",x"38d7",x"3338",x"2aab",x"1e54",x"ba06",x"3d45",x"302e",x"ba14",x"38b9",x"3455",x"2aa5",x"1cb4",x"ba01",x"3d45",x"307d",x"ba66",x"38cb",x"2460",x"2a6e",x"1c77"),
(x"ba01",x"3d45",x"351f",x"a259",x"3bff",x"068d",x"2705",x"2646",x"ba01",x"3d45",x"307d",x"a418",x"3bff",x"9018",x"2b6f",x"2646",x"b9dc",x"3d46",x"2ce6",x"a067",x"3c00",x"1018",x"2c69",x"257f"),
(x"ba06",x"3d45",x"302e",x"2025",x"3bff",x"2025",x"2ba5",x"265f",x"b9dc",x"3d46",x"2ce6",x"a067",x"3c00",x"1018",x"2c69",x"257f",x"ba01",x"3d45",x"307d",x"a418",x"3bff",x"9018",x"2b6f",x"2646"),
(x"ba12",x"3d46",x"2f74",x"1ea7",x"3c00",x"1c67",x"2bf4",x"26a1",x"ba12",x"3d46",x"2ce6",x"0000",x"3c00",x"8000",x"2c69",x"26a1",x"b9dc",x"3d46",x"2ce6",x"a067",x"3c00",x"1018",x"2c69",x"257f"),
(x"ba12",x"4070",x"2f82",x"0000",x"bc00",x"0000",x"2c02",x"26b0",x"b9dc",x"4070",x"2ce6",x"0e8d",x"bc00",x"8000",x"2c74",x"27d3",x"ba12",x"4070",x"2ce6",x"0000",x"bc00",x"0000",x"2c74",x"26b0"),
(x"ba09",x"4070",x"300c",x"0000",x"bc00",x"0000",x"2bd2",x"26e2",x"ba03",x"4070",x"3071",x"0000",x"bc00",x"0000",x"2b8d",x"2702",x"b9dc",x"4070",x"2ce6",x"0e8d",x"bc00",x"8000",x"2c74",x"27d3"),
(x"b9dc",x"4070",x"2ce6",x"0e8d",x"bc00",x"8000",x"2c74",x"27d3",x"ba03",x"4070",x"3071",x"0000",x"bc00",x"0000",x"2b8d",x"2702",x"ba02",x"4070",x"3524",x"128d",x"bc00",x"068d",x"2720",x"2709"),
(x"b9f4",x"3d94",x"3513",x"ba04",x"0000",x"3945",x"31a1",x"3356",x"b9f4",x"4047",x"3513",x"ba04",x"0000",x"3945",x"31a0",x"35aa",x"b9dc",x"404e",x"354b",x"ba04",x"0000",x"3945",x"31ba",x"35b4"),
(x"b9f4",x"3d94",x"30dd",x"ba28",x"b91a",x"0000",x"31e4",x"2aa8",x"b9f4",x"3d94",x"3513",x"ba28",x"b91a",x"0000",x"30fd",x"2aa8",x"b9dc",x"3d85",x"354b",x"ba28",x"b91a",x"0000",x"30ea",x"2b0f"),
(x"b9dc",x"404e",x"3069",x"ba15",x"8000",x"b931",x"3183",x"35b4",x"b9f4",x"4047",x"30dd",x"ba15",x"8000",x"b931",x"319d",x"35aa",x"b9f4",x"3d94",x"30dd",x"ba15",x"8000",x"b931",x"319d",x"3356"),
(x"ba03",x"4070",x"3071",x"ba97",x"b888",x"25b5",x"2a77",x"20ad",x"ba09",x"4070",x"300c",x"ba44",x"b877",x"345b",x"2abd",x"2088",x"ba12",x"4073",x"300a",x"ba59",x"b87c",x"3388",x"2abf",x"1fbf"),
(x"b9f4",x"4047",x"3513",x"bc00",x"0000",x"0000",x"2aa7",x"317f",x"b9f4",x"3d94",x"3513",x"bc00",x"0000",x"0000",x"2aa7",x"2c38",x"b9f4",x"3d94",x"30dd",x"bc00",x"0000",x"0000",x"272f",x"2c38"),
(x"b9dc",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"2b2a",x"b9dc",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"31d6",x"b9dc",x"404e",x"3069",x"bc00",x"0000",x"0000",x"26a2",x"318a"),
(x"ba02",x"4070",x"3524",x"ba76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"ba03",x"4070",x"3071",x"ba97",x"b888",x"25b5",x"2a77",x"20ad",x"ba12",x"4076",x"3076",x"ba76",x"b8b6",x"1fc8",x"2a73",x"1f14"),
(x"b9dc",x"3d85",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"2c24",x"b9dc",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"2c00",x"2b2a",x"b9dc",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"2b2a"),
(x"b9dc",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2465",x"31d6",x"b9dc",x"4070",x"364e",x"bc00",x"0000",x"0000",x"2c00",x"31d6",x"b9dc",x"404e",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"318a"),
(x"b9dc",x"404e",x"354b",x"bc00",x"0000",x"0000",x"2ad8",x"318a",x"b9dc",x"4070",x"364e",x"bc00",x"0000",x"0000",x"2c00",x"31d6",x"b9dc",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"2c00",x"2b2a"),
(x"ba05",x"4070",x"3553",x"ba14",x"b8d9",x"b37c",x"2475",x"2093",x"ba02",x"4070",x"3524",x"ba76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"ba12",x"4076",x"3532",x"ba50",x"b8e8",x"a587",x"24d1",x"1f14"),
(x"b9dc",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"3138",x"2cf5",x"b9dc",x"4070",x"364e",x"0000",x"8000",x"bc00",x"3138",x"3350",x"ba12",x"4070",x"364e",x"0000",x"8000",x"bc00",x"315d",x"3350"),
(x"b9dc",x"3d46",x"364e",x"9e0a",x"3c00",x"91bc",x"2392",x"257f",x"ba12",x"3d46",x"364e",x"0000",x"3c00",x"8000",x"2392",x"26a2",x"ba12",x"3d46",x"3587",x"204d",x"3c00",x"9cb5",x"25e8",x"26a2"),
(x"ba07",x"3d45",x"3551",x"14ea",x"3c00",x"9dd6",x"267b",x"2668",x"ba01",x"3d45",x"351f",x"a259",x"3bff",x"068d",x"2705",x"2646",x"b9dc",x"3d46",x"364e",x"9e0a",x"3c00",x"91bc",x"2392",x"257f"),
(x"b9dc",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3",x"ba12",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2cc3",x"ba12",x"3d7a",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2d50"),
(x"ba08",x"3d84",x"2ce6",x"0000",x"0000",x"3c00",x"3169",x"2d69",x"ba01",x"3d90",x"2ce6",x"0000",x"0000",x"3c00",x"316e",x"2d8c",x"b9dc",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"b9dc",x"404e",x"354b",x"ba28",x"391a",x"0000",x"30ea",x"2b16",x"b9f4",x"4047",x"3513",x"ba28",x"391a",x"0000",x"30fd",x"2b7e",x"b9f4",x"4047",x"30dd",x"ba28",x"391a",x"0000",x"31e4",x"2b7e"),
(x"ba12",x"4070",x"3587",x"0e8d",x"bc00",x"0a8d",x"2613",x"26b0",x"ba12",x"4070",x"364e",x"11bc",x"bc00",x"8000",x"23e8",x"26b0",x"b9dc",x"4070",x"364e",x"11bc",x"bc00",x"8000",x"23e8",x"27d3"),
(x"b9dc",x"4070",x"364e",x"11bc",x"bc00",x"8000",x"23e8",x"27d3",x"ba02",x"4070",x"3524",x"128d",x"bc00",x"068d",x"2720",x"2709",x"ba05",x"4070",x"3553",x"10ea",x"bc00",x"068d",x"26a2",x"26f5"),
(x"ba12",x"3d84",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"32ed",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1",x"ba12",x"3d7a",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32e0"),
(x"ba12",x"3d84",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"32ed",x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"ba12",x"3d85",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"32ee",x"ba12",x"3d7a",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32e1",x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1"),
(x"ba12",x"3d92",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"32fe",x"ba12",x"404b",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"3555",x"ba12",x"3d92",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"32fe"),
(x"ba12",x"404f",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"355a",x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583",x"ba12",x"404b",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"3555"),
(x"ba12",x"404f",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"355a",x"ba12",x"404b",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"3555",x"ba12",x"404b",x"abe1",x"bc00",x"0000",x"0000",x"2c5b",x"3555"),
(x"ba12",x"3d84",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"32ed",x"ba12",x"3d85",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"32ee",x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1"),
(x"ba12",x"3d84",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"32ed",x"ba12",x"3d92",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"32fe",x"ba12",x"3d85",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"32ee"),
(x"ba12",x"3d92",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"32fe",x"ba12",x"3d92",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"32fe",x"ba12",x"3d84",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"32ed"),
(x"ba12",x"3d92",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"32fe",x"ba12",x"404b",x"abe1",x"bc00",x"0000",x"0000",x"2c5b",x"3555",x"ba12",x"404b",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"3555"),
(x"b9ff",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1",x"b9dc",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"b9dc",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"ba03",x"404f",x"2ce6",x"0000",x"0000",x"3c00",x"316c",x"32dd",x"b9dc",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"b9ff",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1"),
(x"ba12",x"4056",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"32f1",x"ba12",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"3337",x"b9dc",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337"),
(x"ba12",x"3d85",x"2c89",x"b9d0",x"342d",x"3915",x"31f9",x"3351",x"ba12",x"3d92",x"2c35",x"ba20",x"184d",x"3924",x"31f3",x"3363",x"ba01",x"3d90",x"2ce6",x"ba49",x"1ec2",x"38f2",x"3206",x"3362"),
(x"ba12",x"3d92",x"2c35",x"ba20",x"184d",x"3924",x"31f3",x"3363",x"ba12",x"404b",x"2c40",x"b9f4",x"9af6",x"3957",x"31f3",x"35b7",x"b9ff",x"404a",x"2ce6",x"ba20",x"935f",x"3925",x"3206",x"35b6"),
(x"ba12",x"404b",x"2c40",x"b9f4",x"9af6",x"3957",x"31f3",x"35b7",x"ba12",x"404e",x"2c57",x"b9db",x"b485",x"38f4",x"31f4",x"35bc",x"ba03",x"404f",x"2ce6",x"b9e5",x"b3cc",x"390b",x"3204",x"35bc"),
(x"ba05",x"3507",x"b544",x"ba14",x"38d9",x"337c",x"3214",x"2c6a",x"ba02",x"3507",x"b515",x"ba7c",x"38ae",x"1c81",x"3204",x"2c67",x"ba12",x"34dc",x"b522",x"ba50",x"38e8",x"2604",x"3209",x"2c8b"),
(x"ba02",x"3507",x"b515",x"ba7c",x"38ae",x"1c81",x"3204",x"2c67",x"ba03",x"3506",x"b075",x"baa1",x"3878",x"a594",x"310b",x"2c66",x"ba12",x"34d8",x"b07b",x"ba7d",x"38ad",x"9e59",x"310c",x"2c8b"),
(x"ba03",x"3506",x"b075",x"baa1",x"3878",x"a594",x"310b",x"2c66",x"ba09",x"3506",x"b010",x"ba5f",x"3855",x"b446",x"30f9",x"2c6a",x"ba12",x"34eb",x"b00e",x"ba6d",x"3864",x"b364",x"30f9",x"2c80"),
(x"b9dc",x"3507",x"aca4",x"9d38",x"3c00",x"8cea",x"2c87",x"224e",x"ba03",x"3506",x"b075",x"a4a8",x"3bff",x"1481",x"2d42",x"23ef",x"ba02",x"3507",x"b515",x"9f10",x"3c00",x"1018",x"2f35",x"23e3"),
(x"ba12",x"3507",x"af74",x"1f79",x"3c00",x"9c81",x"2d02",x"244a",x"b9dc",x"3507",x"aca4",x"9d38",x"3c00",x"8cea",x"2c87",x"224e",x"ba12",x"3507",x"aca4",x"0000",x"3c00",x"8000",x"2c87",x"244a"),
(x"ba09",x"3506",x"b010",x"20d0",x"3bff",x"a081",x"2d20",x"2418",x"ba03",x"3506",x"b075",x"a4a8",x"3bff",x"1481",x"2d42",x"23ef",x"b9dc",x"3507",x"aca4",x"9d38",x"3c00",x"8cea",x"2c87",x"224e"),
(x"ba09",x"3cac",x"b010",x"0000",x"bc00",x"0000",x"262a",x"247f",x"b9dc",x"3cac",x"aca4",x"0e8d",x"bc00",x"8000",x"2392",x"2570",x"ba03",x"3cac",x"b075",x"0000",x"bc00",x"0000",x"26b4",x"249f"),
(x"ba12",x"3cac",x"af8a",x"0000",x"bc00",x"0000",x"25c3",x"244d",x"ba12",x"3cac",x"aca4",x"0000",x"bc00",x"0000",x"2392",x"244d",x"b9dc",x"3cac",x"aca4",x"0e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"ba02",x"3cac",x"b515",x"128d",x"bc00",x"868d",x"2b3f",x"24a6",x"ba03",x"3cac",x"b075",x"0000",x"bc00",x"0000",x"26b4",x"249f",x"b9dc",x"3cac",x"aca4",x"0e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"b9f4",x"3c5a",x"b504",x"ba04",x"8000",x"b945",x"3140",x"3598",x"b9f4",x"3638",x"b504",x"ba04",x"8000",x"b945",x"3140",x"336f",x"b9dc",x"35ff",x"b53c",x"ba04",x"8000",x"b945",x"3127",x"335c"),
(x"b9f4",x"3638",x"b0a7",x"ba0b",x"b93d",x"0000",x"30fe",x"2bf4",x"b9dc",x"35ff",x"b032",x"ba0b",x"b93d",x"0000",x"30ea",x"2c2c",x"b9dc",x"35ff",x"b53c",x"ba0b",x"b93d",x"0000",x"31fc",x"2c2c"),
(x"b9f4",x"3c5a",x"b0a7",x"ba1b",x"0000",x"392a",x"30ec",x"3598",x"b9dc",x"3c69",x"b032",x"ba1b",x"0000",x"392a",x"3106",x"35a2",x"b9dc",x"35ff",x"b032",x"ba1b",x"0000",x"392a",x"3106",x"335c"),
(x"ba12",x"3cb3",x"b00e",x"ba59",x"b87c",x"b388",x"2447",x"2120",x"ba09",x"3cac",x"b010",x"ba44",x"b877",x"b45c",x"244b",x"21c8",x"ba03",x"3cac",x"b075",x"ba96",x"b888",x"a5cf",x"24d8",x"21ed"),
(x"b9f4",x"3638",x"b0a7",x"bc00",x"0000",x"0000",x"2ac8",x"330c",x"b9f4",x"3638",x"b504",x"bc00",x"0000",x"0000",x"26b9",x"330c",x"b9f4",x"3c5a",x"b504",x"bc00",x"0000",x"0000",x"26b9",x"3545"),
(x"b9dc",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"32d0",x"b9dc",x"35ff",x"b032",x"bc00",x"0000",x"0000",x"3036",x"331b",x"b9dc",x"3c69",x"b032",x"bc00",x"0000",x"0000",x"3036",x"354d"),
(x"ba12",x"3cb8",x"b07b",x"ba77",x"b8b5",x"9fc8",x"24df",x"20ca",x"ba03",x"3cac",x"b075",x"ba96",x"b888",x"a5cf",x"24d8",x"21ed",x"ba02",x"3cac",x"b515",x"ba76",x"b8b6",x"1ac2",x"2a51",x"21ed"),
(x"b9dc",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"32d0",x"b9dc",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2ddb",x"32d0",x"b9dc",x"35ff",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"331b"),
(x"b9dc",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"3080",x"3575",x"b9dc",x"3c69",x"b032",x"bc00",x"0000",x"0000",x"3036",x"354d",x"b9dc",x"3c69",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"354d"),
(x"b9dc",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2ddb",x"32d0",x"b9dc",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2ddb",x"3575",x"b9dc",x"3c69",x"b53c",x"bc00",x"0000",x"0000",x"2e82",x"354d"),
(x"ba12",x"3cb7",x"b522",x"ba50",x"b8e8",x"25a8",x"2a63",x"20cc",x"ba02",x"3cac",x"b515",x"ba76",x"b8b6",x"1ac2",x"2a51",x"21ed",x"ba05",x"3cac",x"b544",x"ba14",x"b8d9",x"337c",x"2a90",x"21d6"),
(x"b9dc",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"2d4a",x"ba12",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"2d4a",x"ba12",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"333a"),
(x"ba12",x"3507",x"b578",x"0000",x"3c00",x"8000",x"2f78",x"244a",x"ba12",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"244a",x"b9dc",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e"),
(x"b9dc",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"ba02",x"3507",x"b515",x"9f10",x"3c00",x"1018",x"2f35",x"23e3",x"ba05",x"3507",x"b544",x"0000",x"3c00",x"8000",x"2f54",x"2404"),
(x"ba12",x"35d5",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2dd4",x"ba12",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2d4a",x"b9dc",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"b9dc",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a",x"b9ff",x"3631",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"2e12",x"ba07",x"35fb",x"aca4",x"0000",x"8000",x"bc00",x"31fc",x"2dee"),
(x"b9f4",x"3c5a",x"b0a7",x"ba28",x"391a",x"0000",x"30fe",x"2a76",x"b9f4",x"3c5a",x"b504",x"ba28",x"391a",x"0000",x"31e9",x"2a76",x"b9dc",x"3c69",x"b53c",x"ba28",x"391a",x"0000",x"31fc",x"2a0f"),
(x"b9dc",x"3cac",x"b64e",x"11bc",x"bc00",x"8000",x"2c74",x"2570",x"ba12",x"3cac",x"b64e",x"11bc",x"bc00",x"8000",x"2c74",x"244d",x"ba12",x"3cac",x"b578",x"0e8d",x"bc00",x"8a8d",x"2bc6",x"244d"),
(x"ba05",x"3cac",x"b544",x"10ea",x"bc00",x"868d",x"2b7e",x"2492",x"ba02",x"3cac",x"b515",x"128d",x"bc00",x"868d",x"2b3f",x"24a6",x"b9dc",x"3cac",x"b64e",x"11bc",x"bc00",x"8000",x"2c74",x"2570"),
(x"b9ff",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"b9ff",x"3631",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"2e12",x"b9dc",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"ba12",x"3c7a",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"32f6",x"b9dc",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"ba12",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"333a"),
(x"ba02",x"3c6a",x"aca4",x"0000",x"8000",x"bc00",x"31f9",x"32e0",x"b9ff",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"b9dc",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a"),
(x"ba12",x"35fe",x"ac3b",x"b9ce",x"340f",x"b91d",x"3219",x"3351",x"ba07",x"35fb",x"aca4",x"b9a1",x"3488",x"b935",x"320d",x"3350",x"b9ff",x"3631",x"aca4",x"ba3a",x"1e8d",x"b905",x"320a",x"3363"),
(x"ba12",x"3635",x"abd9",x"ba32",x"1818",x"b90f",x"321e",x"3364",x"b9ff",x"3631",x"aca4",x"ba3a",x"1e8d",x"b905",x"320a",x"3363",x"b9ff",x"3c61",x"aca4",x"ba32",x"9624",x"b90f",x"320a",x"3597"),
(x"ba12",x"3c6a",x"ac0f",x"b9ea",x"b3b0",x"b908",x"321c",x"359d",x"ba12",x"3c61",x"abe1",x"ba2a",x"97c8",x"b918",x"321e",x"3597",x"b9ff",x"3c61",x"aca4",x"ba32",x"9624",x"b90f",x"320a",x"3597"),
(x"ba12",x"34db",x"3523",x"ba4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"ba01",x"3506",x"351f",x"ba5d",x"38d8",x"9f93",x"2b9a",x"1c77",x"ba07",x"3505",x"3551",x"ba36",x"38b3",x"b345",x"2b55",x"1cd0"),
(x"ba12",x"34d8",x"3099",x"ba5b",x"38da",x"1d38",x"2dba",x"1ed9",x"ba01",x"3506",x"307d",x"ba66",x"38cb",x"2460",x"2dc4",x"1c77",x"ba01",x"3506",x"351f",x"ba5d",x"38d8",x"9f93",x"2b9a",x"1c77"),
(x"ba12",x"34e8",x"3026",x"ba1b",x"38d7",x"3338",x"2de2",x"1e54",x"ba06",x"3506",x"302e",x"ba14",x"38b9",x"3455",x"2ddf",x"1cb4",x"ba01",x"3506",x"307d",x"ba66",x"38cb",x"2460",x"2dc4",x"1c77"),
(x"ba01",x"3506",x"351f",x"a259",x"3bff",x"868d",x"2d56",x"2651",x"ba01",x"3506",x"307d",x"a404",x"3bff",x"8e8d",x"2f4d",x"2652",x"b9dc",x"3507",x"2ce6",x"a067",x"3c00",x"1018",x"2fff",x"258a"),
(x"ba06",x"3506",x"302e",x"2032",x"3bff",x"2025",x"2f68",x"266a",x"b9dc",x"3507",x"2ce6",x"a067",x"3c00",x"1018",x"2fff",x"258a",x"ba01",x"3506",x"307d",x"a404",x"3bff",x"8e8d",x"2f4d",x"2652"),
(x"ba12",x"3507",x"2f74",x"1ea7",x"3c00",x"1c67",x"2f8f",x"26ad",x"ba12",x"3507",x"2ce6",x"0000",x"3c00",x"8000",x"2fff",x"26ad",x"b9dc",x"3507",x"2ce6",x"a067",x"3c00",x"1018",x"2fff",x"258a"),
(x"ba12",x"3cac",x"2f82",x"0000",x"bc00",x"0000",x"2f8d",x"26bb",x"b9dc",x"3cac",x"2ce6",x"0e8d",x"bc00",x"8000",x"2fff",x"27de",x"ba12",x"3cac",x"2ce6",x"0000",x"bc00",x"0000",x"2fff",x"26bb"),
(x"ba09",x"3cac",x"300c",x"0000",x"bc00",x"0000",x"2f73",x"26ed",x"ba03",x"3cac",x"3071",x"0000",x"bc00",x"0000",x"2f51",x"270e",x"b9dc",x"3cac",x"2ce6",x"0e8d",x"bc00",x"8000",x"2fff",x"27de"),
(x"b9dc",x"3cac",x"2ce6",x"0e8d",x"bc00",x"8000",x"2fff",x"27de",x"ba03",x"3cac",x"3071",x"0000",x"bc00",x"0000",x"2f51",x"270e",x"ba02",x"3cac",x"3524",x"128d",x"bc00",x"068d",x"2d52",x"2714"),
(x"b9dc",x"3600",x"354b",x"ba04",x"0000",x"3945",x"315d",x"335c",x"b9f4",x"3639",x"3513",x"ba04",x"0000",x"3945",x"3144",x"3370",x"b9f4",x"3c5a",x"3513",x"ba04",x"0000",x"3945",x"3144",x"3597"),
(x"b9f4",x"3639",x"30dd",x"ba0f",x"b938",x"0000",x"31e4",x"2c30",x"b9f4",x"3639",x"3513",x"ba0f",x"b938",x"0000",x"30fd",x"2c30",x"b9dc",x"3600",x"354b",x"ba0f",x"b938",x"0000",x"30ea",x"2c62"),
(x"b9f4",x"3c5a",x"30dd",x"ba15",x"8000",x"b931",x"3123",x"3597",x"b9f4",x"3639",x"30dd",x"ba15",x"8000",x"b931",x"3123",x"3370",x"b9dc",x"3600",x"3069",x"ba15",x"8000",x"b931",x"3109",x"335c"),
(x"ba03",x"3cac",x"3071",x"ba97",x"b888",x"25b5",x"2dc8",x"20ad",x"ba09",x"3cac",x"300c",x"ba44",x"b877",x"345c",x"2deb",x"2088",x"ba12",x"3cb3",x"300a",x"ba59",x"b87c",x"3388",x"2dec",x"1fbf"),
(x"b9f4",x"3c5a",x"3513",x"bc00",x"0000",x"0000",x"3028",x"3547",x"b9f4",x"3639",x"3513",x"bc00",x"0000",x"0000",x"3028",x"3323",x"b9f4",x"3639",x"30dd",x"bc00",x"0000",x"0000",x"2eaa",x"3323"),
(x"b9dc",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"32b8",x"b9dc",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"3573",x"b9dc",x"3c69",x"3069",x"bc00",x"0000",x"0000",x"2658",x"354a"),
(x"ba02",x"3cac",x"3524",x"ba76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"ba03",x"3cac",x"3071",x"ba97",x"b888",x"25b5",x"2dc8",x"20ad",x"ba12",x"3cb8",x"3076",x"ba76",x"b8b6",x"1fc8",x"2dc6",x"1f14"),
(x"b9dc",x"3600",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"3304",x"b9dc",x"3507",x"364e",x"bc00",x"0000",x"0000",x"2c23",x"32b8",x"b9dc",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"32b8"),
(x"b9dc",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"23ce",x"3573",x"b9dc",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"2c23",x"3573",x"b9dc",x"3c69",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"354a"),
(x"b9dc",x"3c69",x"354b",x"bc00",x"0000",x"0000",x"2b04",x"354a",x"b9dc",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"2c23",x"3573",x"b9dc",x"3507",x"364e",x"bc00",x"0000",x"0000",x"2c23",x"32b8"),
(x"ba05",x"3cac",x"3553",x"ba14",x"b8d9",x"b37c",x"2b54",x"2093",x"ba02",x"3cac",x"3524",x"ba76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"ba12",x"3cb7",x"3532",x"ba50",x"b8e8",x"a587",x"2b82",x"1f14"),
(x"b9dc",x"3507",x"364e",x"0000",x"8000",x"bc00",x"318d",x"2d4a",x"b9dc",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"318d",x"333a",x"ba12",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"333a"),
(x"b9dc",x"3507",x"364e",x"9e0a",x"3c00",x"91bc",x"2c87",x"258a",x"ba12",x"3507",x"364e",x"0000",x"3c00",x"8000",x"2c87",x"26ad",x"ba12",x"3507",x"3587",x"204d",x"3c00",x"9cb5",x"2d0f",x"26ad"),
(x"ba07",x"3505",x"3551",x"14ea",x"3c00",x"9dd6",x"2d34",x"2673",x"ba01",x"3506",x"351f",x"a259",x"3bff",x"868d",x"2d56",x"2651",x"b9dc",x"3507",x"364e",x"9e0a",x"3c00",x"91bc",x"2c87",x"258a"),
(x"b9dc",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a",x"ba12",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2d4a",x"ba12",x"35d7",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2dd5"),
(x"ba08",x"35fd",x"2ce6",x"0000",x"0000",x"3c00",x"31bd",x"2def",x"ba01",x"3630",x"2ce6",x"0000",x"0000",x"3c00",x"31c2",x"2e11",x"b9dc",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"b9dc",x"3c69",x"354b",x"ba28",x"391a",x"0000",x"30ea",x"2b85",x"b9f4",x"3c5a",x"3513",x"ba28",x"391a",x"0000",x"30fd",x"2bed",x"b9f4",x"3c5a",x"30dd",x"ba28",x"391a",x"0000",x"31e4",x"2bed"),
(x"ba12",x"3cac",x"3587",x"0e8d",x"bc00",x"0a8d",x"2d0f",x"26bb",x"ba12",x"3cac",x"364e",x"11bc",x"bc00",x"8000",x"2c87",x"26bb",x"b9dc",x"3cac",x"364e",x"11bc",x"bc00",x"8000",x"2c87",x"27de"),
(x"b9dc",x"3cac",x"364e",x"11bc",x"bc00",x"8000",x"2c87",x"27de",x"ba02",x"3cac",x"3524",x"128d",x"bc00",x"068d",x"2d52",x"2714",x"ba05",x"3cac",x"3553",x"10ea",x"bc00",x"068d",x"2d33",x"2701"),
(x"ba12",x"35fe",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"2c0f",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0",x"ba12",x"35d5",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2beb"),
(x"ba12",x"35fe",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"2c0f",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"ba12",x"3601",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"2c10",x"ba12",x"35d7",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2bee",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0"),
(x"ba12",x"3635",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"2c30",x"ba12",x"3c61",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"318b",x"ba12",x"3635",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"2c30"),
(x"ba12",x"3c6a",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"3195",x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3c61",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"318b"),
(x"ba12",x"3c6a",x"ac0f",x"bc00",x"0000",x"0000",x"2c56",x"3195",x"ba12",x"3c61",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"318b",x"ba12",x"3c61",x"abe1",x"bc00",x"0000",x"0000",x"2c5b",x"318b"),
(x"ba12",x"35fe",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"2c0f",x"ba12",x"3601",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"2c10",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0"),
(x"ba12",x"35fe",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"2c0f",x"ba12",x"3635",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"2c30",x"ba12",x"3601",x"2c89",x"bc00",x"0000",x"0000",x"2dbb",x"2c10"),
(x"ba12",x"3635",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"2c30",x"ba12",x"3635",x"2c35",x"bc00",x"0000",x"0000",x"2dad",x"2c30",x"ba12",x"35fe",x"ac3b",x"bc00",x"0000",x"0000",x"2c4f",x"2c0f"),
(x"ba12",x"3635",x"abd9",x"bc00",x"0000",x"0000",x"2c5c",x"2c30",x"ba12",x"3c61",x"abe1",x"bc00",x"0000",x"0000",x"2c5b",x"318b",x"ba12",x"3c61",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"318b"),
(x"b9ff",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4",x"b9dc",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"b9dc",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"ba03",x"3c69",x"2ce6",x"0000",x"0000",x"3c00",x"31c0",x"32e0",x"b9dc",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"b9ff",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4"),
(x"ba12",x"3c78",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"32f4",x"ba12",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"333a",x"b9dc",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a"),
(x"ba12",x"3601",x"2c89",x"b9d0",x"342d",x"3915",x"3227",x"3351",x"ba12",x"3635",x"2c35",x"ba20",x"1881",x"3924",x"3221",x"3363",x"ba01",x"3630",x"2ce6",x"ba49",x"1f45",x"38f2",x"3235",x"3362"),
(x"ba12",x"3635",x"2c35",x"ba20",x"1881",x"3924",x"3221",x"3363",x"ba12",x"3c61",x"2c40",x"b9f4",x"9b5f",x"3957",x"3221",x"3597",x"b9ff",x"3c60",x"2ce6",x"ba20",x"9418",x"3925",x"3234",x"3596"),
(x"ba12",x"3c61",x"2c40",x"b9f4",x"9b5f",x"3957",x"3221",x"3597",x"ba12",x"3c69",x"2c57",x"b9db",x"b485",x"38f4",x"3223",x"359c",x"ba03",x"3c69",x"2ce6",x"b9e5",x"b3cd",x"390b",x"3233",x"359c"),
(x"ba12",x"34e8",x"3026",x"bc00",x"868d",x"0000",x"2e57",x"2acb",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0",x"ba12",x"3507",x"2f74",x"bc00",x"0000",x"0000",x"2e33",x"2af0"),
(x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0"),
(x"ba12",x"34d8",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"2ab8",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0",x"ba12",x"34e8",x"3026",x"bc00",x"868d",x"0000",x"2e57",x"2acb"),
(x"ba12",x"34eb",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"2acf",x"ba12",x"3507",x"af74",x"bc00",x"0000",x"0000",x"2b94",x"2af0",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"ba12",x"34d8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"2ab8",x"ba12",x"34eb",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"2acf",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f",x"ba12",x"3507",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"2af0",x"ba12",x"34d8",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"2ab8"),
(x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c",x"ba12",x"34d8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"2ab8",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c",x"ba12",x"3507",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"2af0",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"2af0",x"ba12",x"3507",x"b578",x"bc00",x"0000",x"0000",x"25d1",x"2af0",x"ba12",x"34f4",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"2ad9"),
(x"ba12",x"34f4",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"2ad9",x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c",x"ba12",x"3507",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"2af0"),
(x"ba12",x"34d8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"2ab8",x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c",x"ba12",x"34dc",x"b522",x"bc00",x"0000",x"0000",x"26af",x"2abd"),
(x"ba12",x"34ea",x"3554",x"bc00",x"0000",x"0000",x"3039",x"2ace",x"ba12",x"3507",x"3587",x"bc00",x"0000",x"0000",x"3049",x"2af0",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"34db",x"3523",x"bc00",x"0000",x"0000",x"3029",x"2abb",x"ba12",x"34ea",x"3554",x"bc00",x"0000",x"0000",x"3039",x"2ace",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c",x"ba12",x"34f4",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"2ad9",x"ba12",x"34dc",x"b522",x"bc00",x"0000",x"0000",x"26af",x"2abd"),
(x"ba12",x"3227",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"34c4",x"ba12",x"4062",x"3753",x"2138",x"0000",x"3bff",x"39a1",x"3947",x"b940",x"4062",x"374f",x"1e73",x"9cb5",x"3c00",x"39c7",x"3946"),
(x"ba12",x"0000",x"3753",x"bc00",x"0000",x"0000",x"30de",x"1e82",x"ba12",x"0000",x"364d",x"bc00",x"0000",x"0000",x"3089",x"1e82",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f",x"ba12",x"3507",x"3587",x"bc00",x"0000",x"0000",x"3049",x"2af0",x"ba12",x"3507",x"364e",x"bc00",x"0000",x"0000",x"308a",x"2af0"),
(x"ba12",x"3507",x"364e",x"bc00",x"0000",x"0000",x"308a",x"2af0",x"ba12",x"3227",x"3753",x"bc00",x"0000",x"0000",x"30de",x"2890",x"ba12",x"3154",x"364d",x"bc00",x"0000",x"0000",x"3089",x"280f"),
(x"ba12",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"308a",x"31e6",x"ba12",x"4062",x"3753",x"bc00",x"0000",x"0000",x"30de",x"3572",x"ba12",x"3227",x"3753",x"bc00",x"0000",x"0000",x"30de",x"2890"),
(x"ba12",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"308a",x"31e6",x"ba12",x"3227",x"3753",x"bc00",x"0000",x"0000",x"30de",x"2890",x"ba12",x"3507",x"364e",x"bc00",x"0000",x"0000",x"308a",x"2af0"),
(x"ba12",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"308a",x"32a1",x"ba12",x"4070",x"364e",x"bc00",x"0000",x"0000",x"308a",x"3583",x"ba12",x"4062",x"3753",x"bc00",x"0000",x"0000",x"30de",x"3572"),
(x"ba12",x"3d3e",x"3554",x"bc00",x"0000",x"0000",x"3039",x"3298",x"ba12",x"3d46",x"3587",x"bc00",x"0000",x"0000",x"3049",x"32a1",x"ba12",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"308a",x"32a1"),
(x"ba12",x"3cb1",x"3569",x"bc00",x"0000",x"0000",x"3040",x"31ec",x"ba12",x"3d3e",x"3554",x"bc00",x"0000",x"0000",x"3039",x"3298",x"ba12",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"308a",x"32a1"),
(x"ba12",x"3cb7",x"3532",x"bc00",x"0000",x"0000",x"302e",x"31f3",x"ba12",x"3d3a",x"3523",x"bc00",x"0000",x"0000",x"3029",x"3293",x"ba12",x"3d3e",x"3554",x"bc00",x"0000",x"0000",x"3039",x"3298"),
(x"ba12",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"308a",x"31e6",x"ba12",x"3cac",x"3587",x"bc00",x"0000",x"0000",x"3049",x"31e6",x"ba12",x"3cb1",x"3569",x"bc00",x"0000",x"0000",x"3040",x"31ec"),
(x"ba12",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"308a",x"32a1",x"ba12",x"4062",x"3753",x"bc00",x"0000",x"0000",x"30de",x"3572",x"ba12",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"308a",x"31e6"),
(x"ba12",x"3d3e",x"3554",x"bc00",x"0000",x"0000",x"3039",x"3298",x"ba12",x"3cb1",x"3569",x"bc00",x"0000",x"0000",x"3040",x"31ec",x"ba12",x"3cb7",x"3532",x"bc00",x"0000",x"0000",x"302e",x"31f3"),
(x"ba12",x"3d46",x"364e",x"bc00",x"0000",x"0000",x"308a",x"32a1",x"ba12",x"3cac",x"364e",x"bc00",x"0000",x"0000",x"308a",x"31e6",x"ba12",x"3cb1",x"3569",x"bc00",x"0000",x"0000",x"3040",x"31ec"),
(x"ba12",x"3d3a",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"3293",x"ba12",x"3cb7",x"3532",x"bc00",x"0000",x"0000",x"302e",x"31f3",x"ba12",x"3cb8",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"31f4"),
(x"ba12",x"3d3a",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"3293",x"ba12",x"3d3a",x"3523",x"bc00",x"0000",x"0000",x"3029",x"3293",x"ba12",x"3cb7",x"3532",x"bc00",x"0000",x"0000",x"302e",x"31f3"),
(x"ba12",x"3cb3",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"31ee",x"ba12",x"3cac",x"2f82",x"bc00",x"0000",x"0000",x"2e36",x"31e6",x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6"),
(x"ba12",x"3d3e",x"3026",x"bc00",x"0000",x"0000",x"2e57",x"3297",x"ba12",x"3cb8",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"31f4",x"ba12",x"3cb3",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"31ee"),
(x"ba12",x"3d3e",x"3026",x"bc00",x"0000",x"0000",x"2e57",x"3297",x"ba12",x"3d3a",x"3099",x"bc00",x"0000",x"0000",x"2e7c",x"3293",x"ba12",x"3cb8",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"31f4"),
(x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1",x"ba12",x"3d46",x"2f74",x"bc00",x"0000",x"0000",x"2e33",x"32a1",x"ba12",x"3d3e",x"3026",x"bc00",x"0000",x"0000",x"2e57",x"3297"),
(x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6",x"ba12",x"3c78",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31a6",x"ba12",x"3c69",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"3194"),
(x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1",x"ba12",x"3cb3",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"31ee",x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6"),
(x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1",x"ba12",x"3d3e",x"3026",x"bc00",x"0000",x"0000",x"2e57",x"3297",x"ba12",x"3cb3",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"31ee"),
(x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1",x"ba12",x"3d46",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"32a1"),
(x"ba12",x"3d3f",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3298",x"ba12",x"3d46",x"af74",x"bc00",x"0000",x"0000",x"2b94",x"32a1",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3d3f",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3298",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"ba12",x"3cb8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"31f4",x"ba12",x"3d3a",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"3293",x"ba12",x"3d3f",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3298"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3c69",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"3194",x"ba12",x"3c61",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"318b"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6",x"ba12",x"3c69",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"3194"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3cac",x"af8a",x"bc00",x"0000",x"0000",x"2b8d",x"31e6",x"ba12",x"3cb3",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"31ee"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3d46",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"32a1",x"ba12",x"3cac",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"31e6"),
(x"ba12",x"3cb3",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"31ee",x"ba12",x"3cb8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"31f4",x"ba12",x"3d3f",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3298"),
(x"ba12",x"3cac",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"31e6",x"ba12",x"3cb3",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"31ee",x"ba12",x"3d3f",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3298"),
(x"ba12",x"3cb7",x"b522",x"bc00",x"0000",x"0000",x"26af",x"31f3",x"ba12",x"3d3b",x"b522",x"bc00",x"0000",x"0000",x"26af",x"3294",x"ba12",x"3d3a",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"3293"),
(x"ba12",x"3cb7",x"b522",x"bc00",x"0000",x"0000",x"26af",x"31f3",x"ba12",x"3d3a",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"3293",x"ba12",x"3cb8",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"31f4"),
(x"ba12",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"32a1",x"ba12",x"3d46",x"b578",x"bc00",x"0000",x"0000",x"25d1",x"32a1",x"ba12",x"3d41",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"329b"),
(x"ba12",x"3cb1",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"31ec",x"ba12",x"3d3b",x"b522",x"bc00",x"0000",x"0000",x"26af",x"3294",x"ba12",x"3cb7",x"b522",x"bc00",x"0000",x"0000",x"26af",x"31f3"),
(x"ba12",x"3cb1",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"31ec",x"ba12",x"3d41",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"329b",x"ba12",x"3d3b",x"b522",x"bc00",x"0000",x"0000",x"26af",x"3294"),
(x"ba12",x"3cb1",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"31ec",x"ba12",x"3cac",x"b578",x"bc00",x"0000",x"0000",x"25d1",x"31e6",x"ba12",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"31e6"),
(x"ba12",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"31e6",x"ba12",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"32a1",x"ba12",x"3d41",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"329b"),
(x"ba12",x"8000",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"1e82",x"ba12",x"3154",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"280f",x"ba12",x"314f",x"b64f",x"bc00",x"0000",x"0000",x"234a",x"280c"),
(x"ba12",x"408e",x"3753",x"bc00",x"0000",x"0000",x"30de",x"35a7",x"ba12",x"4062",x"3753",x"bc00",x"0000",x"0000",x"30de",x"3572",x"ba12",x"4070",x"364e",x"bc00",x"0000",x"0000",x"308a",x"3583"),
(x"ba12",x"4073",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"3586",x"ba12",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"3583",x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7"),
(x"ba12",x"4073",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"3586",x"ba12",x"4070",x"b578",x"bc00",x"0000",x"0000",x"25d1",x"3583",x"ba12",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"3583"),
(x"ba12",x"4073",x"3569",x"bc00",x"0000",x"0000",x"3040",x"3586",x"ba12",x"4070",x"364e",x"bc00",x"0000",x"0000",x"308a",x"3583",x"ba12",x"4070",x"3587",x"bc00",x"0000",x"0000",x"3049",x"3583"),
(x"ba12",x"4073",x"3569",x"bc00",x"0000",x"0000",x"3040",x"3586",x"ba12",x"408e",x"3753",x"bc00",x"0000",x"0000",x"30de",x"35a7",x"ba12",x"4070",x"364e",x"bc00",x"0000",x"0000",x"308a",x"3583"),
(x"ba12",x"4076",x"b522",x"bc00",x"0000",x"0000",x"26af",x"3589",x"ba12",x"4073",x"b55a",x"bc00",x"0000",x"0000",x"261e",x"3586",x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7"),
(x"ba12",x"4076",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"358a",x"ba12",x"4076",x"b522",x"bc00",x"0000",x"0000",x"26af",x"3589",x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7"),
(x"ba12",x"408e",x"3753",x"bc00",x"0000",x"0000",x"30de",x"35a7",x"ba12",x"4073",x"3569",x"bc00",x"0000",x"0000",x"3040",x"3586",x"ba12",x"4076",x"3532",x"bc00",x"0000",x"0000",x"302e",x"3589"),
(x"ba12",x"408e",x"3753",x"bc00",x"0000",x"0000",x"30de",x"35a7",x"ba12",x"4076",x"3532",x"bc00",x"0000",x"0000",x"302e",x"3589",x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a"),
(x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a",x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7",x"ba12",x"408e",x"3753",x"bc00",x"0000",x"0000",x"30de",x"35a7"),
(x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a",x"ba12",x"4076",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"358a",x"ba12",x"408e",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"35a7"),
(x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583",x"ba12",x"4070",x"af8a",x"bc00",x"0000",x"0000",x"2b8d",x"3583",x"ba12",x"4073",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3587"),
(x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583",x"ba12",x"4073",x"b00e",x"bc00",x"0000",x"0000",x"2b5d",x"3587",x"ba12",x"4076",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"358a"),
(x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583",x"ba12",x"4076",x"b07b",x"bc00",x"0000",x"0000",x"2b17",x"358a",x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a"),
(x"ba12",x"404e",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"355a",x"ba12",x"404b",x"2c40",x"bc00",x"0000",x"0000",x"2daf",x"3555",x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583"),
(x"ba12",x"4073",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"3587",x"ba12",x"4070",x"2f82",x"bc00",x"0000",x"0000",x"2e36",x"3583",x"ba12",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3583"),
(x"ba12",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3583",x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a",x"ba12",x"4073",x"300a",x"bc00",x"0000",x"0000",x"2e4d",x"3587"),
(x"ba12",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3583",x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583",x"ba12",x"4076",x"3076",x"bc00",x"0000",x"0000",x"2e71",x"358a"),
(x"ba12",x"4070",x"2ce6",x"bc00",x"0000",x"0000",x"2dca",x"3583",x"ba12",x"404e",x"2c57",x"bc00",x"0000",x"0000",x"2db3",x"355a",x"ba12",x"4070",x"aca4",x"bc00",x"0000",x"0000",x"2c3e",x"3583"),
(x"b9b7",x"314b",x"b64f",x"9e3f",x"bc00",x"1418",x"38da",x"3917",x"ba12",x"314f",x"b64f",x"a24c",x"bbff",x"11bc",x"38be",x"3917",x"ba12",x"3154",x"364d",x"9e3f",x"bc00",x"1418",x"38be",x"39de"),
(x"b9b7",x"314b",x"b64f",x"0000",x"0000",x"3c00",x"396a",x"3402",x"b941",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"397d",x"3342",x"ba12",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"395b",x"3342"),
(x"3a12",x"4092",x"b6b0",x"0000",x"8a8d",x"bc00",x"3aed",x"3881",x"b941",x"4092",x"b6b0",x"0000",x"8a8d",x"bc00",x"39fa",x"3881",x"b941",x"3d3f",x"b6b0",x"0000",x"8a8d",x"bc00",x"39fa",x"3929"),
(x"ba12",x"4070",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"3583",x"ba12",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"32a1",x"ba12",x"3d42",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"329d"),
(x"ba12",x"3154",x"b751",x"1018",x"8000",x"bc00",x"3bbf",x"355b",x"ba12",x"8000",x"b751",x"1018",x"8000",x"bc00",x"3bbf",x"34f7",x"b941",x"34e4",x"b751",x"0e8d",x"8000",x"bc00",x"3ba1",x"35af"),
(x"b941",x"34e4",x"b751",x"0e8d",x"8000",x"bc00",x"3ba1",x"35af",x"ba12",x"3cb5",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"37bc",x"ba12",x"3154",x"b751",x"1018",x"8000",x"bc00",x"3bbf",x"355b"),
(x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929",x"ba12",x"3d42",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"3807",x"b941",x"3d3f",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"3807"),
(x"b941",x"3d3f",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"3807",x"ba12",x"3d42",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"3807",x"ba12",x"3cb5",x"b751",x"0cea",x"8000",x"bc00",x"3bbf",x"37bc"),
(x"ba12",x"3d46",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"32a1",x"ba12",x"3cac",x"b64e",x"bc00",x"0000",x"0000",x"2351",x"31e6",x"ba12",x"3cb5",x"b751",x"bc00",x"0000",x"0000",x"1c22",x"31f0"),
(x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af",x"b941",x"34e4",x"b751",x"0e8d",x"8000",x"bc00",x"3ba1",x"35af",x"b941",x"3161",x"b751",x"0cea",x"8000",x"bc00",x"3ba1",x"355c"),
(x"b941",x"34e4",x"b6b0",x"3c00",x"0000",x"0000",x"3b75",x"380d",x"b941",x"3cb4",x"b6af",x"3c00",x"0000",x"0000",x"3b75",x"3926",x"b941",x"3cb4",x"b751",x"3c00",x"0000",x"0000",x"3b80",x"3926"),
(x"b941",x"4092",x"b6b0",x"3c00",x"0000",x"0000",x"3b84",x"391f",x"b941",x"4092",x"b751",x"3c00",x"0000",x"0000",x"3b8e",x"391f",x"b941",x"3d3f",x"b751",x"3c00",x"0000",x"0000",x"3b8e",x"3813"),
(x"ba77",x"40a6",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3938",x"ba77",x"40a4",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3936",x"ba73",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3935"),
(x"ba4d",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"393b",x"ba72",x"40a7",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3938",x"ba73",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"3bce",x"3935"),
(x"ba4b",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba4b",x"409a",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba4a",x"4099",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3930"),
(x"ba49",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba4b",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba47",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc7",x"392f"),
(x"ba4d",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"393b",x"ba49",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"3bc8",x"3931",x"ba30",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc4",x"392f"),
(x"ba29",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"393f",x"ba30",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"3bc4",x"392f",x"ba27",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392e"),
(x"ba26",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"3bc2",x"392c",x"ba29",x"4091",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392b",x"ba27",x"408f",x"b74a",x"0000",x"8000",x"bc00",x"3bc3",x"392a"),
(x"ba21",x"4092",x"b74a",x"b299",x"a65f",x"bbd3",x"3bc2",x"392c",x"ba26",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"3bc2",x"392c",x"ba1f",x"408e",x"b74a",x"b075",x"a386",x"bbeb",x"3bc1",x"3929"),
(x"ba1e",x"40b8",x"b74a",x"9418",x"257a",x"bbff",x"3bc1",x"3942",x"ba22",x"4094",x"b74a",x"b0ee",x"1881",x"bbe7",x"3bc2",x"392d",x"ba12",x"408e",x"b751",x"90ea",x"128d",x"bc00",x"3bbf",x"3929"),
(x"b940",x"4062",x"364d",x"3c00",x"0000",x"0000",x"393e",x"346c",x"b940",x"0000",x"364d",x"3c00",x"0000",x"0000",x"393e",x"3888",x"b940",x"0000",x"374f",x"3c00",x"0000",x"0000",x"394f",x"3888"),
(x"b9b6",x"3154",x"364d",x"1818",x"8000",x"bc00",x"393a",x"3464",x"b940",x"4062",x"364d",x"0a8d",x"068d",x"bc00",x"3928",x"383c",x"b9b7",x"40b6",x"364d",x"068d",x"0000",x"bc00",x"393a",x"3867"),
(x"b9b6",x"3154",x"364d",x"1818",x"8000",x"bc00",x"393a",x"3464",x"b940",x"0000",x"364d",x"1a8d",x"8000",x"bc00",x"3929",x"340e",x"b940",x"4062",x"364d",x"0a8d",x"068d",x"bc00",x"3928",x"383c"),
(x"b9b7",x"40b6",x"b64d",x"3c00",x"0cea",x"8a8d",x"1ca6",x"38e0",x"b9b7",x"314b",x"b64f",x"3c00",x"8000",x"9418",x"1ca0",x"3aac",x"b9b6",x"3154",x"364d",x"3c00",x"0a8d",x"8e8d",x"2d77",x"3aac"),
(x"b9b7",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"396a",x"3887",x"b941",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"397d",x"3887",x"b941",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404"),
(x"ba12",x"0000",x"364d",x"1624",x"8e8d",x"bc00",x"3948",x"340e",x"b9b6",x"3154",x"364d",x"175f",x"8000",x"bc00",x"393a",x"3464",x"ba12",x"3154",x"364d",x"0000",x"8000",x"bc00",x"3948",x"3464"),
(x"b941",x"40b6",x"b694",x"3c00",x"0000",x"0000",x"38b9",x"3bef",x"b941",x"3161",x"b694",x"3c00",x"0000",x"0000",x"38a5",x"3980",x"b941",x"3161",x"b64f",x"3c00",x"0000",x"0000",x"389d",x"3981"),
(x"b941",x"8000",x"b751",x"3c00",x"8000",x"868d",x"38b5",x"3912",x"b941",x"8000",x"b64f",x"3c00",x"8000",x"868d",x"3899",x"3914",x"b941",x"3161",x"b694",x"3c00",x"0000",x"0000",x"38a5",x"3980"),
(x"b9c7",x"3527",x"b696",x"0000",x"3c00",x"8000",x"2de7",x"3ab7",x"3a98",x"3527",x"b696",x"0000",x"3c00",x"8000",x"2de7",x"3bfc",x"3a98",x"3527",x"364c",x"0000",x"3c00",x"8000",x"3199",x"3bfc"),
(x"3a94",x"3488",x"3650",x"0000",x"bc00",x"0000",x"3af7",x"37a8",x"3a94",x"3488",x"b696",x"0000",x"bc00",x"0000",x"3b42",x"37a8",x"b9cb",x"3488",x"b696",x"0000",x"bc00",x"0000",x"3b42",x"3689"),
(x"3a94",x"3488",x"3650",x"0000",x"2631",x"3bff",x"3976",x"39c4",x"b9cb",x"3488",x"3650",x"0000",x"2631",x"3bff",x"3976",x"3b5b",x"b9c7",x"3527",x"364c",x"0000",x"2631",x"3bff",x"398a",x"3b5b"),
(x"b944",x"3499",x"3748",x"0000",x"34bc",x"3ba4",x"393c",x"3b5b",x"b944",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3b5b",x"3a1c",x"34b8",x"372f",x"0000",x"3bf0",x"2ff1",x"3946",x"3a40"),
(x"b944",x"345f",x"3745",x"0000",x"ba15",x"3932",x"3929",x"3b5b",x"3a1c",x"345f",x"3745",x"8000",x"b970",x"39dd",x"3929",x"3a40",x"3a1c",x"3449",x"3727",x"0000",x"ba5c",x"38da",x"3920",x"3a40"),
(x"3aef",x"40b8",x"376a",x"3b44",x"36ae",x"0000",x"3718",x"3ab8",x"3aef",x"40b8",x"b74a",x"3b44",x"36ae",x"0000",x"3718",x"3910",x"3af9",x"40b3",x"b74a",x"3a61",x"38d2",x"0000",x"370a",x"3910"),
(x"ba1e",x"40b8",x"376a",x"0000",x"3587",x"3b81",x"36a6",x"3ab2",x"3aef",x"40b8",x"376a",x"0000",x"3587",x"3b81",x"36a6",x"3868",x"3af9",x"40b3",x"377b",x"8000",x"38b6",x"3a76",x"3692",x"3863"),
(x"3b1e",x"40ab",x"37c7",x"8000",x"3a96",x"388a",x"367e",x"385b",x"ba4d",x"40ab",x"37c7",x"0000",x"3af8",x"37d8",x"367f",x"3abe",x"ba29",x"40b3",x"377b",x"8000",x"39b1",x"399e",x"3692",x"3ab6"),
(x"3b43",x"40a7",x"3805",x"0000",x"3b38",x"36e2",x"366b",x"3852",x"ba72",x"40a7",x"3805",x"8000",x"3ae3",x"3811",x"366b",x"3ac9",x"ba4d",x"40ab",x"37c7",x"0000",x"3af8",x"37d8",x"367f",x"3abe"),
(x"3b48",x"40a6",x"380b",x"0000",x"3824",x"3ad7",x"3656",x"384c",x"ba77",x"40a6",x"380b",x"0000",x"34ea",x"3b9c",x"3656",x"3ad1",x"ba72",x"40a7",x"3805",x"8000",x"3ae3",x"3811",x"366b",x"3ac9"),
(x"3b48",x"40a4",x"380c",x"0000",x"b0b3",x"3be9",x"3642",x"384c",x"ba77",x"40a4",x"380c",x"0000",x"b607",x"3b69",x"3641",x"3ad1",x"ba77",x"40a6",x"380b",x"0000",x"34ea",x"3b9c",x"3656",x"3ad1"),
(x"3b44",x"40a2",x"3807",x"8000",x"ba4c",x"38ee",x"362d",x"3853",x"ba73",x"40a2",x"3807",x"0000",x"ba9a",x"3884",x"362d",x"3acb",x"ba77",x"40a4",x"380c",x"0000",x"b607",x"3b69",x"3641",x"3ad1"),
(x"3b1a",x"409b",x"37ba",x"0000",x"baba",x"3854",x"3619",x"385c",x"ba49",x"409b",x"37ba",x"0000",x"baba",x"3854",x"361a",x"3ac3",x"ba73",x"40a2",x"3807",x"0000",x"ba9a",x"3884",x"362d",x"3acb"),
(x"3b1c",x"409b",x"37bd",x"8000",x"3873",x"3aa5",x"37b7",x"3971",x"ba4b",x"409b",x"37bd",x"0000",x"384b",x"3abf",x"37b7",x"3ad1",x"ba49",x"409b",x"37ba",x"0000",x"3897",x"3a8d",x"37c2",x"3ace"),
(x"3b1c",x"409a",x"37c0",x"0000",x"32ec",x"3bcf",x"37ac",x"3971",x"ba4b",x"409a",x"37c0",x"8000",x"8cea",x"3c00",x"37ac",x"3ad1",x"ba4b",x"409b",x"37bd",x"0000",x"384b",x"3abf",x"37b7",x"3ad1"),
(x"3b1b",x"4099",x"37bf",x"0000",x"b654",x"3b58",x"37a1",x"3972",x"ba4a",x"4099",x"37bf",x"8000",x"b927",x"3a1e",x"37a1",x"3ad1",x"ba4b",x"409a",x"37c0",x"8000",x"8cea",x"3c00",x"37ac",x"3ad1"),
(x"3b18",x"4098",x"37b7",x"0000",x"bbda",x"3211",x"3795",x"3976",x"ba47",x"4098",x"37b7",x"8000",x"bbf8",x"2d73",x"3795",x"3acd",x"ba4a",x"4099",x"37bf",x"8000",x"b927",x"3a1e",x"37a1",x"3ad1"),
(x"3b01",x"4098",x"3785",x"0000",x"bbfe",x"28cc",x"378a",x"397c",x"ba30",x"4098",x"3785",x"0000",x"bbfe",x"28cc",x"378b",x"3ac9",x"ba47",x"4098",x"37b7",x"8000",x"bbf8",x"2d73",x"3795",x"3acd"),
(x"3af8",x"4096",x"3773",x"0000",x"b9da",x"3973",x"3809",x"394c",x"ba27",x"4096",x"3773",x"8000",x"b967",x"39e6",x"3809",x"3ad2",x"ba30",x"4098",x"3785",x"0000",x"ba3a",x"3905",x"380f",x"3ad7"),
(x"3af3",x"4094",x"3767",x"8000",x"b745",x"3b20",x"3802",x"3950",x"ba22",x"4094",x"3767",x"8000",x"b449",x"3bb5",x"3802",x"3acf",x"ba27",x"4096",x"3773",x"8000",x"b967",x"39e6",x"3809",x"3ad2"),
(x"3af1",x"4092",x"3766",x"0000",x"ac55",x"3bfb",x"37f9",x"3951",x"ba21",x"4092",x"3766",x"0000",x"ac55",x"3bfb",x"37f9",x"3ace",x"ba22",x"4094",x"3767",x"8000",x"b449",x"3bb5",x"3802",x"3acf"),
(x"3af6",x"4092",x"3775",x"0000",x"3ba1",x"34ce",x"37ee",x"3983",x"ba26",x"4092",x"3775",x"8000",x"3a53",x"38e6",x"37ee",x"3acc",x"ba21",x"4092",x"3766",x"0000",x"3bf8",x"2d9e",x"37f8",x"3ac8"),
(x"3afa",x"4091",x"3778",x"0000",x"326d",x"3bd6",x"37e3",x"397e",x"ba29",x"4091",x"3778",x"0000",x"26d5",x"3bff",x"37e3",x"3ad1",x"ba26",x"4092",x"3775",x"8000",x"3a53",x"38e6",x"37ee",x"3acc"),
(x"3af8",x"408f",x"3777",x"8000",x"b682",x"3b4e",x"37d8",x"3980",x"ba27",x"408f",x"3777",x"0000",x"b8ed",x"3a4d",x"37d8",x"3acf",x"ba29",x"4091",x"3778",x"0000",x"26d5",x"3bff",x"37e3",x"3ad1"),
(x"3af0",x"408e",x"3769",x"8000",x"bb26",x"372c",x"37cd",x"3985",x"ba1f",x"408e",x"3769",x"0000",x"bbd1",x"32c7",x"37cd",x"3aca",x"ba27",x"408f",x"3777",x"0000",x"b8ed",x"3a4d",x"37d8",x"3acf"),
(x"3af8",x"4096",x"b74a",x"3a2e",x"b913",x"0000",x"382d",x"3888",x"3af3",x"4094",x"b74a",x"3ba9",x"b498",x"0000",x"3829",x"3888",x"3af3",x"4094",x"3767",x"3b41",x"b6be",x"8000",x"3829",x"39a6"),
(x"3b48",x"40a4",x"b74a",x"3b97",x"b50b",x"8000",x"36c9",x"3910",x"3b44",x"40a2",x"b74a",x"3892",x"ba90",x"068d",x"36bb",x"3910",x"3b44",x"40a2",x"3807",x"38f8",x"ba45",x"0000",x"36ba",x"3acd"),
(x"3b01",x"4098",x"b74a",x"391e",x"ba25",x"0000",x"3832",x"3888",x"3af8",x"4096",x"b74a",x"3a2e",x"b913",x"0000",x"382d",x"3888",x"3af8",x"4096",x"3773",x"39a4",x"b9ac",x"0000",x"382d",x"39a9"),
(x"3af0",x"408e",x"b74a",x"31b5",x"bbdf",x"0000",x"3813",x"38cb",x"3ae3",x"408e",x"b751",x"0000",x"bc00",x"0000",x"380f",x"38cb",x"3ae3",x"408e",x"3753",x"0000",x"bc00",x"0000",x"380f",x"39c7"),
(x"3b48",x"40a6",x"380b",x"3bc1",x"33d8",x"8000",x"36d8",x"3ad0",x"3b48",x"40a6",x"b74a",x"3af6",x"37df",x"0000",x"36d8",x"3910",x"3b48",x"40a4",x"b74a",x"3b97",x"b50b",x"8000",x"36c9",x"3910"),
(x"3b18",x"4098",x"b74a",x"2dde",x"bbf7",x"8000",x"3793",x"3872",x"3b01",x"4098",x"b74a",x"2918",x"bbfe",x"0000",x"378b",x"3872",x"3b01",x"4098",x"3785",x"2918",x"bbfe",x"0000",x"378b",x"3968"),
(x"3af8",x"408f",x"b74a",x"399f",x"b9b0",x"068d",x"3817",x"38cc",x"3af0",x"408e",x"b74a",x"31b5",x"bbdf",x"0000",x"3813",x"38cb",x"3af0",x"408e",x"3769",x"361a",x"bb65",x"8000",x"3813",x"39ca"),
(x"3b43",x"40a7",x"3805",x"37c0",x"3aff",x"8000",x"36e6",x"3acb",x"3b43",x"40a7",x"b74a",x"3671",x"3b52",x"0000",x"36e6",x"3910",x"3b48",x"40a6",x"b74a",x"3af6",x"37df",x"0000",x"36d8",x"3910"),
(x"3b1b",x"4099",x"b74a",x"3aa8",x"b86e",x"0000",x"379b",x"3872",x"3b18",x"4098",x"b74a",x"2dde",x"bbf7",x"8000",x"3793",x"3872",x"3b18",x"4098",x"37b7",x"32b5",x"bbd2",x"0000",x"3793",x"396c"),
(x"3afa",x"4091",x"b74a",x"3bdb",x"31fa",x"8000",x"381b",x"38cc",x"3af8",x"408f",x"b74a",x"399f",x"b9b0",x"068d",x"3817",x"38cc",x"3af8",x"408f",x"3777",x"3ac3",x"b845",x"0000",x"3817",x"39cd"),
(x"3b1e",x"40ab",x"37c7",x"379e",x"3b08",x"0000",x"36f6",x"3ac3",x"3b1e",x"40ab",x"b74a",x"3890",x"3a91",x"8000",x"36f6",x"3910",x"3b43",x"40a7",x"b74a",x"3671",x"3b52",x"0000",x"36e6",x"3910"),
(x"3b1c",x"409a",x"b74a",x"3bfc",x"abd5",x"8000",x"37a3",x"3873",x"3b1b",x"4099",x"b74a",x"3aa8",x"b86e",x"0000",x"379b",x"3872",x"3b1b",x"4099",x"37bf",x"3b8d",x"b548",x"8000",x"379b",x"3970"),
(x"3af6",x"4092",x"3775",x"38a6",x"3a82",x"0000",x"381f",x"39cc",x"3af6",x"4092",x"b74a",x"35d6",x"3b72",x"0000",x"3820",x"38cc",x"3afa",x"4091",x"b74a",x"3bdb",x"31fa",x"8000",x"381b",x"38cc"),
(x"3af9",x"40b3",x"377b",x"39af",x"39a0",x"8000",x"370a",x"3aba",x"3af9",x"40b3",x"b74a",x"3a61",x"38d2",x"0000",x"370a",x"3910",x"3b1e",x"40ab",x"b74a",x"3890",x"3a91",x"8000",x"36f6",x"3910"),
(x"3b1c",x"409b",x"37bd",x"3bb8",x"3431",x"8000",x"37ab",x"396e",x"3b1c",x"409b",x"b74a",x"3b4e",x"3681",x"0000",x"37ab",x"3873",x"3b1c",x"409a",x"b74a",x"3bfc",x"abd5",x"8000",x"37a3",x"3873"),
(x"3af1",x"4092",x"3766",x"3033",x"3bee",x"0000",x"3824",x"39c5",x"3af1",x"4092",x"b74a",x"3033",x"3bee",x"0000",x"3824",x"38cc",x"3af6",x"4092",x"b74a",x"35d6",x"3b72",x"0000",x"3820",x"38cc"),
(x"3b1a",x"409b",x"37ba",x"3ad7",x"3825",x"0000",x"37b3",x"396b",x"3b1a",x"409b",x"b74a",x"3ad7",x"3825",x"0000",x"37b3",x"3872",x"3b1c",x"409b",x"b74a",x"3b4e",x"3681",x"0000",x"37ab",x"3873"),
(x"3af3",x"4094",x"b74a",x"3ba9",x"b498",x"0000",x"3829",x"3888",x"3af1",x"4092",x"b74a",x"3be9",x"b0c2",x"0000",x"3824",x"3888",x"3af1",x"4092",x"3766",x"3be9",x"b0c2",x"0000",x"3824",x"39a5"),
(x"3b44",x"40a2",x"b74a",x"3892",x"ba90",x"068d",x"36bb",x"3910",x"3b1a",x"409b",x"b74a",x"3863",x"bab0",x"0000",x"36a6",x"3910",x"3b1a",x"409b",x"37ba",x"3863",x"bab0",x"0000",x"36a6",x"3ac4"),
(x"3ae3",x"408e",x"3753",x"0000",x"bc00",x"0000",x"37c3",x"398c",x"ba12",x"408e",x"3753",x"0000",x"bc00",x"868d",x"37c3",x"3ac4",x"ba1f",x"408e",x"3769",x"0000",x"bbd1",x"32c7",x"37cd",x"3aca"),
(x"3ae3",x"3227",x"3753",x"a138",x"0000",x"3bff",x"3bf9",x"34c4",x"3a11",x"0000",x"374f",x"a138",x"0000",x"3bff",x"3bd3",x"3436",x"3a11",x"4062",x"374f",x"a018",x"9953",x"3c00",x"3bd3",x"3946"),
(x"3a88",x"314b",x"b64f",x"1e3f",x"bc00",x"1418",x"38db",x"3917",x"3a87",x"3154",x"364d",x"0000",x"bc00",x"15bc",x"38db",x"39de",x"3ae3",x"3154",x"364d",x"1e3f",x"bc00",x"1418",x"38f7",x"39de"),
(x"3ae3",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"399f",x"3342",x"3a12",x"8000",x"b64f",x"0000",x"0000",x"3c00",x"397d",x"3342",x"3a88",x"314b",x"b64f",x"0000",x"868d",x"3c00",x"3990",x"3402"),
(x"b941",x"3cb4",x"b6af",x"0000",x"bc00",x"0000",x"39d2",x"34a6",x"3a12",x"3cb4",x"b6af",x"0000",x"bc00",x"0000",x"3bc8",x"34a6",x"3a12",x"3cb4",x"b751",x"0000",x"bc00",x"0000",x"3bc8",x"3494"),
(x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807",x"b941",x"3d3f",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"3807",x"b941",x"3cb4",x"b751",x"0a8d",x"8000",x"bc00",x"3ba1",x"37bb"),
(x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af",x"3ae3",x"8000",x"b751",x"8a8d",x"0a8d",x"bc00",x"39d8",x"34f7",x"3ae3",x"3154",x"b751",x"9018",x"8000",x"bc00",x"39d8",x"355b"),
(x"3ae3",x"3cb5",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"37bc",x"3a12",x"3cb4",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"37bb",x"3a12",x"34e4",x"b751",x"8e8d",x"8000",x"bc00",x"39f6",x"35af"),
(x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3a12",x"4092",x"b751",x"068d",x"21e3",x"bbff",x"39f6",x"392c",x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807"),
(x"3ae3",x"3cb5",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"37bc",x"3ae3",x"3d42",x"b751",x"8cea",x"8000",x"bc00",x"39d8",x"3807",x"3a12",x"3d3f",x"b751",x"8a8d",x"8000",x"bc00",x"39f6",x"3807"),
(x"3a12",x"34e4",x"b6b0",x"0000",x"3c00",x"8000",x"3bc8",x"34a6",x"b941",x"34e4",x"b6b0",x"0000",x"3c00",x"8000",x"39d2",x"34a6",x"b941",x"34e4",x"b751",x"0000",x"3c00",x"8000",x"39d2",x"34b8"),
(x"3a12",x"3cb4",x"b751",x"bc00",x"0000",x"0000",x"3b69",x"3926",x"3a12",x"3cb4",x"b6af",x"bc00",x"0000",x"0000",x"3b75",x"3926",x"3a12",x"34e4",x"b6b0",x"bc00",x"0000",x"0000",x"3b75",x"380d"),
(x"3a12",x"4092",x"b6b0",x"bc00",x"0000",x"0000",x"3b9e",x"3922",x"3a12",x"3d3f",x"b6b0",x"bc00",x"0000",x"0000",x"3b9e",x"3814",x"3a12",x"3d3f",x"b751",x"bc00",x"0000",x"0000",x"3b90",x"3814"),
(x"3a12",x"4092",x"b6b0",x"0000",x"bc00",x"0000",x"3bcd",x"3475",x"3a12",x"4092",x"b751",x"0000",x"bc00",x"0000",x"3bcd",x"345e",x"b941",x"4092",x"b751",x"0000",x"bc00",x"0000",x"39ce",x"345e"),
(x"b940",x"4062",x"374f",x"1e73",x"9cb5",x"3c00",x"39c7",x"3946",x"ba12",x"408e",x"3753",x"10ea",x"a1e3",x"3bff",x"39a1",x"3966",x"3ae3",x"408e",x"3753",x"8cea",x"a1fd",x"3bff",x"3bf9",x"3966"),
(x"3b48",x"40a6",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3938",x"3b43",x"40a7",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3938",x"3b44",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3935"),
(x"3b44",x"40a2",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3935",x"3b43",x"40a7",x"b74a",x"0000",x"8000",x"bc00",x"39c9",x"3938",x"3b1e",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"393b"),
(x"3b1b",x"4099",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3930",x"3b1c",x"409a",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3931",x"3b1c",x"409b",x"b74a",x"068d",x"0000",x"bc00",x"39cf",x"3931"),
(x"3b18",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d0",x"392f",x"3b1c",x"409b",x"b74a",x"068d",x"0000",x"bc00",x"39cf",x"3931",x"3b1a",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3931"),
(x"3b01",x"4098",x"b74a",x"0000",x"8000",x"bc00",x"39d3",x"392f",x"3b1a",x"409b",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"3931",x"3b1e",x"40ab",x"b74a",x"0000",x"8000",x"bc00",x"39cf",x"393b"),
(x"3af9",x"40b3",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"393f",x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942",x"3af8",x"4096",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392e"),
(x"3af8",x"408f",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392a",x"3afa",x"4091",x"b74a",x"0000",x"8000",x"bc00",x"39d4",x"392b",x"3af6",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"39d5",x"392c"),
(x"3af0",x"408e",x"b74a",x"3075",x"a386",x"bbeb",x"39d6",x"3929",x"3af6",x"4092",x"b74a",x"0000",x"8000",x"bc00",x"39d5",x"392c",x"3af1",x"4092",x"b74a",x"3299",x"a666",x"bbd3",x"39d5",x"392c"),
(x"3ae3",x"408e",x"b751",x"10ea",x"128d",x"bc00",x"39d8",x"3929",x"3af3",x"4094",x"b74a",x"30ed",x"1881",x"bbe7",x"39d5",x"392d",x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942"),
(x"3aef",x"40b8",x"376a",x"0000",x"3c00",x"8000",x"316c",x"38f0",x"ba1e",x"40b8",x"376a",x"0000",x"3c00",x"8000",x"316c",x"3a98",x"ba1e",x"40b8",x"b74a",x"0000",x"3c00",x"8000",x"346a",x"3a98"),
(x"3aef",x"40b8",x"b74a",x"1018",x"2581",x"bbff",x"39d6",x"3942",x"ba1e",x"40b8",x"b74a",x"9418",x"257a",x"bbff",x"3bc1",x"3942",x"b941",x"4092",x"b751",x"0000",x"23e2",x"bbff",x"3ba1",x"392c"),
(x"3a12",x"34e4",x"b6b0",x"0000",x"0cea",x"bc00",x"3aed",x"37b1",x"3a12",x"3cb4",x"b6af",x"0000",x"0cea",x"bc00",x"3aed",x"3687",x"b941",x"3cb4",x"b6af",x"0000",x"0cea",x"bc00",x"39fa",x"3687"),
(x"3a11",x"4062",x"364d",x"0000",x"bc00",x"0000",x"3166",x"38eb",x"b940",x"4062",x"364d",x"0000",x"bc00",x"0000",x"3592",x"38eb",x"b940",x"4062",x"374f",x"0000",x"bc00",x"0000",x"3592",x"38dd"),
(x"3a11",x"40b6",x"364d",x"0000",x"8000",x"bc00",x"36e3",x"3866",x"b940",x"40b6",x"364d",x"0000",x"8000",x"bc00",x"3928",x"3867",x"b940",x"4062",x"364d",x"0a8d",x"068d",x"bc00",x"3928",x"383c"),
(x"3a11",x"0000",x"374f",x"bc00",x"0000",x"0000",x"3953",x"3861",x"3a11",x"0000",x"364d",x"bc00",x"0000",x"0000",x"3964",x"3861",x"3a11",x"4062",x"364d",x"bc00",x"0000",x"0000",x"3964",x"341e"),
(x"3a12",x"40b6",x"b694",x"0000",x"068d",x"3c00",x"2da6",x"38d9",x"3a12",x"3161",x"b694",x"0000",x"068d",x"3c00",x"3501",x"38d9",x"b941",x"3161",x"b694",x"0000",x"068d",x"3c00",x"3501",x"375f"),
(x"3a87",x"3154",x"364d",x"96f6",x"0000",x"bc00",x"36c0",x"3464",x"3a11",x"4062",x"364d",x"9018",x"8000",x"bc00",x"36e3",x"383c",x"3a11",x"0000",x"364d",x"9ac2",x"8000",x"bc00",x"36e3",x"340e"),
(x"3a87",x"3154",x"364d",x"96f6",x"0000",x"bc00",x"36c0",x"3464",x"3a88",x"40b6",x"364d",x"8e8d",x"068d",x"bc00",x"36bf",x"3866",x"3a11",x"4062",x"364d",x"9018",x"8000",x"bc00",x"36e3",x"383c"),
(x"3a87",x"3154",x"364d",x"bc00",x"0a8d",x"8e8d",x"315f",x"38e0",x"3a88",x"314b",x"b64f",x"bc00",x"8000",x"9418",x"2d91",x"38e0",x"3a88",x"40b6",x"b64d",x"bc00",x"0cea",x"8a8d",x"2d91",x"3aac"),
(x"3a88",x"40b6",x"b64d",x"0000",x"8a8d",x"3c00",x"3990",x"3887",x"3a88",x"314b",x"b64f",x"0000",x"868d",x"3c00",x"3990",x"3402",x"3a12",x"3161",x"b64f",x"0000",x"868d",x"3c00",x"397d",x"3404"),
(x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd",x"b940",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"38cd",x"3a11",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"374a"),
(x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd",x"b9b7",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"38d9",x"b940",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"38cd"),
(x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd",x"b9b7",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38d9",x"b9b7",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"38d9"),
(x"3a12",x"40b6",x"b694",x"0000",x"bc00",x"0000",x"1c61",x"374a",x"b941",x"40b6",x"b694",x"0000",x"bc00",x"0000",x"1c61",x"38cd",x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd"),
(x"3a88",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"3732",x"3a88",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"3732",x"3a12",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"374a"),
(x"3a12",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"374a",x"3a12",x"40b6",x"b694",x"0000",x"bc00",x"0000",x"1c61",x"374a",x"b941",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"38cd"),
(x"3a11",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"374a",x"3a88",x"40b6",x"364d",x"0000",x"bc00",x"0000",x"2d97",x"3732",x"3a12",x"40b6",x"b64d",x"0000",x"bc00",x"0000",x"1ef8",x"374a"),
(x"3a12",x"3161",x"b751",x"0000",x"bc00",x"0000",x"3bc8",x"347e",x"b941",x"3161",x"b751",x"0000",x"bc00",x"0000",x"39d2",x"347e",x"b941",x"3161",x"b694",x"0000",x"bc00",x"0000",x"39d2",x"3494"),
(x"3a12",x"40b6",x"b694",x"bc00",x"0000",x"0000",x"3879",x"3bef",x"3a12",x"40b6",x"b64d",x"bc00",x"0000",x"0000",x"3881",x"3bf0",x"3a12",x"3161",x"b64f",x"bc00",x"0000",x"0000",x"3895",x"3981"),
(x"3a12",x"8000",x"b751",x"bc00",x"8000",x"868d",x"387d",x"3912",x"3a12",x"3161",x"b751",x"bc00",x"0000",x"0000",x"3879",x"397f",x"3a12",x"3161",x"b694",x"bc00",x"0000",x"0000",x"388e",x"3980"),
(x"b941",x"3d3f",x"b751",x"0000",x"3c00",x"8000",x"39ce",x"345e",x"3a12",x"3d3f",x"b751",x"0000",x"3c00",x"8000",x"3bcd",x"345e",x"3a12",x"3d3f",x"b6b0",x"0000",x"3c00",x"8000",x"3bcd",x"3447"),
(x"3ad6",x"3d46",x"b544",x"3a14",x"38d9",x"337c",x"2dd6",x"20e8",x"3ae3",x"3d46",x"b578",x"39e8",x"3889",x"35d4",x"2dfc",x"2140",x"3ae3",x"3d41",x"b55a",x"39cc",x"38ee",x"34e9",x"2de7",x"218f"),
(x"3ad6",x"3d46",x"b544",x"3a14",x"38d9",x"337c",x"2dd6",x"20e8",x"3ae3",x"3d41",x"b55a",x"39cc",x"38ee",x"34e9",x"2de7",x"218f",x"3ae3",x"3d3b",x"b522",x"3a50",x"38e8",x"2604",x"2dbf",x"21f1"),
(x"3ad2",x"3d46",x"b515",x"3a7c",x"38ae",x"1c81",x"2db6",x"20d0",x"3ae3",x"3d3b",x"b522",x"3a50",x"38e8",x"2604",x"2dbf",x"21f1",x"3ae3",x"3d3a",x"b07b",x"3a7d",x"38ad",x"9e59",x"2b8b",x"21f1"),
(x"3ae3",x"3d3f",x"b00e",x"3a6d",x"3864",x"b364",x"2b40",x"219c",x"3ae3",x"3d46",x"af74",x"3a37",x"3832",x"b58f",x"2b03",x"211f",x"3ada",x"3d45",x"b010",x"3a60",x"3855",x"b446",x"2b42",x"20ee"),
(x"3ad4",x"3d45",x"b075",x"3aa1",x"3878",x"a594",x"2b88",x"20ca",x"3ae3",x"3d3a",x"b07b",x"3a7d",x"38ad",x"9e59",x"2b8b",x"21f1",x"3ae3",x"3d3f",x"b00e",x"3a6d",x"3864",x"b364",x"2b40",x"219c"),
(x"3aad",x"3d46",x"aca4",x"1d38",x"3c00",x"8cea",x"2392",x"2238",x"3aad",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"3ad2",x"3d46",x"b515",x"1f10",x"3c00",x"1018",x"2b3f",x"23cc"),
(x"3ae3",x"3d46",x"af74",x"9f79",x"3c00",x"9c81",x"25b4",x"243e",x"3aad",x"3d46",x"aca4",x"1d38",x"3c00",x"8cea",x"2392",x"2238",x"3ada",x"3d45",x"b010",x"a0d0",x"3bff",x"a081",x"262a",x"240d"),
(x"3aad",x"4070",x"aca4",x"8e8d",x"bc00",x"8000",x"2c87",x"257b",x"3ae3",x"4070",x"af8a",x"0000",x"bc00",x"0000",x"2d06",x"2458",x"3ada",x"4070",x"b010",x"0000",x"bc00",x"0000",x"2d20",x"248a"),
(x"3ad2",x"4070",x"b515",x"928d",x"bc00",x"868d",x"2f35",x"24b1",x"3aad",x"4070",x"b64e",x"91bc",x"bc00",x"8000",x"3005",x"257b",x"3aad",x"4070",x"aca4",x"8e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"3ac5",x"3d94",x"b504",x"3a04",x"8000",x"b945",x"31d8",x"3356",x"3ac5",x"4047",x"b504",x"3a04",x"8000",x"b945",x"31d7",x"35aa",x"3aad",x"404e",x"b53c",x"3a04",x"8000",x"b945",x"31be",x"35b4"),
(x"3ac5",x"3d94",x"b0a7",x"3a28",x"b91a",x"0000",x"30f8",x"290c",x"3ac5",x"3d94",x"b504",x"3a28",x"b91a",x"0000",x"31e3",x"290c",x"3aad",x"3d85",x"b53c",x"3a28",x"b91a",x"0000",x"31f6",x"2973"),
(x"3ac5",x"3d94",x"b0a7",x"3a1b",x"0000",x"392a",x"3165",x"3356",x"3aad",x"3d85",x"b032",x"3a1b",x"0000",x"392a",x"317f",x"3342",x"3aad",x"404e",x"b032",x"3a1b",x"0000",x"392a",x"317f",x"35b4"),
(x"3ae3",x"4073",x"b00e",x"3a59",x"b87c",x"b388",x"30f7",x"2c99",x"3ae3",x"4076",x"b07b",x"3a76",x"b8b6",x"9ffc",x"310a",x"2c8f",x"3ad4",x"4070",x"b075",x"3a96",x"b888",x"a5cf",x"3109",x"2cb3"),
(x"3ae3",x"4070",x"af8a",x"3a0f",x"b848",x"b5fa",x"30ea",x"2ca7",x"3ae3",x"4073",x"b00e",x"3a59",x"b87c",x"b388",x"30f7",x"2c99",x"3ada",x"4070",x"b010",x"3a44",x"b877",x"b45c",x"30f8",x"2cae"),
(x"3ac5",x"3d94",x"b0a7",x"3c00",x"0000",x"0000",x"301e",x"2c2f",x"3ac5",x"4047",x"b0a7",x"3c00",x"0000",x"0000",x"301e",x"3185",x"3ac5",x"4047",x"b504",x"3c00",x"0000",x"0000",x"2ea8",x"3185"),
(x"3aad",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"2b18",x"3aad",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"31dc",x"3aad",x"404e",x"b032",x"3c00",x"0000",x"0000",x"302e",x"318f"),
(x"3ae3",x"4076",x"b07b",x"3a76",x"b8b6",x"9ffc",x"310a",x"2c8f",x"3ae3",x"4076",x"b522",x"3a50",x"b8e8",x"25a8",x"3207",x"2c8f",x"3ad2",x"4070",x"b515",x"3a76",x"b8b6",x"1ac2",x"3203",x"2cb3"),
(x"3aad",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"2b18",x"3aad",x"3d85",x"b032",x"3c00",x"0000",x"0000",x"302e",x"2c1c",x"3aad",x"3d85",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"2c1c"),
(x"3aad",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"31dc",x"3aad",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2def",x"31dc",x"3aad",x"404e",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"318f"),
(x"3aad",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2def",x"2b18",x"3aad",x"3d85",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"2c1c",x"3aad",x"404e",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"318f"),
(x"3ae3",x"4076",x"b522",x"3a50",x"b8e8",x"25a8",x"3207",x"2c8f",x"3ae3",x"4073",x"b55a",x"39cc",x"b8ee",x"34e9",x"321b",x"2c9b",x"3ad6",x"4070",x"b544",x"3a14",x"b8d9",x"337c",x"3212",x"2cb0"),
(x"3ae3",x"4070",x"b578",x"39e8",x"b889",x"35d4",x"3226",x"2ca5",x"3ad6",x"4070",x"b544",x"3a14",x"b8d9",x"337c",x"3212",x"2cb0",x"3ae3",x"4073",x"b55a",x"39cc",x"b8ee",x"34e9",x"321b",x"2c9b"),
(x"3aad",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"2cf5",x"3aad",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"3350",x"3ae3",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"3350"),
(x"3ad6",x"3d46",x"b544",x"0000",x"3c00",x"8000",x"2b7e",x"23f3",x"3aad",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"3ae3",x"3d46",x"b578",x"0000",x"3c00",x"8000",x"2bc6",x"243e"),
(x"3ad7",x"3d83",x"aca4",x"0000",x"8000",x"bc00",x"312d",x"2d9a",x"3aad",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"3ae3",x"3d7a",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2d80"),
(x"3ac5",x"4047",x"b0a7",x"3a28",x"391a",x"0000",x"30f8",x"29e2",x"3aad",x"404e",x"b032",x"3a28",x"391a",x"0000",x"30e4",x"297b",x"3aad",x"404e",x"b53c",x"3a28",x"391a",x"0000",x"31f6",x"297b"),
(x"3ad6",x"4070",x"b544",x"90ea",x"bc00",x"868d",x"2f54",x"249e",x"3ae3",x"4070",x"b578",x"8e8d",x"bc00",x"868d",x"2f78",x"2458",x"3aad",x"4070",x"b64e",x"91bc",x"bc00",x"8000",x"3005",x"257b"),
(x"3ae3",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"2af0",x"3ae3",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"31e6",x"3ae3",x"3cb5",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"31f0"),
(x"3ae3",x"3d84",x"ac3b",x"39ce",x"340f",x"b91d",x"31ea",x"3351",x"3ad7",x"3d83",x"aca4",x"39a1",x"3488",x"b935",x"31de",x"3350",x"3ae3",x"3d7a",x"aca4",x"3950",x"3666",x"b90d",x"31e3",x"3342"),
(x"3aad",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"3aad",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"3ad0",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe"),
(x"3ae3",x"4057",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"330c",x"3aad",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"3ad3",x"404f",x"aca4",x"0000",x"8000",x"bc00",x"312a",x"32f6"),
(x"3ae3",x"3d84",x"ac3b",x"39ce",x"340f",x"b91d",x"31ea",x"3351",x"3ae3",x"3d92",x"abd9",x"3a32",x"17c8",x"b90f",x"31ef",x"3364",x"3ad0",x"3d91",x"aca4",x"3a39",x"1e0a",x"b906",x"31db",x"3363"),
(x"3ae3",x"3d92",x"abd9",x"3a32",x"17c8",x"b90f",x"31ef",x"3364",x"3ae3",x"404b",x"abe1",x"3a2a",x"975f",x"b918",x"31ef",x"35b8",x"3ad0",x"404b",x"aca4",x"3a32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"3ae3",x"404f",x"ac0f",x"39ea",x"b3b0",x"b908",x"31ed",x"35bd",x"3ad3",x"404f",x"aca4",x"39d3",x"b46b",x"b903",x"31dc",x"35bd",x"3ad0",x"404b",x"aca4",x"3a32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"3ae3",x"404f",x"ac0f",x"39ea",x"b3b0",x"b908",x"31ed",x"35bd",x"3ae3",x"4057",x"aca4",x"39ad",x"b59c",x"b8e3",x"31e3",x"35c9",x"3ad3",x"404f",x"aca4",x"39d3",x"b46b",x"b903",x"31dc",x"35bd"),
(x"3ae3",x"3d46",x"3587",x"3a16",x"3888",x"b50c",x"23b9",x"1d50",x"3ad8",x"3d45",x"3551",x"3a36",x"38b3",x"b345",x"2477",x"1cd0",x"3ae3",x"3d3e",x"3554",x"3a2c",x"38a8",x"b41a",x"246e",x"1e40"),
(x"3ae3",x"3d3a",x"3523",x"3a4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"3ae3",x"3d3e",x"3554",x"3a2c",x"38a8",x"b41a",x"246e",x"1e40",x"3ad8",x"3d45",x"3551",x"3a36",x"38b3",x"b345",x"2477",x"1cd0"),
(x"3ae3",x"3d3a",x"3099",x"3a5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"3ae3",x"3d3a",x"3523",x"3a4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"3ad2",x"3d45",x"351f",x"3a5d",x"38d8",x"9f93",x"2503",x"1c77"),
(x"3ae3",x"3d46",x"2f74",x"39ff",x"3898",x"3541",x"2af9",x"1d4d",x"3ae3",x"3d3e",x"3026",x"3a1b",x"38d7",x"3338",x"2aab",x"1e54",x"3ad7",x"3d45",x"302e",x"3a14",x"38b9",x"3455",x"2aa5",x"1cb4"),
(x"3ae3",x"3d3e",x"3026",x"3a1b",x"38d7",x"3338",x"2aab",x"1e54",x"3ae3",x"3d3a",x"3099",x"3a5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"3ad2",x"3d45",x"307d",x"3a66",x"38cb",x"2460",x"2a6e",x"1c77"),
(x"3ad2",x"3d45",x"351f",x"224c",x"3bff",x"0a8d",x"2705",x"2646",x"3aad",x"3d46",x"364e",x"1e0a",x"3c00",x"91bc",x"2392",x"257f",x"3aad",x"3d46",x"2ce6",x"2067",x"3c00",x"1018",x"2c69",x"257f"),
(x"3aad",x"3d46",x"2ce6",x"2067",x"3c00",x"1018",x"2c69",x"257f",x"3ae3",x"3d46",x"2f74",x"9ea7",x"3c00",x"1c67",x"2bf4",x"26a1",x"3ad7",x"3d45",x"302e",x"a025",x"3bff",x"2025",x"2ba5",x"265f"),
(x"3ae3",x"4070",x"2f82",x"0000",x"bc00",x"0000",x"2c02",x"26b0",x"3aad",x"4070",x"2ce6",x"8e8d",x"bc00",x"8000",x"2c74",x"27d3",x"3ada",x"4070",x"300c",x"0000",x"bc00",x"0000",x"2bd2",x"26e2"),
(x"3aad",x"4070",x"2ce6",x"8e8d",x"bc00",x"8000",x"2c74",x"27d3",x"3aad",x"4070",x"364e",x"91bc",x"bc00",x"8000",x"23e8",x"27d3",x"3ad2",x"4070",x"3524",x"928d",x"bc00",x"068d",x"2720",x"2709"),
(x"3ac5",x"3d94",x"3513",x"3a04",x"0000",x"3945",x"31a1",x"3356",x"3aad",x"3d85",x"354b",x"3a04",x"0000",x"3945",x"31ba",x"3342",x"3aad",x"404e",x"354b",x"3a04",x"0000",x"3945",x"31ba",x"35b4"),
(x"3ac5",x"3d94",x"30dd",x"3a28",x"b91a",x"0000",x"31e4",x"2aa8",x"3aad",x"3d85",x"3069",x"3a28",x"b91a",x"0000",x"31f8",x"2b0f",x"3aad",x"3d85",x"354b",x"3a28",x"b91a",x"0000",x"30ea",x"2b0f"),
(x"3aad",x"404e",x"3069",x"3a15",x"8000",x"b931",x"3183",x"35b4",x"3aad",x"3d85",x"3069",x"3a15",x"8000",x"b931",x"3183",x"3342",x"3ac5",x"3d94",x"30dd",x"3a15",x"8000",x"b931",x"319d",x"3356"),
(x"3ad4",x"4070",x"3071",x"3a97",x"b888",x"25b5",x"2a77",x"20ad",x"3ae3",x"4076",x"3076",x"3a77",x"b8b5",x"1f93",x"2a73",x"1f14",x"3ae3",x"4073",x"300a",x"3a59",x"b87c",x"3388",x"2abf",x"1fbf"),
(x"3ae3",x"4073",x"300a",x"3a59",x"b87c",x"3388",x"2abf",x"1fbf",x"3ae3",x"4070",x"2f82",x"3a0f",x"b848",x"35fa",x"2af4",x"2050",x"3ada",x"4070",x"300c",x"3a44",x"b877",x"345b",x"2abd",x"2088"),
(x"3ac5",x"4047",x"3513",x"3c00",x"0000",x"0000",x"2aa7",x"317f",x"3ac5",x"4047",x"30dd",x"3c00",x"0000",x"0000",x"272f",x"317f",x"3ac5",x"3d94",x"30dd",x"3c00",x"0000",x"0000",x"272f",x"2c38"),
(x"3aad",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"2b2a",x"3aad",x"3d85",x"3069",x"3c00",x"0000",x"0000",x"26a2",x"2c24",x"3aad",x"404e",x"3069",x"3c00",x"0000",x"0000",x"26a2",x"318a"),
(x"3ad2",x"4070",x"3524",x"3a76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"3ae3",x"4076",x"3532",x"3a50",x"b8e8",x"a587",x"24d1",x"1f14",x"3ae3",x"4076",x"3076",x"3a77",x"b8b5",x"1f93",x"2a73",x"1f14"),
(x"3aad",x"3d85",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"2c24",x"3aad",x"3d85",x"3069",x"3c00",x"0000",x"0000",x"26a2",x"2c24",x"3aad",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"2b2a"),
(x"3aad",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"31d6",x"3aad",x"404e",x"3069",x"3c00",x"0000",x"0000",x"26a2",x"318a",x"3aad",x"404e",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"318a"),
(x"3aad",x"404e",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"318a",x"3aad",x"3d85",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"2c24",x"3aad",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"2c00",x"2b2a"),
(x"3ad6",x"4070",x"3553",x"3a14",x"b8d9",x"b37c",x"2475",x"2093",x"3ae3",x"4073",x"3569",x"39cc",x"b8ee",x"b4e9",x"2433",x"1fda",x"3ae3",x"4076",x"3532",x"3a50",x"b8e8",x"a587",x"24d1",x"1f14"),
(x"3ad6",x"4070",x"3553",x"3a14",x"b8d9",x"b37c",x"2475",x"2093",x"3ae3",x"4070",x"3587",x"39e8",x"b889",x"b5d4",x"23b9",x"203c",x"3ae3",x"4073",x"3569",x"39cc",x"b8ee",x"b4e9",x"2433",x"1fda"),
(x"3aad",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"3138",x"2cf5",x"3ae3",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"315d",x"2cf5",x"3ae3",x"4070",x"364e",x"0000",x"8000",x"bc00",x"315d",x"3350"),
(x"3ad8",x"3d45",x"3551",x"94ea",x"3c00",x"9dd6",x"267b",x"2668",x"3ae3",x"3d46",x"3587",x"a04d",x"3c00",x"9cb5",x"25e8",x"26a2",x"3aad",x"3d46",x"364e",x"1e0a",x"3c00",x"91bc",x"2392",x"257f"),
(x"3ad9",x"3d84",x"2ce6",x"0000",x"0000",x"3c00",x"3169",x"2d69",x"3ae3",x"3d7a",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2d50",x"3aad",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"3aad",x"404e",x"354b",x"3a28",x"391a",x"0000",x"30ea",x"2b16",x"3aad",x"404e",x"3069",x"3a28",x"391a",x"0000",x"31f8",x"2b16",x"3ac5",x"4047",x"30dd",x"3a28",x"391a",x"0000",x"31e4",x"2b7e"),
(x"3ad6",x"4070",x"3553",x"90ea",x"bc00",x"068d",x"26a2",x"26f5",x"3aad",x"4070",x"364e",x"91bc",x"bc00",x"8000",x"23e8",x"27d3",x"3ae3",x"4070",x"3587",x"8e8d",x"bc00",x"0a8d",x"2613",x"26b0"),
(x"3ae3",x"4057",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3564",x"3ae3",x"404f",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"355a",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583"),
(x"3ad9",x"3d84",x"2ce6",x"39a5",x"3468",x"3938",x"3203",x"3350",x"3ae3",x"3d85",x"2c89",x"39d0",x"342d",x"3915",x"31f9",x"3351",x"3ae3",x"3d7a",x"2ce6",x"396d",x"35b1",x"3924",x"31ff",x"3342"),
(x"3ad0",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1",x"3ad1",x"3d90",x"2ce6",x"0000",x"0000",x"3c00",x"316e",x"2d8c",x"3aad",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"3aad",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"3ae3",x"4056",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"32f1",x"3ad4",x"404f",x"2ce6",x"0000",x"0000",x"3c00",x"316c",x"32dd"),
(x"3ae3",x"3d85",x"2c89",x"39d0",x"342d",x"3915",x"31f9",x"3351",x"3ad9",x"3d84",x"2ce6",x"39a5",x"3468",x"3938",x"3203",x"3350",x"3ad1",x"3d90",x"2ce6",x"3a4a",x"1ef6",x"38f1",x"3206",x"3362"),
(x"3ae3",x"3d92",x"2c35",x"3a20",x"184d",x"3924",x"31f3",x"3363",x"3ad1",x"3d90",x"2ce6",x"3a4a",x"1ef6",x"38f1",x"3206",x"3362",x"3ad0",x"404a",x"2ce6",x"3a20",x"935f",x"3925",x"3206",x"35b6"),
(x"3ae3",x"404b",x"2c40",x"39f4",x"9af6",x"3957",x"31f3",x"35b7",x"3ad0",x"404a",x"2ce6",x"3a20",x"935f",x"3925",x"3206",x"35b6",x"3ad4",x"404f",x"2ce6",x"39e5",x"b3cd",x"390b",x"3204",x"35bc"),
(x"3ae3",x"4056",x"2ce6",x"39b2",x"b5ad",x"38d8",x"31fe",x"35c7",x"3ae3",x"404e",x"2c57",x"39db",x"b485",x"38f4",x"31f4",x"35bc",x"3ad4",x"404f",x"2ce6",x"39e5",x"b3cd",x"390b",x"3204",x"35bc"),
(x"3ad6",x"3507",x"b544",x"3a14",x"38d9",x"337c",x"3214",x"2c6a",x"3ae3",x"3507",x"b578",x"39e8",x"3889",x"35d4",x"3227",x"2c75",x"3ae3",x"34f4",x"b55a",x"39cc",x"38ee",x"34e9",x"321c",x"2c7f"),
(x"3ad6",x"3507",x"b544",x"3a14",x"38d9",x"337c",x"3214",x"2c6a",x"3ae3",x"34f4",x"b55a",x"39cc",x"38ee",x"34e9",x"321c",x"2c7f",x"3ae3",x"34dc",x"b522",x"3a50",x"38e8",x"2604",x"3209",x"2c8b"),
(x"3ad2",x"3507",x"b515",x"3a7c",x"38ae",x"1c81",x"3204",x"2c67",x"3ae3",x"34dc",x"b522",x"3a50",x"38e8",x"2604",x"3209",x"2c8b",x"3ae3",x"34d8",x"b07b",x"3a7d",x"38ad",x"9e59",x"310c",x"2c8b"),
(x"3ae3",x"34eb",x"b00e",x"3a6d",x"3864",x"b364",x"30f9",x"2c80",x"3ae3",x"3507",x"af74",x"3a37",x"3832",x"b58f",x"30ea",x"2c71",x"3ada",x"3506",x"b010",x"3a5f",x"3855",x"b446",x"30f9",x"2c6a"),
(x"3ad4",x"3506",x"b075",x"3aa1",x"3878",x"a594",x"310b",x"2c66",x"3ae3",x"34d8",x"b07b",x"3a7d",x"38ad",x"9e59",x"310c",x"2c8b",x"3ae3",x"34eb",x"b00e",x"3a6d",x"3864",x"b364",x"30f9",x"2c80"),
(x"3aad",x"3507",x"aca4",x"1d38",x"3c00",x"8cea",x"2c87",x"224e",x"3aad",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"3ad2",x"3507",x"b515",x"1f10",x"3c00",x"1018",x"2f35",x"23e3"),
(x"3ae3",x"3507",x"af74",x"9f79",x"3c00",x"9c81",x"2d02",x"244a",x"3aad",x"3507",x"aca4",x"1d38",x"3c00",x"8cea",x"2c87",x"224e",x"3ada",x"3506",x"b010",x"a0d0",x"3bff",x"a081",x"2d20",x"2418"),
(x"3aad",x"3cac",x"aca4",x"8e8d",x"bc00",x"8000",x"2392",x"2570",x"3ae3",x"3cac",x"af8a",x"0000",x"bc00",x"0000",x"25c3",x"244d",x"3ada",x"3cac",x"b010",x"0000",x"bc00",x"0000",x"262a",x"247f"),
(x"3ad2",x"3cac",x"b515",x"928d",x"bc00",x"868d",x"2b3f",x"24a6",x"3aad",x"3cac",x"b64e",x"91bc",x"bc00",x"8000",x"2c74",x"2570",x"3aad",x"3cac",x"aca4",x"8e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"3ac5",x"3c5a",x"b504",x"3a04",x"8000",x"b945",x"3140",x"3598",x"3aad",x"3c69",x"b53c",x"3a04",x"8000",x"b945",x"3127",x"35a2",x"3aad",x"35ff",x"b53c",x"3a04",x"8000",x"b945",x"3127",x"335c"),
(x"3ac5",x"3638",x"b0a7",x"3a0b",x"b93d",x"0000",x"30fe",x"2bf4",x"3ac5",x"3638",x"b504",x"3a0b",x"b93d",x"0000",x"31e9",x"2bf4",x"3aad",x"35ff",x"b53c",x"3a0b",x"b93d",x"0000",x"31fc",x"2c2c"),
(x"3ac5",x"3c5a",x"b0a7",x"3a1b",x"0000",x"392a",x"30ec",x"3598",x"3ac5",x"3638",x"b0a7",x"3a1b",x"0000",x"392a",x"30ec",x"336f",x"3aad",x"35ff",x"b032",x"3a1b",x"0000",x"392a",x"3106",x"335c"),
(x"3ae3",x"3cb3",x"b00e",x"3a59",x"b87c",x"b388",x"2447",x"2120",x"3ae3",x"3cb8",x"b07b",x"3a76",x"b8b6",x"9fe2",x"24df",x"20ca",x"3ad4",x"3cac",x"b075",x"3a96",x"b888",x"a5d6",x"24d8",x"21ed"),
(x"3ae3",x"3cac",x"af8a",x"3a0f",x"b848",x"b5fa",x"23b9",x"2190",x"3ae3",x"3cb3",x"b00e",x"3a59",x"b87c",x"b388",x"2447",x"2120",x"3ada",x"3cac",x"b010",x"3a44",x"b877",x"b45c",x"244b",x"21c8"),
(x"3ac5",x"3638",x"b0a7",x"3c00",x"0000",x"0000",x"2ac8",x"330c",x"3ac5",x"3c5a",x"b0a7",x"3c00",x"0000",x"0000",x"2ac8",x"3545",x"3ac5",x"3c5a",x"b504",x"3c00",x"0000",x"0000",x"26b9",x"3545"),
(x"3aad",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"32d0",x"3aad",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"3575",x"3aad",x"3c69",x"b032",x"3c00",x"0000",x"0000",x"3036",x"354d"),
(x"3ae3",x"3cb8",x"b07b",x"3a76",x"b8b6",x"9fe2",x"24df",x"20ca",x"3ae3",x"3cb7",x"b522",x"3a50",x"b8e8",x"25a8",x"2a63",x"20cc",x"3ad2",x"3cac",x"b515",x"3a76",x"b8b6",x"1ac2",x"2a51",x"21ed"),
(x"3aad",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"32d0",x"3aad",x"35ff",x"b032",x"3c00",x"0000",x"0000",x"3036",x"331b",x"3aad",x"35ff",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"331b"),
(x"3aad",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"3575",x"3aad",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2ddb",x"3575",x"3aad",x"3c69",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"354d"),
(x"3aad",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2ddb",x"32d0",x"3aad",x"35ff",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"331b",x"3aad",x"3c69",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"354d"),
(x"3ae3",x"3cb7",x"b522",x"3a50",x"b8e8",x"25a8",x"2a63",x"20cc",x"3ae3",x"3cb1",x"b55a",x"39cc",x"b8ee",x"34e9",x"2ab1",x"212f",x"3ad6",x"3cac",x"b544",x"3a14",x"b8d9",x"337c",x"2a90",x"21d6"),
(x"3ae3",x"3cac",x"b578",x"39e8",x"b889",x"35d4",x"2add",x"217f",x"3ad6",x"3cac",x"b544",x"3a14",x"b8d9",x"337c",x"2a90",x"21d6",x"3ae3",x"3cb1",x"b55a",x"39cc",x"b8ee",x"34e9",x"2ab1",x"212f"),
(x"3aad",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"2d4a",x"3aad",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"333a",x"3ae3",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"333a"),
(x"3ad6",x"3507",x"b544",x"0000",x"3c00",x"8000",x"2f54",x"2404",x"3aad",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"3ae3",x"3507",x"b578",x"0000",x"3c00",x"8000",x"2f78",x"244a"),
(x"3ad7",x"35fb",x"aca4",x"0000",x"8000",x"bc00",x"31fc",x"2dee",x"3aad",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a",x"3ae3",x"35d5",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2dd4"),
(x"3ac5",x"3c5a",x"b0a7",x"3a28",x"391a",x"0000",x"30fe",x"2a76",x"3aad",x"3c69",x"b032",x"3a28",x"391a",x"0000",x"30ea",x"2a0f",x"3aad",x"3c69",x"b53c",x"3a28",x"391a",x"0000",x"31fc",x"2a0f"),
(x"3ad6",x"3cac",x"b544",x"90ea",x"bc00",x"868d",x"2b7e",x"2492",x"3ae3",x"3cac",x"b578",x"8e8d",x"bc00",x"8a8d",x"2bc6",x"244d",x"3aad",x"3cac",x"b64e",x"91bc",x"bc00",x"8000",x"2c74",x"2570"),
(x"3ae3",x"35fe",x"ac3b",x"39ce",x"340f",x"b91d",x"3219",x"3351",x"3ad7",x"35fb",x"aca4",x"39a1",x"3488",x"b935",x"320d",x"3350",x"3ae3",x"35d5",x"aca4",x"3950",x"3666",x"b90d",x"3212",x"3342"),
(x"3ad0",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"3aad",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"3aad",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"3ae3",x"3c7a",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"32f6",x"3aad",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"3ad3",x"3c6a",x"aca4",x"0000",x"8000",x"bc00",x"31f9",x"32e0"),
(x"3ae3",x"35fe",x"ac3b",x"39ce",x"340f",x"b91d",x"3219",x"3351",x"3ae3",x"3635",x"abd9",x"3a32",x"1818",x"b90f",x"321e",x"3364",x"3ad0",x"3631",x"aca4",x"3a39",x"1e59",x"b906",x"320a",x"3363"),
(x"3ae3",x"3635",x"abd9",x"3a32",x"1818",x"b90f",x"321e",x"3364",x"3ae3",x"3c61",x"abe1",x"3a2a",x"97c8",x"b918",x"321e",x"3597",x"3ad0",x"3c61",x"aca4",x"3a32",x"95bc",x"b90f",x"320a",x"3597"),
(x"3ae3",x"3c6a",x"ac0f",x"39ea",x"b3b0",x"b908",x"321c",x"359d",x"3ad3",x"3c6a",x"aca4",x"39d3",x"b46b",x"b903",x"320b",x"359d",x"3ad0",x"3c61",x"aca4",x"3a32",x"95bc",x"b90f",x"320a",x"3597"),
(x"3ae3",x"3c6a",x"ac0f",x"39ea",x"b3b0",x"b908",x"321c",x"359d",x"3ae3",x"3c7a",x"aca4",x"39ad",x"b59c",x"b8e3",x"3212",x"35a9",x"3ad3",x"3c6a",x"aca4",x"39d3",x"b46b",x"b903",x"320b",x"359d"),
(x"3ae3",x"3507",x"3587",x"3a16",x"3888",x"b50c",x"2b07",x"1d50",x"3ad8",x"3505",x"3551",x"3a36",x"38b3",x"b345",x"2b55",x"1cd0",x"3ae3",x"34ea",x"3554",x"3a2c",x"38a8",x"b41a",x"2b50",x"1e40"),
(x"3ae3",x"34db",x"3523",x"3a4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"3ae3",x"34ea",x"3554",x"3a2c",x"38a8",x"b41a",x"2b50",x"1e40",x"3ad8",x"3505",x"3551",x"3a36",x"38b3",x"b345",x"2b55",x"1cd0"),
(x"3ae3",x"34d8",x"3099",x"3a5b",x"38da",x"1d38",x"2dba",x"1ed9",x"3ae3",x"34db",x"3523",x"3a4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"3ad2",x"3506",x"351f",x"3a5d",x"38d8",x"9f93",x"2b9a",x"1c77"),
(x"3ae3",x"3507",x"2f74",x"39ff",x"3898",x"3541",x"2e09",x"1d4d",x"3ae3",x"34e8",x"3026",x"3a1b",x"38d7",x"3338",x"2de2",x"1e54",x"3ad7",x"3506",x"302e",x"3a14",x"38b9",x"3455",x"2ddf",x"1cb4"),
(x"3ae3",x"34e8",x"3026",x"3a1b",x"38d7",x"3338",x"2de2",x"1e54",x"3ae3",x"34d8",x"3099",x"3a5b",x"38da",x"1d38",x"2dba",x"1ed9",x"3ad2",x"3506",x"307d",x"3a66",x"38cb",x"2460",x"2dc4",x"1c77"),
(x"3ad2",x"3506",x"351f",x"2259",x"3bff",x"068d",x"2d56",x"2651",x"3aad",x"3507",x"364e",x"1e0a",x"3c00",x"91bc",x"2c87",x"258a",x"3aad",x"3507",x"2ce6",x"2067",x"3c00",x"1018",x"2fff",x"258a"),
(x"3aad",x"3507",x"2ce6",x"2067",x"3c00",x"1018",x"2fff",x"258a",x"3ae3",x"3507",x"2f74",x"9ea7",x"3c00",x"1c67",x"2f8f",x"26ad",x"3ad7",x"3506",x"302e",x"a032",x"3bff",x"2025",x"2f68",x"266a"),
(x"3ae3",x"3cac",x"2f82",x"0000",x"bc00",x"0000",x"2f8d",x"26bb",x"3aad",x"3cac",x"2ce6",x"8e8d",x"bc00",x"8000",x"2fff",x"27de",x"3ada",x"3cac",x"300c",x"0000",x"bc00",x"0000",x"2f73",x"26ed"),
(x"3aad",x"3cac",x"2ce6",x"8e8d",x"bc00",x"8000",x"2fff",x"27de",x"3aad",x"3cac",x"364e",x"91bc",x"bc00",x"8000",x"2c87",x"27de",x"3ad2",x"3cac",x"3524",x"928d",x"bc00",x"068d",x"2d52",x"2714"),
(x"3aad",x"3600",x"354b",x"3a04",x"0000",x"3945",x"315d",x"335c",x"3aad",x"3c69",x"354b",x"3a04",x"0000",x"3945",x"315d",x"35a1",x"3ac5",x"3c5a",x"3513",x"3a04",x"0000",x"3945",x"3144",x"3597"),
(x"3ac5",x"3639",x"30dd",x"3a0f",x"b938",x"0000",x"31e4",x"2c30",x"3aad",x"3600",x"3069",x"3a0f",x"b938",x"0000",x"31f8",x"2c62",x"3aad",x"3600",x"354b",x"3a0f",x"b938",x"0000",x"30ea",x"2c62"),
(x"3ac5",x"3c5a",x"30dd",x"3a15",x"8000",x"b931",x"3123",x"3597",x"3aad",x"3c69",x"3069",x"3a15",x"8000",x"b931",x"3109",x"35a1",x"3aad",x"3600",x"3069",x"3a15",x"8000",x"b931",x"3109",x"335c"),
(x"3ad4",x"3cac",x"3071",x"3a96",x"b888",x"25b5",x"2dc8",x"20ad",x"3ae3",x"3cb8",x"3076",x"3a77",x"b8b5",x"1f93",x"2dc6",x"1f14",x"3ae3",x"3cb3",x"300a",x"3a59",x"b87c",x"3388",x"2dec",x"1fbf"),
(x"3ae3",x"3cb3",x"300a",x"3a59",x"b87c",x"3388",x"2dec",x"1fbf",x"3ae3",x"3cac",x"2f82",x"3a0f",x"b848",x"35fa",x"2e07",x"2050",x"3ada",x"3cac",x"300c",x"3a44",x"b877",x"345c",x"2deb",x"2088"),
(x"3ac5",x"3c5a",x"3513",x"3c00",x"0000",x"0000",x"3028",x"3547",x"3ac5",x"3c5a",x"30dd",x"3c00",x"0000",x"0000",x"2eaa",x"3547",x"3ac5",x"3639",x"30dd",x"3c00",x"0000",x"0000",x"2eaa",x"3323"),
(x"3aad",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"32b8",x"3aad",x"3600",x"3069",x"3c00",x"0000",x"0000",x"2658",x"3304",x"3aad",x"3c69",x"3069",x"3c00",x"0000",x"0000",x"2658",x"354a"),
(x"3ad2",x"3cac",x"3524",x"3a76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"3ae3",x"3cb7",x"3532",x"3a50",x"b8e8",x"a587",x"2b82",x"1f14",x"3ae3",x"3cb8",x"3076",x"3a77",x"b8b5",x"1f93",x"2dc6",x"1f14"),
(x"3aad",x"3600",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"3304",x"3aad",x"3600",x"3069",x"3c00",x"0000",x"0000",x"2658",x"3304",x"3aad",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"32b8"),
(x"3aad",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"3573",x"3aad",x"3c69",x"3069",x"3c00",x"0000",x"0000",x"2658",x"354a",x"3aad",x"3c69",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"354a"),
(x"3aad",x"3c69",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"354a",x"3aad",x"3600",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"3304",x"3aad",x"3507",x"364e",x"3c00",x"0000",x"0000",x"2c23",x"32b8"),
(x"3ad6",x"3cac",x"3553",x"3a14",x"b8d9",x"b37c",x"2b54",x"2093",x"3ae3",x"3cb1",x"3569",x"39cc",x"b8ee",x"b4e9",x"2b33",x"1fda",x"3ae3",x"3cb7",x"3532",x"3a50",x"b8e8",x"a587",x"2b82",x"1f14"),
(x"3ad6",x"3cac",x"3553",x"3a14",x"b8d9",x"b37c",x"2b54",x"2093",x"3ae3",x"3cac",x"3587",x"39e8",x"b889",x"b5d4",x"2b07",x"203c",x"3ae3",x"3cb1",x"3569",x"39cc",x"b8ee",x"b4e9",x"2b33",x"1fda"),
(x"3aad",x"3507",x"364e",x"0000",x"8000",x"bc00",x"318d",x"2d4a",x"3ae3",x"3507",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"2d4a",x"3ae3",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"333a"),
(x"3ad8",x"3505",x"3551",x"94ea",x"3c00",x"9dd6",x"2d34",x"2673",x"3ae3",x"3507",x"3587",x"a04d",x"3c00",x"9cb5",x"2d0f",x"26ad",x"3aad",x"3507",x"364e",x"1e0a",x"3c00",x"91bc",x"2c87",x"258a"),
(x"3ad9",x"35fd",x"2ce6",x"0000",x"0000",x"3c00",x"31bd",x"2def",x"3ae3",x"35d7",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2dd5",x"3aad",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"3aad",x"3c69",x"354b",x"3a28",x"391a",x"0000",x"30ea",x"2b85",x"3aad",x"3c69",x"3069",x"3a28",x"391a",x"0000",x"31f8",x"2b85",x"3ac5",x"3c5a",x"30dd",x"3a28",x"391a",x"0000",x"31e4",x"2bed"),
(x"3ad6",x"3cac",x"3553",x"8a8d",x"bc00",x"0cea",x"2d33",x"2701",x"3aad",x"3cac",x"364e",x"91bc",x"bc00",x"8000",x"2c87",x"27de",x"3ae3",x"3cac",x"3587",x"8e8d",x"bc00",x"0a8d",x"2d0f",x"26bb"),
(x"3ae3",x"3c7a",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31a9",x"3ae3",x"3c6a",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"3195",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6"),
(x"3ad9",x"35fd",x"2ce6",x"39a5",x"3468",x"3938",x"3231",x"3350",x"3ae3",x"3601",x"2c89",x"39d0",x"342d",x"3915",x"3227",x"3351",x"3ae3",x"35d7",x"2ce6",x"396d",x"35b1",x"3924",x"322d",x"3342"),
(x"3ad0",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4",x"3ad1",x"3630",x"2ce6",x"0000",x"0000",x"3c00",x"31c2",x"2e11",x"3aad",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"3aad",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"3ae3",x"3c78",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"32f4",x"3ad4",x"3c69",x"2ce6",x"0000",x"0000",x"3c00",x"31c0",x"32e0"),
(x"3ae3",x"3601",x"2c89",x"39d0",x"342d",x"3915",x"3227",x"3351",x"3ad9",x"35fd",x"2ce6",x"39a5",x"3468",x"3938",x"3231",x"3350",x"3ad1",x"3630",x"2ce6",x"3a4a",x"1f5f",x"38f1",x"3235",x"3362"),
(x"3ae3",x"3635",x"2c35",x"3a20",x"1881",x"3924",x"3221",x"3363",x"3ad1",x"3630",x"2ce6",x"3a4a",x"1f5f",x"38f1",x"3235",x"3362",x"3ad0",x"3c60",x"2ce6",x"3a20",x"9418",x"3925",x"3234",x"3596"),
(x"3ae3",x"3c61",x"2c40",x"39f4",x"9b5f",x"3957",x"3221",x"3597",x"3ad0",x"3c60",x"2ce6",x"3a20",x"9418",x"3925",x"3234",x"3596",x"3ad4",x"3c69",x"2ce6",x"39e5",x"b3cc",x"390b",x"3233",x"359c"),
(x"3ae3",x"3c78",x"2ce6",x"39b2",x"b5ad",x"38d8",x"322c",x"35a7",x"3ae3",x"3c69",x"2c57",x"39db",x"b485",x"38f4",x"3223",x"359c",x"3ad4",x"3c69",x"2ce6",x"39e5",x"b3cc",x"390b",x"3233",x"359c"),
(x"3ae3",x"34db",x"3523",x"3c00",x"0000",x"0000",x"3029",x"2abb",x"3ae3",x"34d8",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"2ab8",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"0000",x"3753",x"3c00",x"0000",x"0000",x"30de",x"1e82",x"3ae3",x"3227",x"3753",x"3c00",x"0000",x"0000",x"30de",x"2890",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"31e6",x"3ae3",x"3cb1",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"31ec",x"3ae3",x"3d41",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"329b"),
(x"3ae3",x"8000",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"1e82",x"3ae3",x"8000",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"1e82",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c"),
(x"3ae3",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"2af0",x"3ae3",x"3154",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"280f",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c"),
(x"3ae3",x"4056",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3563",x"3ae3",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3583",x"3ae3",x"404e",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"355a"),
(x"3ae3",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"3583",x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7",x"3ae3",x"3d42",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"329d"),
(x"3ae3",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"32a1",x"3ae3",x"3d42",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"329d",x"3ae3",x"3cb5",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"31f0"),
(x"3ad2",x"3d46",x"b515",x"3a7c",x"38ae",x"1c81",x"2db6",x"20d0",x"3ad6",x"3d46",x"b544",x"3a14",x"38d9",x"337c",x"2dd6",x"20e8",x"3ae3",x"3d3b",x"b522",x"3a50",x"38e8",x"2604",x"2dbf",x"21f1"),
(x"3ad4",x"3d45",x"b075",x"3aa1",x"3878",x"a594",x"2b88",x"20ca",x"3ad2",x"3d46",x"b515",x"3a7c",x"38ae",x"1c81",x"2db6",x"20d0",x"3ae3",x"3d3a",x"b07b",x"3a7d",x"38ad",x"9e59",x"2b8b",x"21f1"),
(x"3ada",x"3d45",x"b010",x"3a60",x"3855",x"b446",x"2b42",x"20ee",x"3ad4",x"3d45",x"b075",x"3aa1",x"3878",x"a594",x"2b88",x"20ca",x"3ae3",x"3d3f",x"b00e",x"3a6d",x"3864",x"b364",x"2b40",x"219c"),
(x"3ad4",x"3d45",x"b075",x"24a2",x"3bff",x"1481",x"26b4",x"23d9",x"3aad",x"3d46",x"aca4",x"1d38",x"3c00",x"8cea",x"2392",x"2238",x"3ad2",x"3d46",x"b515",x"1f10",x"3c00",x"1018",x"2b3f",x"23cc"),
(x"3aad",x"3d46",x"aca4",x"1d38",x"3c00",x"8cea",x"2392",x"2238",x"3ae3",x"3d46",x"af74",x"9f79",x"3c00",x"9c81",x"25b4",x"243e",x"3ae3",x"3d46",x"aca4",x"0000",x"3c00",x"8000",x"2392",x"243e"),
(x"3ad4",x"3d45",x"b075",x"24a2",x"3bff",x"1481",x"26b4",x"23d9",x"3ada",x"3d45",x"b010",x"a0d0",x"3bff",x"a081",x"262a",x"240d",x"3aad",x"3d46",x"aca4",x"1d38",x"3c00",x"8cea",x"2392",x"2238"),
(x"3aad",x"4070",x"aca4",x"8e8d",x"bc00",x"8000",x"2c87",x"257b",x"3ada",x"4070",x"b010",x"0000",x"bc00",x"0000",x"2d20",x"248a",x"3ad4",x"4070",x"b075",x"0000",x"bc00",x"0000",x"2d42",x"24ab"),
(x"3ae3",x"4070",x"aca4",x"0000",x"bc00",x"0000",x"2c87",x"2458",x"3ae3",x"4070",x"af8a",x"0000",x"bc00",x"0000",x"2d06",x"2458",x"3aad",x"4070",x"aca4",x"8e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"3ad4",x"4070",x"b075",x"0000",x"bc00",x"0000",x"2d42",x"24ab",x"3ad2",x"4070",x"b515",x"928d",x"bc00",x"868d",x"2f35",x"24b1",x"3aad",x"4070",x"aca4",x"8e8d",x"bc00",x"8000",x"2c87",x"257b"),
(x"3aad",x"3d85",x"b53c",x"3a04",x"8000",x"b945",x"31be",x"3342",x"3ac5",x"3d94",x"b504",x"3a04",x"8000",x"b945",x"31d8",x"3356",x"3aad",x"404e",x"b53c",x"3a04",x"8000",x"b945",x"31be",x"35b4"),
(x"3aad",x"3d85",x"b032",x"3a28",x"b91a",x"0000",x"30e4",x"2973",x"3ac5",x"3d94",x"b0a7",x"3a28",x"b91a",x"0000",x"30f8",x"290c",x"3aad",x"3d85",x"b53c",x"3a28",x"b91a",x"0000",x"31f6",x"2973"),
(x"3ac5",x"4047",x"b0a7",x"3a1b",x"0000",x"392a",x"3165",x"35aa",x"3ac5",x"3d94",x"b0a7",x"3a1b",x"0000",x"392a",x"3165",x"3356",x"3aad",x"404e",x"b032",x"3a1b",x"0000",x"392a",x"317f",x"35b4"),
(x"3ada",x"4070",x"b010",x"3a44",x"b877",x"b45c",x"30f8",x"2cae",x"3ae3",x"4073",x"b00e",x"3a59",x"b87c",x"b388",x"30f7",x"2c99",x"3ad4",x"4070",x"b075",x"3a96",x"b888",x"a5cf",x"3109",x"2cb3"),
(x"3ac5",x"3d94",x"b504",x"3c00",x"0000",x"0000",x"2ea9",x"2c2f",x"3ac5",x"3d94",x"b0a7",x"3c00",x"0000",x"0000",x"301e",x"2c2f",x"3ac5",x"4047",x"b504",x"3c00",x"0000",x"0000",x"2ea8",x"3185"),
(x"3aad",x"3d85",x"b032",x"3c00",x"0000",x"0000",x"302e",x"2c1c",x"3aad",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"2b18",x"3aad",x"404e",x"b032",x"3c00",x"0000",x"0000",x"302e",x"318f"),
(x"3ad4",x"4070",x"b075",x"3a96",x"b888",x"a5cf",x"3109",x"2cb3",x"3ae3",x"4076",x"b07b",x"3a76",x"b8b6",x"9ffc",x"310a",x"2c8f",x"3ad2",x"4070",x"b515",x"3a76",x"b8b6",x"1ac2",x"3203",x"2cb3"),
(x"3aad",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2def",x"2b18",x"3aad",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"2b18",x"3aad",x"3d85",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"2c1c"),
(x"3aad",x"404e",x"b032",x"3c00",x"0000",x"0000",x"302e",x"318f",x"3aad",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"3073",x"31dc",x"3aad",x"404e",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"318f"),
(x"3aad",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2def",x"31dc",x"3aad",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2def",x"2b18",x"3aad",x"404e",x"b53c",x"3c00",x"0000",x"0000",x"2e8c",x"318f"),
(x"3ad2",x"4070",x"b515",x"3a76",x"b8b6",x"1ac2",x"3203",x"2cb3",x"3ae3",x"4076",x"b522",x"3a50",x"b8e8",x"25a8",x"3207",x"2c8f",x"3ad6",x"4070",x"b544",x"3a14",x"b8d9",x"337c",x"3212",x"2cb0"),
(x"3ae3",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"2cf5",x"3aad",x"3d46",x"b64e",x"0000",x"0000",x"3c00",x"310c",x"2cf5",x"3ae3",x"4070",x"b64e",x"0000",x"0000",x"3c00",x"30e7",x"3350"),
(x"3ae3",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"243e",x"3ae3",x"3d46",x"b578",x"0000",x"3c00",x"8000",x"2bc6",x"243e",x"3aad",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238"),
(x"3ad2",x"3d46",x"b515",x"1f10",x"3c00",x"1018",x"2b3f",x"23cc",x"3aad",x"3d46",x"b64e",x"0000",x"3c00",x"8000",x"2c74",x"2238",x"3ad6",x"3d46",x"b544",x"0000",x"3c00",x"8000",x"2b7e",x"23f3"),
(x"3ae3",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2cf5",x"3ae3",x"3d7a",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"2d80",x"3aad",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5"),
(x"3ad0",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe",x"3aad",x"3d46",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"2cf5",x"3ad7",x"3d83",x"aca4",x"0000",x"8000",x"bc00",x"312d",x"2d9a"),
(x"3ac5",x"4047",x"b504",x"3a28",x"391a",x"0000",x"31e3",x"29e2",x"3ac5",x"4047",x"b0a7",x"3a28",x"391a",x"0000",x"30f8",x"29e2",x"3aad",x"404e",x"b53c",x"3a28",x"391a",x"0000",x"31f6",x"297b"),
(x"3ae3",x"4070",x"b64e",x"91bc",x"bc00",x"8000",x"3005",x"2458",x"3aad",x"4070",x"b64e",x"91bc",x"bc00",x"8000",x"3005",x"257b",x"3ae3",x"4070",x"b578",x"8e8d",x"bc00",x"868d",x"2f78",x"2458"),
(x"3ad2",x"4070",x"b515",x"928d",x"bc00",x"868d",x"2f35",x"24b1",x"3ad6",x"4070",x"b544",x"90ea",x"bc00",x"868d",x"2f54",x"249e",x"3aad",x"4070",x"b64e",x"91bc",x"bc00",x"8000",x"3005",x"257b"),
(x"3ae3",x"3154",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"280f",x"3ae3",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"2af0",x"3ae3",x"3cb5",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"31f0"),
(x"3ad0",x"404b",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"32eb",x"3aad",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"3ad0",x"3d91",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"2dbe"),
(x"3aad",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350",x"3ae3",x"4057",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"330c",x"3ae3",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3135",x"3350"),
(x"3ad0",x"404b",x"aca4",x"0000",x"8000",x"bc00",x"3128",x"32eb",x"3ad3",x"404f",x"aca4",x"0000",x"8000",x"bc00",x"312a",x"32f6",x"3aad",x"4070",x"aca4",x"0000",x"8000",x"bc00",x"3110",x"3350"),
(x"3ad7",x"3d83",x"aca4",x"39a1",x"3488",x"b935",x"31de",x"3350",x"3ae3",x"3d84",x"ac3b",x"39ce",x"340f",x"b91d",x"31ea",x"3351",x"3ad0",x"3d91",x"aca4",x"3a39",x"1e0a",x"b906",x"31db",x"3363"),
(x"3ad0",x"3d91",x"aca4",x"3a39",x"1e0a",x"b906",x"31db",x"3363",x"3ae3",x"3d92",x"abd9",x"3a32",x"17c8",x"b90f",x"31ef",x"3364",x"3ad0",x"404b",x"aca4",x"3a32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"3ae3",x"404b",x"abe1",x"3a2a",x"975f",x"b918",x"31ef",x"35b8",x"3ae3",x"404f",x"ac0f",x"39ea",x"b3b0",x"b908",x"31ed",x"35bd",x"3ad0",x"404b",x"aca4",x"3a32",x"95bc",x"b90f",x"31db",x"35b8"),
(x"3ad2",x"3d45",x"351f",x"3a5d",x"38d8",x"9f93",x"2503",x"1c77",x"3ae3",x"3d3a",x"3523",x"3a4f",x"38ea",x"a57a",x"24f8",x"1ec7",x"3ad8",x"3d45",x"3551",x"3a36",x"38b3",x"b345",x"2477",x"1cd0"),
(x"3ad2",x"3d45",x"307d",x"3a66",x"38cb",x"2460",x"2a6e",x"1c77",x"3ae3",x"3d3a",x"3099",x"3a5b",x"38da",x"1d38",x"2a5b",x"1ed9",x"3ad2",x"3d45",x"351f",x"3a5d",x"38d8",x"9f93",x"2503",x"1c77"),
(x"3ad7",x"3d45",x"302e",x"3a14",x"38b9",x"3455",x"2aa5",x"1cb4",x"3ae3",x"3d3e",x"3026",x"3a1b",x"38d7",x"3338",x"2aab",x"1e54",x"3ad2",x"3d45",x"307d",x"3a66",x"38cb",x"2460",x"2a6e",x"1c77"),
(x"3ad2",x"3d45",x"307d",x"2404",x"3bff",x"8e8d",x"2b6f",x"2646",x"3ad2",x"3d45",x"351f",x"224c",x"3bff",x"0a8d",x"2705",x"2646",x"3aad",x"3d46",x"2ce6",x"2067",x"3c00",x"1018",x"2c69",x"257f"),
(x"3aad",x"3d46",x"2ce6",x"2067",x"3c00",x"1018",x"2c69",x"257f",x"3ad7",x"3d45",x"302e",x"a025",x"3bff",x"2025",x"2ba5",x"265f",x"3ad2",x"3d45",x"307d",x"2404",x"3bff",x"8e8d",x"2b6f",x"2646"),
(x"3ae3",x"3d46",x"2ce6",x"0000",x"3c00",x"8000",x"2c69",x"26a1",x"3ae3",x"3d46",x"2f74",x"9ea7",x"3c00",x"1c67",x"2bf4",x"26a1",x"3aad",x"3d46",x"2ce6",x"2067",x"3c00",x"1018",x"2c69",x"257f"),
(x"3aad",x"4070",x"2ce6",x"8e8d",x"bc00",x"8000",x"2c74",x"27d3",x"3ae3",x"4070",x"2f82",x"0000",x"bc00",x"0000",x"2c02",x"26b0",x"3ae3",x"4070",x"2ce6",x"0000",x"bc00",x"0000",x"2c74",x"26b0"),
(x"3ad4",x"4070",x"3071",x"0000",x"bc00",x"0000",x"2b8d",x"2702",x"3ada",x"4070",x"300c",x"0000",x"bc00",x"0000",x"2bd2",x"26e2",x"3aad",x"4070",x"2ce6",x"8e8d",x"bc00",x"8000",x"2c74",x"27d3"),
(x"3ad4",x"4070",x"3071",x"0000",x"bc00",x"0000",x"2b8d",x"2702",x"3aad",x"4070",x"2ce6",x"8e8d",x"bc00",x"8000",x"2c74",x"27d3",x"3ad2",x"4070",x"3524",x"928d",x"bc00",x"068d",x"2720",x"2709"),
(x"3ac5",x"4047",x"3513",x"3a04",x"0000",x"3945",x"31a0",x"35aa",x"3ac5",x"3d94",x"3513",x"3a04",x"0000",x"3945",x"31a1",x"3356",x"3aad",x"404e",x"354b",x"3a04",x"0000",x"3945",x"31ba",x"35b4"),
(x"3ac5",x"3d94",x"3513",x"3a28",x"b91a",x"0000",x"30fd",x"2aa8",x"3ac5",x"3d94",x"30dd",x"3a28",x"b91a",x"0000",x"31e4",x"2aa8",x"3aad",x"3d85",x"354b",x"3a28",x"b91a",x"0000",x"30ea",x"2b0f"),
(x"3ac5",x"4047",x"30dd",x"3a15",x"8000",x"b931",x"319d",x"35aa",x"3aad",x"404e",x"3069",x"3a15",x"8000",x"b931",x"3183",x"35b4",x"3ac5",x"3d94",x"30dd",x"3a15",x"8000",x"b931",x"319d",x"3356"),
(x"3ada",x"4070",x"300c",x"3a44",x"b877",x"345b",x"2abd",x"2088",x"3ad4",x"4070",x"3071",x"3a97",x"b888",x"25b5",x"2a77",x"20ad",x"3ae3",x"4073",x"300a",x"3a59",x"b87c",x"3388",x"2abf",x"1fbf"),
(x"3ac5",x"3d94",x"3513",x"3c00",x"0000",x"0000",x"2aa7",x"2c38",x"3ac5",x"4047",x"3513",x"3c00",x"0000",x"0000",x"2aa7",x"317f",x"3ac5",x"3d94",x"30dd",x"3c00",x"0000",x"0000",x"272f",x"2c38"),
(x"3aad",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"31d6",x"3aad",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"2b2a",x"3aad",x"404e",x"3069",x"3c00",x"0000",x"0000",x"26a2",x"318a"),
(x"3ad4",x"4070",x"3071",x"3a97",x"b888",x"25b5",x"2a77",x"20ad",x"3ad2",x"4070",x"3524",x"3a76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"3ae3",x"4076",x"3076",x"3a77",x"b8b5",x"1f93",x"2a73",x"1f14"),
(x"3aad",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"2c00",x"2b2a",x"3aad",x"3d85",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"2c24",x"3aad",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"2b2a"),
(x"3aad",x"4070",x"364e",x"3c00",x"0000",x"0000",x"2c00",x"31d6",x"3aad",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2465",x"31d6",x"3aad",x"404e",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"318a"),
(x"3aad",x"4070",x"364e",x"3c00",x"0000",x"0000",x"2c00",x"31d6",x"3aad",x"404e",x"354b",x"3c00",x"0000",x"0000",x"2ad8",x"318a",x"3aad",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"2c00",x"2b2a"),
(x"3ad2",x"4070",x"3524",x"3a76",x"b8b6",x"9a8d",x"24f4",x"20ab",x"3ad6",x"4070",x"3553",x"3a14",x"b8d9",x"b37c",x"2475",x"2093",x"3ae3",x"4076",x"3532",x"3a50",x"b8e8",x"a587",x"24d1",x"1f14"),
(x"3aad",x"4070",x"364e",x"0000",x"8000",x"bc00",x"3138",x"3350",x"3aad",x"3d46",x"364e",x"0000",x"8000",x"bc00",x"3138",x"2cf5",x"3ae3",x"4070",x"364e",x"0000",x"8000",x"bc00",x"315d",x"3350"),
(x"3ae3",x"3d46",x"364e",x"0000",x"3c00",x"8000",x"2392",x"26a2",x"3aad",x"3d46",x"364e",x"1e0a",x"3c00",x"91bc",x"2392",x"257f",x"3ae3",x"3d46",x"3587",x"a04d",x"3c00",x"9cb5",x"25e8",x"26a2"),
(x"3ad2",x"3d45",x"351f",x"224c",x"3bff",x"0a8d",x"2705",x"2646",x"3ad8",x"3d45",x"3551",x"94ea",x"3c00",x"9dd6",x"267b",x"2668",x"3aad",x"3d46",x"364e",x"1e0a",x"3c00",x"91bc",x"2392",x"257f"),
(x"3ae3",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2cc3",x"3aad",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3",x"3ae3",x"3d7a",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"2d50"),
(x"3ad1",x"3d90",x"2ce6",x"0000",x"0000",x"3c00",x"316e",x"2d8c",x"3ad9",x"3d84",x"2ce6",x"0000",x"0000",x"3c00",x"3169",x"2d69",x"3aad",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"3ac5",x"4047",x"3513",x"3a28",x"391a",x"0000",x"30fd",x"2b7e",x"3aad",x"404e",x"354b",x"3a28",x"391a",x"0000",x"30ea",x"2b16",x"3ac5",x"4047",x"30dd",x"3a28",x"391a",x"0000",x"31e4",x"2b7e"),
(x"3ae3",x"4070",x"364e",x"91bc",x"bc00",x"8000",x"23e8",x"26b0",x"3ae3",x"4070",x"3587",x"8e8d",x"bc00",x"0a8d",x"2613",x"26b0",x"3aad",x"4070",x"364e",x"91bc",x"bc00",x"8000",x"23e8",x"27d3"),
(x"3ad2",x"4070",x"3524",x"928d",x"bc00",x"068d",x"2720",x"2709",x"3aad",x"4070",x"364e",x"91bc",x"bc00",x"8000",x"23e8",x"27d3",x"3ad6",x"4070",x"3553",x"90ea",x"bc00",x"068d",x"26a2",x"26f5"),
(x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1",x"3ae3",x"3d84",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"32ed",x"3ae3",x"3d7a",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32e0"),
(x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1",x"3ae3",x"3d84",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"32ed",x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"3ae3",x"3d7a",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32e1",x"3ae3",x"3d85",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"32ee",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1"),
(x"3ae3",x"404b",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"3555",x"3ae3",x"3d92",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"32fe",x"3ae3",x"3d92",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"32fe"),
(x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583",x"3ae3",x"404f",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"355a",x"3ae3",x"404b",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"3555"),
(x"3ae3",x"404b",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"3555",x"3ae3",x"404f",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"355a",x"3ae3",x"404b",x"abe1",x"3c00",x"0000",x"0000",x"2c5b",x"3555"),
(x"3ae3",x"3d85",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"32ee",x"3ae3",x"3d84",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"32ed",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1"),
(x"3ae3",x"3d92",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"32fe",x"3ae3",x"3d84",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"32ed",x"3ae3",x"3d85",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"32ee"),
(x"3ae3",x"3d92",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"32fe",x"3ae3",x"3d92",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"32fe",x"3ae3",x"3d84",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"32ed"),
(x"3ae3",x"404b",x"abe1",x"3c00",x"0000",x"0000",x"2c5b",x"3555",x"3ae3",x"3d92",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"32fe",x"3ae3",x"404b",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"3555"),
(x"3aad",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"3ad0",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1",x"3aad",x"3d46",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"2cc3"),
(x"3aad",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337",x"3ad4",x"404f",x"2ce6",x"0000",x"0000",x"3c00",x"316c",x"32dd",x"3ad0",x"404a",x"2ce6",x"0000",x"0000",x"3c00",x"316f",x"32d1"),
(x"3ae3",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"3337",x"3ae3",x"4056",x"2ce6",x"0000",x"0000",x"3c00",x"3162",x"32f1",x"3aad",x"4070",x"2ce6",x"0000",x"0000",x"3c00",x"3187",x"3337"),
(x"3ae3",x"3d92",x"2c35",x"3a20",x"184d",x"3924",x"31f3",x"3363",x"3ae3",x"3d85",x"2c89",x"39d0",x"342d",x"3915",x"31f9",x"3351",x"3ad1",x"3d90",x"2ce6",x"3a4a",x"1ef6",x"38f1",x"3206",x"3362"),
(x"3ae3",x"404b",x"2c40",x"39f4",x"9af6",x"3957",x"31f3",x"35b7",x"3ae3",x"3d92",x"2c35",x"3a20",x"184d",x"3924",x"31f3",x"3363",x"3ad0",x"404a",x"2ce6",x"3a20",x"935f",x"3925",x"3206",x"35b6"),
(x"3ae3",x"404e",x"2c57",x"39db",x"b485",x"38f4",x"31f4",x"35bc",x"3ae3",x"404b",x"2c40",x"39f4",x"9af6",x"3957",x"31f3",x"35b7",x"3ad4",x"404f",x"2ce6",x"39e5",x"b3cd",x"390b",x"3204",x"35bc"),
(x"3ad2",x"3507",x"b515",x"3a7c",x"38ae",x"1c81",x"3204",x"2c67",x"3ad6",x"3507",x"b544",x"3a14",x"38d9",x"337c",x"3214",x"2c6a",x"3ae3",x"34dc",x"b522",x"3a50",x"38e8",x"2604",x"3209",x"2c8b"),
(x"3ad4",x"3506",x"b075",x"3aa1",x"3878",x"a594",x"310b",x"2c66",x"3ad2",x"3507",x"b515",x"3a7c",x"38ae",x"1c81",x"3204",x"2c67",x"3ae3",x"34d8",x"b07b",x"3a7d",x"38ad",x"9e59",x"310c",x"2c8b"),
(x"3ada",x"3506",x"b010",x"3a5f",x"3855",x"b446",x"30f9",x"2c6a",x"3ad4",x"3506",x"b075",x"3aa1",x"3878",x"a594",x"310b",x"2c66",x"3ae3",x"34eb",x"b00e",x"3a6d",x"3864",x"b364",x"30f9",x"2c80"),
(x"3ad4",x"3506",x"b075",x"249b",x"3bff",x"1418",x"2d42",x"23ef",x"3aad",x"3507",x"aca4",x"1d38",x"3c00",x"8cea",x"2c87",x"224e",x"3ad2",x"3507",x"b515",x"1f10",x"3c00",x"1018",x"2f35",x"23e3"),
(x"3aad",x"3507",x"aca4",x"1d38",x"3c00",x"8cea",x"2c87",x"224e",x"3ae3",x"3507",x"af74",x"9f79",x"3c00",x"9c81",x"2d02",x"244a",x"3ae3",x"3507",x"aca4",x"0000",x"3c00",x"8000",x"2c87",x"244a"),
(x"3ad4",x"3506",x"b075",x"249b",x"3bff",x"1418",x"2d42",x"23ef",x"3ada",x"3506",x"b010",x"a0d0",x"3bff",x"a081",x"2d20",x"2418",x"3aad",x"3507",x"aca4",x"1d38",x"3c00",x"8cea",x"2c87",x"224e"),
(x"3aad",x"3cac",x"aca4",x"8e8d",x"bc00",x"8000",x"2392",x"2570",x"3ada",x"3cac",x"b010",x"0000",x"bc00",x"0000",x"262a",x"247f",x"3ad4",x"3cac",x"b075",x"0000",x"bc00",x"0000",x"26b4",x"249f"),
(x"3ae3",x"3cac",x"aca4",x"0000",x"bc00",x"0000",x"2392",x"244d",x"3ae3",x"3cac",x"af8a",x"0000",x"bc00",x"0000",x"25c3",x"244d",x"3aad",x"3cac",x"aca4",x"8e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"3ad4",x"3cac",x"b075",x"0000",x"bc00",x"0000",x"26b4",x"249f",x"3ad2",x"3cac",x"b515",x"928d",x"bc00",x"868d",x"2b3f",x"24a6",x"3aad",x"3cac",x"aca4",x"8e8d",x"bc00",x"8000",x"2392",x"2570"),
(x"3ac5",x"3638",x"b504",x"3a04",x"8000",x"b945",x"3140",x"336f",x"3ac5",x"3c5a",x"b504",x"3a04",x"8000",x"b945",x"3140",x"3598",x"3aad",x"35ff",x"b53c",x"3a04",x"8000",x"b945",x"3127",x"335c"),
(x"3aad",x"35ff",x"b032",x"3a0b",x"b93d",x"0000",x"30ea",x"2c2c",x"3ac5",x"3638",x"b0a7",x"3a0b",x"b93d",x"0000",x"30fe",x"2bf4",x"3aad",x"35ff",x"b53c",x"3a0b",x"b93d",x"0000",x"31fc",x"2c2c"),
(x"3aad",x"3c69",x"b032",x"3a1b",x"0000",x"392a",x"3106",x"35a2",x"3ac5",x"3c5a",x"b0a7",x"3a1b",x"0000",x"392a",x"30ec",x"3598",x"3aad",x"35ff",x"b032",x"3a1b",x"0000",x"392a",x"3106",x"335c"),
(x"3ada",x"3cac",x"b010",x"3a44",x"b877",x"b45c",x"244b",x"21c8",x"3ae3",x"3cb3",x"b00e",x"3a59",x"b87c",x"b388",x"2447",x"2120",x"3ad4",x"3cac",x"b075",x"3a96",x"b888",x"a5d6",x"24d8",x"21ed"),
(x"3ac5",x"3638",x"b504",x"3c00",x"0000",x"0000",x"26b9",x"330c",x"3ac5",x"3638",x"b0a7",x"3c00",x"0000",x"0000",x"2ac8",x"330c",x"3ac5",x"3c5a",x"b504",x"3c00",x"0000",x"0000",x"26b9",x"3545"),
(x"3aad",x"35ff",x"b032",x"3c00",x"0000",x"0000",x"3036",x"331b",x"3aad",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"32d0",x"3aad",x"3c69",x"b032",x"3c00",x"0000",x"0000",x"3036",x"354d"),
(x"3ad4",x"3cac",x"b075",x"3a96",x"b888",x"a5d6",x"24d8",x"21ed",x"3ae3",x"3cb8",x"b07b",x"3a76",x"b8b6",x"9fe2",x"24df",x"20ca",x"3ad2",x"3cac",x"b515",x"3a76",x"b8b6",x"1ac2",x"2a51",x"21ed"),
(x"3aad",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2ddb",x"32d0",x"3aad",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"32d0",x"3aad",x"35ff",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"331b"),
(x"3aad",x"3c69",x"b032",x"3c00",x"0000",x"0000",x"3036",x"354d",x"3aad",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"3080",x"3575",x"3aad",x"3c69",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"354d"),
(x"3aad",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2ddb",x"3575",x"3aad",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2ddb",x"32d0",x"3aad",x"3c69",x"b53c",x"3c00",x"0000",x"0000",x"2e82",x"354d"),
(x"3ad2",x"3cac",x"b515",x"3a76",x"b8b6",x"1ac2",x"2a51",x"21ed",x"3ae3",x"3cb7",x"b522",x"3a50",x"b8e8",x"25a8",x"2a63",x"20cc",x"3ad6",x"3cac",x"b544",x"3a14",x"b8d9",x"337c",x"2a90",x"21d6"),
(x"3ae3",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"2d4a",x"3aad",x"3507",x"b64e",x"0000",x"0000",x"3c00",x"322c",x"2d4a",x"3ae3",x"3cac",x"b64e",x"0000",x"0000",x"3c00",x"3207",x"333a"),
(x"3ae3",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"244a",x"3ae3",x"3507",x"b578",x"0000",x"3c00",x"8000",x"2f78",x"244a",x"3aad",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e"),
(x"3ad2",x"3507",x"b515",x"1f10",x"3c00",x"1018",x"2f35",x"23e3",x"3aad",x"3507",x"b64e",x"0000",x"3c00",x"8000",x"3005",x"224e",x"3ad6",x"3507",x"b544",x"0000",x"3c00",x"8000",x"2f54",x"2404"),
(x"3ae3",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2d4a",x"3ae3",x"35d5",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"2dd4",x"3aad",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"3ad0",x"3631",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"2e12",x"3aad",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a",x"3ad7",x"35fb",x"aca4",x"0000",x"8000",x"bc00",x"31fc",x"2dee"),
(x"3ac5",x"3c5a",x"b504",x"3a28",x"391a",x"0000",x"31e9",x"2a76",x"3ac5",x"3c5a",x"b0a7",x"3a28",x"391a",x"0000",x"30fe",x"2a76",x"3aad",x"3c69",x"b53c",x"3a28",x"391a",x"0000",x"31fc",x"2a0f"),
(x"3ae3",x"3cac",x"b64e",x"91bc",x"bc00",x"8000",x"2c74",x"244d",x"3aad",x"3cac",x"b64e",x"91bc",x"bc00",x"8000",x"2c74",x"2570",x"3ae3",x"3cac",x"b578",x"8e8d",x"bc00",x"8a8d",x"2bc6",x"244d"),
(x"3ad2",x"3cac",x"b515",x"928d",x"bc00",x"868d",x"2b3f",x"24a6",x"3ad6",x"3cac",x"b544",x"90ea",x"bc00",x"868d",x"2b7e",x"2492",x"3aad",x"3cac",x"b64e",x"91bc",x"bc00",x"8000",x"2c74",x"2570"),
(x"3ad0",x"3631",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"2e12",x"3ad0",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"3aad",x"3507",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"2d4a"),
(x"3aad",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a",x"3ae3",x"3c7a",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"32f6",x"3ae3",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"3203",x"333a"),
(x"3ad0",x"3c61",x"aca4",x"0000",x"8000",x"bc00",x"31f7",x"32d5",x"3ad3",x"3c6a",x"aca4",x"0000",x"8000",x"bc00",x"31f9",x"32e0",x"3aad",x"3cac",x"aca4",x"0000",x"8000",x"bc00",x"31de",x"333a"),
(x"3ad7",x"35fb",x"aca4",x"39a1",x"3488",x"b935",x"320d",x"3350",x"3ae3",x"35fe",x"ac3b",x"39ce",x"340f",x"b91d",x"3219",x"3351",x"3ad0",x"3631",x"aca4",x"3a39",x"1e59",x"b906",x"320a",x"3363"),
(x"3ad0",x"3631",x"aca4",x"3a39",x"1e59",x"b906",x"320a",x"3363",x"3ae3",x"3635",x"abd9",x"3a32",x"1818",x"b90f",x"321e",x"3364",x"3ad0",x"3c61",x"aca4",x"3a32",x"95bc",x"b90f",x"320a",x"3597"),
(x"3ae3",x"3c61",x"abe1",x"3a2a",x"97c8",x"b918",x"321e",x"3597",x"3ae3",x"3c6a",x"ac0f",x"39ea",x"b3b0",x"b908",x"321c",x"359d",x"3ad0",x"3c61",x"aca4",x"3a32",x"95bc",x"b90f",x"320a",x"3597"),
(x"3ad2",x"3506",x"351f",x"3a5d",x"38d8",x"9f93",x"2b9a",x"1c77",x"3ae3",x"34db",x"3523",x"3a4f",x"38ea",x"a57a",x"2b95",x"1ec7",x"3ad8",x"3505",x"3551",x"3a36",x"38b3",x"b345",x"2b55",x"1cd0"),
(x"3ad2",x"3506",x"307d",x"3a66",x"38cb",x"2460",x"2dc4",x"1c77",x"3ae3",x"34d8",x"3099",x"3a5b",x"38da",x"1d38",x"2dba",x"1ed9",x"3ad2",x"3506",x"351f",x"3a5d",x"38d8",x"9f93",x"2b9a",x"1c77"),
(x"3ad7",x"3506",x"302e",x"3a14",x"38b9",x"3455",x"2ddf",x"1cb4",x"3ae3",x"34e8",x"3026",x"3a1b",x"38d7",x"3338",x"2de2",x"1e54",x"3ad2",x"3506",x"307d",x"3a66",x"38cb",x"2460",x"2dc4",x"1c77"),
(x"3ad2",x"3506",x"307d",x"23e2",x"3bff",x"8cea",x"2f4d",x"2652",x"3ad2",x"3506",x"351f",x"2259",x"3bff",x"068d",x"2d56",x"2651",x"3aad",x"3507",x"2ce6",x"2067",x"3c00",x"1018",x"2fff",x"258a"),
(x"3aad",x"3507",x"2ce6",x"2067",x"3c00",x"1018",x"2fff",x"258a",x"3ad7",x"3506",x"302e",x"a032",x"3bff",x"2025",x"2f68",x"266a",x"3ad2",x"3506",x"307d",x"23e2",x"3bff",x"8cea",x"2f4d",x"2652"),
(x"3ae3",x"3507",x"2ce6",x"0000",x"3c00",x"8000",x"2fff",x"26ad",x"3ae3",x"3507",x"2f74",x"9ea7",x"3c00",x"1c67",x"2f8f",x"26ad",x"3aad",x"3507",x"2ce6",x"2067",x"3c00",x"1018",x"2fff",x"258a"),
(x"3aad",x"3cac",x"2ce6",x"8e8d",x"bc00",x"8000",x"2fff",x"27de",x"3ae3",x"3cac",x"2f82",x"0000",x"bc00",x"0000",x"2f8d",x"26bb",x"3ae3",x"3cac",x"2ce6",x"0000",x"bc00",x"0000",x"2fff",x"26bb"),
(x"3ad4",x"3cac",x"3071",x"0000",x"bc00",x"0000",x"2f51",x"270e",x"3ada",x"3cac",x"300c",x"0000",x"bc00",x"0000",x"2f73",x"26ed",x"3aad",x"3cac",x"2ce6",x"8e8d",x"bc00",x"8000",x"2fff",x"27de"),
(x"3ad4",x"3cac",x"3071",x"0000",x"bc00",x"0000",x"2f51",x"270e",x"3aad",x"3cac",x"2ce6",x"8e8d",x"bc00",x"8000",x"2fff",x"27de",x"3ad2",x"3cac",x"3524",x"928d",x"bc00",x"068d",x"2d52",x"2714"),
(x"3ac5",x"3639",x"3513",x"3a04",x"0000",x"3945",x"3144",x"3370",x"3aad",x"3600",x"354b",x"3a04",x"0000",x"3945",x"315d",x"335c",x"3ac5",x"3c5a",x"3513",x"3a04",x"0000",x"3945",x"3144",x"3597"),
(x"3ac5",x"3639",x"3513",x"3a0f",x"b938",x"0000",x"30fd",x"2c30",x"3ac5",x"3639",x"30dd",x"3a0f",x"b938",x"0000",x"31e4",x"2c30",x"3aad",x"3600",x"354b",x"3a0f",x"b938",x"0000",x"30ea",x"2c62"),
(x"3ac5",x"3639",x"30dd",x"3a15",x"8000",x"b931",x"3123",x"3370",x"3ac5",x"3c5a",x"30dd",x"3a15",x"8000",x"b931",x"3123",x"3597",x"3aad",x"3600",x"3069",x"3a15",x"8000",x"b931",x"3109",x"335c"),
(x"3ada",x"3cac",x"300c",x"3a44",x"b877",x"345c",x"2deb",x"2088",x"3ad4",x"3cac",x"3071",x"3a96",x"b888",x"25b5",x"2dc8",x"20ad",x"3ae3",x"3cb3",x"300a",x"3a59",x"b87c",x"3388",x"2dec",x"1fbf"),
(x"3ac5",x"3639",x"3513",x"3c00",x"0000",x"0000",x"3028",x"3323",x"3ac5",x"3c5a",x"3513",x"3c00",x"0000",x"0000",x"3028",x"3547",x"3ac5",x"3639",x"30dd",x"3c00",x"0000",x"0000",x"2eaa",x"3323"),
(x"3aad",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"3573",x"3aad",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"32b8",x"3aad",x"3c69",x"3069",x"3c00",x"0000",x"0000",x"2658",x"354a"),
(x"3ad4",x"3cac",x"3071",x"3a96",x"b888",x"25b5",x"2dc8",x"20ad",x"3ad2",x"3cac",x"3524",x"3a76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"3ae3",x"3cb8",x"3076",x"3a77",x"b8b5",x"1f93",x"2dc6",x"1f14"),
(x"3aad",x"3507",x"364e",x"3c00",x"0000",x"0000",x"2c23",x"32b8",x"3aad",x"3600",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"3304",x"3aad",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"32b8"),
(x"3aad",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"2c23",x"3573",x"3aad",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"23ce",x"3573",x"3aad",x"3c69",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"354a"),
(x"3aad",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"2c23",x"3573",x"3aad",x"3c69",x"354b",x"3c00",x"0000",x"0000",x"2b04",x"354a",x"3aad",x"3507",x"364e",x"3c00",x"0000",x"0000",x"2c23",x"32b8"),
(x"3ad2",x"3cac",x"3524",x"3a76",x"b8b6",x"9a8d",x"2b93",x"20ab",x"3ad6",x"3cac",x"3553",x"3a14",x"b8d9",x"b37c",x"2b54",x"2093",x"3ae3",x"3cb7",x"3532",x"3a50",x"b8e8",x"a587",x"2b82",x"1f14"),
(x"3aad",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"318d",x"333a",x"3aad",x"3507",x"364e",x"0000",x"8000",x"bc00",x"318d",x"2d4a",x"3ae3",x"3cac",x"364e",x"0000",x"8000",x"bc00",x"31b2",x"333a"),
(x"3ae3",x"3507",x"364e",x"0000",x"3c00",x"8000",x"2c87",x"26ad",x"3aad",x"3507",x"364e",x"1e0a",x"3c00",x"91bc",x"2c87",x"258a",x"3ae3",x"3507",x"3587",x"a04d",x"3c00",x"9cb5",x"2d0f",x"26ad"),
(x"3ad2",x"3506",x"351f",x"2259",x"3bff",x"068d",x"2d56",x"2651",x"3ad8",x"3505",x"3551",x"94ea",x"3c00",x"9dd6",x"2d34",x"2673",x"3aad",x"3507",x"364e",x"1e0a",x"3c00",x"91bc",x"2c87",x"258a"),
(x"3ae3",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2d4a",x"3aad",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a",x"3ae3",x"35d7",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"2dd5"),
(x"3ad1",x"3630",x"2ce6",x"0000",x"0000",x"3c00",x"31c2",x"2e11",x"3ad9",x"35fd",x"2ce6",x"0000",x"0000",x"3c00",x"31bd",x"2def",x"3aad",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"3ac5",x"3c5a",x"3513",x"3a28",x"391a",x"0000",x"30fd",x"2bed",x"3aad",x"3c69",x"354b",x"3a28",x"391a",x"0000",x"30ea",x"2b85",x"3ac5",x"3c5a",x"30dd",x"3a28",x"391a",x"0000",x"31e4",x"2bed"),
(x"3ae3",x"3cac",x"364e",x"91bc",x"bc00",x"8000",x"2c87",x"26bb",x"3ae3",x"3cac",x"3587",x"8e8d",x"bc00",x"0a8d",x"2d0f",x"26bb",x"3aad",x"3cac",x"364e",x"91bc",x"bc00",x"8000",x"2c87",x"27de"),
(x"3ad2",x"3cac",x"3524",x"928d",x"bc00",x"068d",x"2d52",x"2714",x"3aad",x"3cac",x"364e",x"91bc",x"bc00",x"8000",x"2c87",x"27de",x"3ad6",x"3cac",x"3553",x"8a8d",x"bc00",x"0cea",x"2d33",x"2701"),
(x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0",x"3ae3",x"35fe",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"2c0f",x"3ae3",x"35d5",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2beb"),
(x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0",x"3ae3",x"35fe",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"2c0f",x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"3ae3",x"35d7",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2bee",x"3ae3",x"3601",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"2c10",x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0"),
(x"3ae3",x"3c61",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"318b",x"3ae3",x"3635",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"2c30",x"3ae3",x"3635",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"2c30"),
(x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3c6a",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"3195",x"3ae3",x"3c61",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"318b"),
(x"3ae3",x"3c61",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"318b",x"3ae3",x"3c6a",x"ac0f",x"3c00",x"0000",x"0000",x"2c56",x"3195",x"3ae3",x"3c61",x"abe1",x"3c00",x"0000",x"0000",x"2c5b",x"318b"),
(x"3ae3",x"3601",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"2c10",x"3ae3",x"35fe",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"2c0f",x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0"),
(x"3ae3",x"3635",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"2c30",x"3ae3",x"35fe",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"2c0f",x"3ae3",x"3601",x"2c89",x"3c00",x"0000",x"0000",x"2dbb",x"2c10"),
(x"3ae3",x"3635",x"2c35",x"3c00",x"0000",x"0000",x"2dad",x"2c30",x"3ae3",x"3635",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"2c30",x"3ae3",x"35fe",x"ac3b",x"3c00",x"0000",x"0000",x"2c4f",x"2c0f"),
(x"3ae3",x"3c61",x"abe1",x"3c00",x"0000",x"0000",x"2c5b",x"318b",x"3ae3",x"3635",x"abd9",x"3c00",x"0000",x"0000",x"2c5c",x"2c30",x"3ae3",x"3c61",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"318b"),
(x"3aad",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"3ad0",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4",x"3aad",x"3507",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"2d4a"),
(x"3aad",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a",x"3ad4",x"3c69",x"2ce6",x"0000",x"0000",x"3c00",x"31c0",x"32e0",x"3ad0",x"3c60",x"2ce6",x"0000",x"0000",x"3c00",x"31c3",x"32d4"),
(x"3ae3",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"333a",x"3ae3",x"3c78",x"2ce6",x"0000",x"0000",x"3c00",x"31b6",x"32f4",x"3aad",x"3cac",x"2ce6",x"0000",x"0000",x"3c00",x"31db",x"333a"),
(x"3ae3",x"3635",x"2c35",x"3a20",x"1881",x"3924",x"3221",x"3363",x"3ae3",x"3601",x"2c89",x"39d0",x"342d",x"3915",x"3227",x"3351",x"3ad1",x"3630",x"2ce6",x"3a4a",x"1f5f",x"38f1",x"3235",x"3362"),
(x"3ae3",x"3c61",x"2c40",x"39f4",x"9b5f",x"3957",x"3221",x"3597",x"3ae3",x"3635",x"2c35",x"3a20",x"1881",x"3924",x"3221",x"3363",x"3ad0",x"3c60",x"2ce6",x"3a20",x"9418",x"3925",x"3234",x"3596"),
(x"3ae3",x"3c69",x"2c57",x"39db",x"b485",x"38f4",x"3223",x"359c",x"3ae3",x"3c61",x"2c40",x"39f4",x"9b5f",x"3957",x"3221",x"3597",x"3ad4",x"3c69",x"2ce6",x"39e5",x"b3cc",x"390b",x"3233",x"359c"),
(x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0",x"3ae3",x"34e8",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"2acb",x"3ae3",x"3507",x"2f74",x"3c00",x"0000",x"0000",x"2e33",x"2af0"),
(x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f",x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0"),
(x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0",x"3ae3",x"34d8",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"2ab8",x"3ae3",x"34e8",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"2acb"),
(x"3ae3",x"3507",x"af74",x"3c00",x"0000",x"0000",x"2b94",x"2af0",x"3ae3",x"34eb",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"2acf",x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"3ae3",x"34eb",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"2acf",x"3ae3",x"34d8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"2ab8",x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"3ae3",x"3507",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"2af0",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f",x"3ae3",x"34d8",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"2ab8"),
(x"3ae3",x"34d8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"2ab8",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c",x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0"),
(x"3ae3",x"3507",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"2af0",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"3507",x"b578",x"3c00",x"0000",x"0000",x"25d1",x"2af0",x"3ae3",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"2af0",x"3ae3",x"34f4",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"2ad9"),
(x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c",x"3ae3",x"34f4",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"2ad9",x"3ae3",x"3507",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"2af0"),
(x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c",x"3ae3",x"34d8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"2ab8",x"3ae3",x"34dc",x"b522",x"3c00",x"0000",x"0000",x"26af",x"2abd"),
(x"3ae3",x"3507",x"3587",x"3c00",x"0000",x"0000",x"3049",x"2af0",x"3ae3",x"34ea",x"3554",x"3c00",x"0000",x"0000",x"3039",x"2ace",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"34ea",x"3554",x"3c00",x"0000",x"0000",x"3039",x"2ace",x"3ae3",x"34db",x"3523",x"3c00",x"0000",x"0000",x"3029",x"2abb",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"34f4",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"2ad9",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c",x"3ae3",x"34dc",x"b522",x"3c00",x"0000",x"0000",x"26af",x"2abd"),
(x"3ae3",x"0000",x"364d",x"3c00",x"0000",x"0000",x"3089",x"1e82",x"3ae3",x"0000",x"3753",x"3c00",x"0000",x"0000",x"30de",x"1e82",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"3507",x"3587",x"3c00",x"0000",x"0000",x"3049",x"2af0",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f",x"3ae3",x"3507",x"364e",x"3c00",x"0000",x"0000",x"308a",x"2af0"),
(x"3ae3",x"3227",x"3753",x"3c00",x"0000",x"0000",x"30de",x"2890",x"3ae3",x"3507",x"364e",x"3c00",x"0000",x"0000",x"308a",x"2af0",x"3ae3",x"3154",x"364d",x"3c00",x"0000",x"0000",x"3089",x"280f"),
(x"3ae3",x"4062",x"3753",x"3c00",x"0000",x"0000",x"30de",x"3572",x"3ae3",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"308a",x"31e6",x"3ae3",x"3227",x"3753",x"3c00",x"0000",x"0000",x"30de",x"2890"),
(x"3ae3",x"3227",x"3753",x"3c00",x"0000",x"0000",x"30de",x"2890",x"3ae3",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"308a",x"31e6",x"3ae3",x"3507",x"364e",x"3c00",x"0000",x"0000",x"308a",x"2af0"),
(x"3ae3",x"4070",x"364e",x"3c00",x"0000",x"0000",x"308a",x"3583",x"3ae3",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"308a",x"32a1",x"3ae3",x"4062",x"3753",x"3c00",x"0000",x"0000",x"30de",x"3572"),
(x"3ae3",x"3d46",x"3587",x"3c00",x"0000",x"0000",x"3049",x"32a1",x"3ae3",x"3d3e",x"3554",x"3c00",x"0000",x"0000",x"3039",x"3298",x"3ae3",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"308a",x"32a1"),
(x"3ae3",x"3d3e",x"3554",x"3c00",x"0000",x"0000",x"3039",x"3298",x"3ae3",x"3cb1",x"3569",x"3c00",x"0000",x"0000",x"3040",x"31ec",x"3ae3",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"308a",x"32a1"),
(x"3ae3",x"3d3a",x"3523",x"3c00",x"0000",x"0000",x"3029",x"3293",x"3ae3",x"3cb7",x"3532",x"3c00",x"0000",x"0000",x"302e",x"31f3",x"3ae3",x"3d3e",x"3554",x"3c00",x"0000",x"0000",x"3039",x"3298"),
(x"3ae3",x"3cac",x"3587",x"3c00",x"0000",x"0000",x"3049",x"31e6",x"3ae3",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"308a",x"31e6",x"3ae3",x"3cb1",x"3569",x"3c00",x"0000",x"0000",x"3040",x"31ec"),
(x"3ae3",x"4062",x"3753",x"3c00",x"0000",x"0000",x"30de",x"3572",x"3ae3",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"308a",x"32a1",x"3ae3",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"308a",x"31e6"),
(x"3ae3",x"3cb1",x"3569",x"3c00",x"0000",x"0000",x"3040",x"31ec",x"3ae3",x"3d3e",x"3554",x"3c00",x"0000",x"0000",x"3039",x"3298",x"3ae3",x"3cb7",x"3532",x"3c00",x"0000",x"0000",x"302e",x"31f3"),
(x"3ae3",x"3cac",x"364e",x"3c00",x"0000",x"0000",x"308a",x"31e6",x"3ae3",x"3d46",x"364e",x"3c00",x"0000",x"0000",x"308a",x"32a1",x"3ae3",x"3cb1",x"3569",x"3c00",x"0000",x"0000",x"3040",x"31ec"),
(x"3ae3",x"3cb7",x"3532",x"3c00",x"0000",x"0000",x"302e",x"31f3",x"3ae3",x"3d3a",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"3293",x"3ae3",x"3cb8",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"31f4"),
(x"3ae3",x"3d3a",x"3523",x"3c00",x"0000",x"0000",x"3029",x"3293",x"3ae3",x"3d3a",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"3293",x"3ae3",x"3cb7",x"3532",x"3c00",x"0000",x"0000",x"302e",x"31f3"),
(x"3ae3",x"3cac",x"2f82",x"3c00",x"0000",x"0000",x"2e36",x"31e6",x"3ae3",x"3cb3",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"31ee",x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6"),
(x"3ae3",x"3cb8",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"31f4",x"3ae3",x"3d3e",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"3297",x"3ae3",x"3cb3",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"31ee"),
(x"3ae3",x"3d3a",x"3099",x"3c00",x"0000",x"0000",x"2e7c",x"3293",x"3ae3",x"3d3e",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"3297",x"3ae3",x"3cb8",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"31f4"),
(x"3ae3",x"3d46",x"2f74",x"3c00",x"0000",x"0000",x"2e33",x"32a1",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1",x"3ae3",x"3d3e",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"3297"),
(x"3ae3",x"3c78",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31a6",x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6",x"3ae3",x"3c69",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"3194"),
(x"3ae3",x"3cb3",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"31ee",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1",x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6"),
(x"3ae3",x"3d3e",x"3026",x"3c00",x"0000",x"0000",x"2e57",x"3297",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1",x"3ae3",x"3cb3",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"31ee"),
(x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1",x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6",x"3ae3",x"3d46",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"32a1"),
(x"3ae3",x"3d46",x"af74",x"3c00",x"0000",x"0000",x"2b94",x"32a1",x"3ae3",x"3d3f",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3298",x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"3ae3",x"3d3f",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3298",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1"),
(x"3ae3",x"3d3a",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"3293",x"3ae3",x"3cb8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"31f4",x"3ae3",x"3d3f",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3298"),
(x"3ae3",x"3c69",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"3194",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3c61",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"318b"),
(x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3c69",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"3194"),
(x"3ae3",x"3cac",x"af8a",x"3c00",x"0000",x"0000",x"2b8d",x"31e6",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3cb3",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"31ee"),
(x"3ae3",x"3d46",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"32a1",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3cac",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"31e6"),
(x"3ae3",x"3cb8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"31f4",x"3ae3",x"3cb3",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"31ee",x"3ae3",x"3d3f",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3298"),
(x"3ae3",x"3cb3",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"31ee",x"3ae3",x"3cac",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"31e6",x"3ae3",x"3d3f",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3298"),
(x"3ae3",x"3d3b",x"b522",x"3c00",x"0000",x"0000",x"26af",x"3294",x"3ae3",x"3cb7",x"b522",x"3c00",x"0000",x"0000",x"26af",x"31f3",x"3ae3",x"3d3a",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"3293"),
(x"3ae3",x"3d3a",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"3293",x"3ae3",x"3cb7",x"b522",x"3c00",x"0000",x"0000",x"26af",x"31f3",x"3ae3",x"3cb8",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"31f4"),
(x"3ae3",x"3d46",x"b578",x"3c00",x"0000",x"0000",x"25d1",x"32a1",x"3ae3",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"32a1",x"3ae3",x"3d41",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"329b"),
(x"3ae3",x"3d3b",x"b522",x"3c00",x"0000",x"0000",x"26af",x"3294",x"3ae3",x"3cb1",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"31ec",x"3ae3",x"3cb7",x"b522",x"3c00",x"0000",x"0000",x"26af",x"31f3"),
(x"3ae3",x"3d41",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"329b",x"3ae3",x"3cb1",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"31ec",x"3ae3",x"3d3b",x"b522",x"3c00",x"0000",x"0000",x"26af",x"3294"),
(x"3ae3",x"3cac",x"b578",x"3c00",x"0000",x"0000",x"25d1",x"31e6",x"3ae3",x"3cb1",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"31ec",x"3ae3",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"31e6"),
(x"3ae3",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"32a1",x"3ae3",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"31e6",x"3ae3",x"3d41",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"329b"),
(x"3ae3",x"3154",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"280f",x"3ae3",x"8000",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"1e82",x"3ae3",x"314f",x"b64f",x"3c00",x"0000",x"0000",x"234a",x"280c"),
(x"3ae3",x"4062",x"3753",x"3c00",x"0000",x"0000",x"30de",x"3572",x"3ae3",x"408e",x"3753",x"3c00",x"0000",x"0000",x"30de",x"35a7",x"3ae3",x"4070",x"364e",x"3c00",x"0000",x"0000",x"308a",x"3583"),
(x"3ae3",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"3583",x"3ae3",x"4073",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"3586",x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7"),
(x"3ae3",x"4070",x"b578",x"3c00",x"0000",x"0000",x"25d1",x"3583",x"3ae3",x"4073",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"3586",x"3ae3",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"3583"),
(x"3ae3",x"4070",x"364e",x"3c00",x"0000",x"0000",x"308a",x"3583",x"3ae3",x"4073",x"3569",x"3c00",x"0000",x"0000",x"3040",x"3586",x"3ae3",x"4070",x"3587",x"3c00",x"0000",x"0000",x"3049",x"3583"),
(x"3ae3",x"408e",x"3753",x"3c00",x"0000",x"0000",x"30de",x"35a7",x"3ae3",x"4073",x"3569",x"3c00",x"0000",x"0000",x"3040",x"3586",x"3ae3",x"4070",x"364e",x"3c00",x"0000",x"0000",x"308a",x"3583"),
(x"3ae3",x"4073",x"b55a",x"3c00",x"0000",x"0000",x"261e",x"3586",x"3ae3",x"4076",x"b522",x"3c00",x"0000",x"0000",x"26af",x"3589",x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7"),
(x"3ae3",x"4076",x"b522",x"3c00",x"0000",x"0000",x"26af",x"3589",x"3ae3",x"4076",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"358a",x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7"),
(x"3ae3",x"4073",x"3569",x"3c00",x"0000",x"0000",x"3040",x"3586",x"3ae3",x"408e",x"3753",x"3c00",x"0000",x"0000",x"30de",x"35a7",x"3ae3",x"4076",x"3532",x"3c00",x"0000",x"0000",x"302e",x"3589"),
(x"3ae3",x"4076",x"3532",x"3c00",x"0000",x"0000",x"302e",x"3589",x"3ae3",x"408e",x"3753",x"3c00",x"0000",x"0000",x"30de",x"35a7",x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a"),
(x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7",x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a",x"3ae3",x"408e",x"3753",x"3c00",x"0000",x"0000",x"30de",x"35a7"),
(x"3ae3",x"4076",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"358a",x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a",x"3ae3",x"408e",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"35a7"),
(x"3ae3",x"4070",x"af8a",x"3c00",x"0000",x"0000",x"2b8d",x"3583",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583",x"3ae3",x"4073",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3587"),
(x"3ae3",x"4073",x"b00e",x"3c00",x"0000",x"0000",x"2b5d",x"3587",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583",x"3ae3",x"4076",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"358a"),
(x"3ae3",x"4076",x"b07b",x"3c00",x"0000",x"0000",x"2b17",x"358a",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583",x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a"),
(x"3ae3",x"404b",x"2c40",x"3c00",x"0000",x"0000",x"2daf",x"3555",x"3ae3",x"404e",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"355a",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583"),
(x"3ae3",x"4070",x"2f82",x"3c00",x"0000",x"0000",x"2e36",x"3583",x"3ae3",x"4073",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"3587",x"3ae3",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3583"),
(x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a",x"3ae3",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3583",x"3ae3",x"4073",x"300a",x"3c00",x"0000",x"0000",x"2e4d",x"3587"),
(x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583",x"3ae3",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3583",x"3ae3",x"4076",x"3076",x"3c00",x"0000",x"0000",x"2e71",x"358a"),
(x"3ae3",x"404e",x"2c57",x"3c00",x"0000",x"0000",x"2db3",x"355a",x"3ae3",x"4070",x"2ce6",x"3c00",x"0000",x"0000",x"2dca",x"3583",x"3ae3",x"4070",x"aca4",x"3c00",x"0000",x"0000",x"2c3e",x"3583"),
(x"3ae3",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"32a1",x"3ae3",x"4070",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"3583",x"3ae3",x"3d42",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"329d"),
(x"3ae3",x"3cac",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"31e6",x"3ae3",x"3d46",x"b64e",x"3c00",x"0000",x"0000",x"2351",x"32a1",x"3ae3",x"3cb5",x"b751",x"3c00",x"0000",x"0000",x"1c22",x"31f0"),
(x"ba24",x"3d17",x"b69f",x"baa3",x"3877",x"8a8d",x"3820",x"360d",x"ba22",x"3d1b",x"b69c",x"bbe0",x"3192",x"868d",x"381a",x"360e",x"ba24",x"3d17",x"3793",x"bab4",x"385d",x"0000",x"3820",x"381b"),
(x"ba22",x"3d1b",x"3791",x"adff",x"3bf6",x"1c32",x"3821",x"35db",x"ba22",x"3d1b",x"b69c",x"ae6e",x"3bf5",x"8000",x"3823",x"3361",x"ba0f",x"3d1c",x"3751",x"ae0a",x"3bf6",x"1b93",x"3826",x"35cd"),
(x"ba73",x"3cfa",x"b73d",x"bb54",x"b669",x"068d",x"3847",x"35de",x"ba72",x"3cfe",x"b739",x"bb04",x"37ae",x"0a8d",x"3840",x"35e1",x"ba73",x"3cf9",x"381a",x"bb62",x"b628",x"8cea",x"3846",x"3833"),
(x"ba72",x"3cfe",x"b739",x"bb04",x"37ae",x"0a8d",x"3840",x"35e1",x"ba66",x"3d02",x"b720",x"b74f",x"3b1d",x"8000",x"3839",x"35eb",x"ba73",x"3cfd",x"3819",x"ba34",x"390d",x"8e8d",x"3840",x"3833"),
(x"ba6d",x"3cf5",x"3814",x"b8f1",x"ba4a",x"8a8d",x"384d",x"3830",x"ba69",x"3cf4",x"b72a",x"b902",x"ba3c",x"8000",x"384e",x"35e5",x"ba73",x"3cf9",x"381a",x"bb62",x"b628",x"8cea",x"3846",x"3833"),
(x"ba6c",x"3d01",x"3812",x"b7d0",x"3afb",x"8e8d",x"3839",x"382f",x"ba66",x"3d02",x"b720",x"b74f",x"3b1d",x"8000",x"3839",x"35eb",x"ba59",x"3d04",x"37fb",x"b62b",x"3b61",x"868d",x"3832",x"3829"),
(x"ba57",x"3cee",x"b704",x"b85c",x"bab4",x"0a8d",x"3854",x"35ee",x"ba69",x"3cf4",x"b72a",x"b902",x"ba3c",x"8000",x"384e",x"35e5",x"ba59",x"3cef",x"3800",x"b852",x"babb",x"0a8d",x"3854",x"382c"),
(x"ba59",x"3d04",x"37fb",x"b62b",x"3b61",x"868d",x"3832",x"3829",x"ba51",x"3d06",x"b6f9",x"b6de",x"3b39",x"8000",x"3833",x"35f5",x"ba3f",x"3d0b",x"37cd",x"b82f",x"3ad1",x"8000",x"382c",x"3824"),
(x"ba45",x"3ce8",x"b6e1",x"b8fd",x"ba41",x"8000",x"385a",x"35f7",x"ba57",x"3cee",x"b704",x"b85c",x"bab4",x"0a8d",x"3854",x"35ee",x"ba48",x"3ce9",x"37dc",x"b8b5",x"ba78",x"8000",x"385a",x"3827"),
(x"ba3f",x"3d0b",x"37cd",x"b82f",x"3ad1",x"8000",x"382c",x"3824",x"ba3e",x"3d0b",x"b6d2",x"b8d1",x"3a62",x"0a8d",x"382c",x"35fe",x"ba2f",x"3d12",x"37ac",x"b96f",x"39de",x"0a8d",x"3826",x"3820"),
(x"ba31",x"3cdf",x"b6b8",x"b9a0",x"b9b0",x"0a8d",x"3860",x"35ff",x"ba45",x"3ce8",x"b6e1",x"b8fd",x"ba41",x"8000",x"385a",x"35f7",x"ba30",x"3cdf",x"37af",x"b96d",x"b9e0",x"068d",x"3861",x"3823"),
(x"ba2f",x"3d12",x"37ac",x"b96f",x"39de",x"0a8d",x"3826",x"3820",x"ba30",x"3d12",x"b6b5",x"b995",x"39ba",x"0a8d",x"3826",x"3606",x"ba24",x"3d17",x"3793",x"bab4",x"385d",x"0000",x"3820",x"381b"),
(x"ba1f",x"3cd6",x"b693",x"b9b2",x"b99d",x"0000",x"3867",x"3607",x"ba31",x"3cdf",x"b6b8",x"b9a0",x"b9b0",x"0a8d",x"3860",x"35ff",x"ba1e",x"3cd6",x"3788",x"b9be",x"b991",x"0a8d",x"3867",x"381f"),
(x"ba1e",x"3cd6",x"3788",x"b099",x"bbea",x"1e0a",x"3827",x"35c9",x"ba11",x"3cd5",x"374e",x"aca7",x"bbfa",x"1d04",x"382b",x"35b5",x"ba1f",x"3cd6",x"b693",x"ad09",x"bbf9",x"91bc",x"382a",x"3380"),
(x"ba73",x"3cfa",x"b73d",x"8000",x"b59f",x"bb7d",x"38b4",x"359e",x"ba11",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b4",x"3573",x"ba72",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b2",x"359d"),
(x"ba72",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b2",x"359d",x"ba11",x"3cfe",x"b739",x"0000",x"39e6",x"b967",x"38b1",x"3573",x"ba66",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38ae",x"3598"),
(x"ba11",x"3cf4",x"b72a",x"0000",x"ba78",x"b8b3",x"38b8",x"3573",x"ba11",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b4",x"3573",x"ba69",x"3cf4",x"b72a",x"0000",x"b9ee",x"b95e",x"38b8",x"3599"),
(x"ba66",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38ae",x"3598",x"ba11",x"3d02",x"b720",x"8000",x"3b4b",x"b68f",x"38ad",x"3573",x"ba51",x"3d06",x"b6f9",x"0000",x"3b4f",x"b67f",x"38a8",x"358f"),
(x"ba11",x"3cee",x"b704",x"8000",x"baba",x"b853",x"38bd",x"3573",x"ba11",x"3cf4",x"b72a",x"0000",x"ba78",x"b8b3",x"38b8",x"3573",x"ba57",x"3cee",x"b704",x"0000",x"bacf",x"b832",x"38be",x"3592"),
(x"ba51",x"3d06",x"b6f9",x"0000",x"3b4f",x"b67f",x"38a8",x"358f",x"ba11",x"3d06",x"b6f9",x"0000",x"3b21",x"b73f",x"38a8",x"3573",x"ba3e",x"3d0b",x"b6d2",x"0000",x"3ab8",x"b856",x"38a2",x"3587"),
(x"ba11",x"3ce8",x"b6e1",x"8000",x"ba3a",x"b904",x"38c3",x"3573",x"ba11",x"3cee",x"b704",x"8000",x"baba",x"b853",x"38bd",x"3573",x"ba45",x"3ce8",x"b6e1",x"8000",x"ba6e",x"b8c2",x"38c3",x"3589"),
(x"ba3e",x"3d0b",x"b6d2",x"0000",x"3ab8",x"b856",x"38a2",x"3587",x"ba11",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bd",x"38a2",x"3573",x"ba30",x"3d12",x"b6b5",x"8000",x"39f0",x"b95c",x"389d",x"3581"),
(x"ba11",x"3cdf",x"b6b8",x"0000",x"b9cc",x"b983",x"38ca",x"3573",x"ba11",x"3ce8",x"b6e1",x"8000",x"ba3a",x"b904",x"38c3",x"3573",x"ba31",x"3cdf",x"b6b8",x"0000",x"b9ea",x"b962",x"38ca",x"3581"),
(x"ba30",x"3d12",x"b6b5",x"8000",x"39f0",x"b95c",x"389d",x"3581",x"ba11",x"3d12",x"b6b5",x"0000",x"39c3",x"b98b",x"389d",x"3574",x"ba24",x"3d17",x"b69f",x"0000",x"38fa",x"ba43",x"3899",x"357c"),
(x"ba11",x"3cd6",x"b693",x"0000",x"b9a2",x"b9ad",x"38d1",x"3573",x"ba11",x"3cdf",x"b6b8",x"0000",x"b9cc",x"b983",x"38ca",x"3573",x"ba1f",x"3cd6",x"b693",x"0000",x"b9a2",x"b9ad",x"38d1",x"3579"),
(x"b9d3",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38d1",x"359f",x"b9d3",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38cf",x"359f",x"ba22",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38d1",x"35c1"),
(x"ba1e",x"3cd6",x"3788",x"b099",x"bbea",x"1e0a",x"3827",x"35c9",x"b9d3",x"3cd6",x"3788",x"0000",x"bbfa",x"2ca7",x"383d",x"35c7",x"ba11",x"3cd5",x"374e",x"aca7",x"bbfa",x"1d04",x"382b",x"35b5"),
(x"b9d3",x"3d1c",x"3751",x"0000",x"3bfc",x"2bc8",x"3833",x"35d2",x"b9d3",x"3d1b",x"3791",x"0000",x"3bfc",x"2bc8",x"3831",x"35dd",x"ba0f",x"3d1c",x"3751",x"ae0a",x"3bf6",x"1b93",x"3826",x"35cd"),
(x"ba73",x"3cfd",x"3819",x"8000",x"3707",x"3b2f",x"38b5",x"35e4",x"b9d3",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38b5",x"359f",x"ba73",x"3cf9",x"381a",x"0000",x"b15c",x"3be2",x"38b4",x"35e4"),
(x"b9d3",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b8",x"359f",x"b9d3",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38b5",x"359f",x"ba6c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b8",x"35e1"),
(x"ba73",x"3cf9",x"381a",x"0000",x"b15c",x"3be2",x"38b4",x"35e4",x"b9d3",x"3cf9",x"381a",x"868d",x"b62d",x"3b61",x"38b4",x"359f",x"ba6d",x"3cf5",x"3814",x"0000",x"b9d2",x"397b",x"38b1",x"35e1"),
(x"b9d3",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38be",x"359f",x"b9d3",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b8",x"359f",x"ba59",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38be",x"35d9"),
(x"ba6d",x"3cf5",x"3814",x"0000",x"b9d2",x"397b",x"38b1",x"35e1",x"b9d3",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38b1",x"359f",x"ba59",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38ab",x"35d9"),
(x"b9d3",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38c5",x"359f",x"b9d3",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38be",x"359f",x"ba3f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c5",x"35ce"),
(x"ba59",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38ab",x"35d9",x"b9d3",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38ab",x"359f",x"ba48",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a5",x"35d1"),
(x"b9d3",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38ca",x"359f",x"b9d3",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38c5",x"359f",x"ba2f",x"3d12",x"37ac",x"8000",x"3a00",x"3949",x"38ca",x"35c6"),
(x"ba48",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a5",x"35d1",x"b9d3",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"38a5",x"359f",x"ba30",x"3cdf",x"37af",x"0000",x"b9ed",x"395f",x"389e",x"35c7"),
(x"b9d3",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38cf",x"359f",x"b9d3",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38ca",x"359f",x"ba24",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cf",x"35c2"),
(x"ba30",x"3cdf",x"37af",x"0000",x"b9ed",x"395f",x"389e",x"35c7",x"b9d3",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"389e",x"359f",x"ba1e",x"3cd6",x"3788",x"0000",x"b9c4",x"398a",x"3896",x"35bf"),
(x"b94c",x"3d2f",x"364c",x"0000",x"3c00",x"1818",x"3819",x"3833",x"3a1b",x"3d2f",x"364c",x"0000",x"3c00",x"1818",x"3819",x"34a2",x"b94c",x"3d2f",x"3730",x"868d",x"3bfc",x"2baa",x"3803",x"3833"),
(x"b94c",x"3cef",x"37de",x"8000",x"baca",x"383b",x"373b",x"3833",x"3a1b",x"3cef",x"37de",x"0000",x"bacd",x"3836",x"373b",x"3574",x"b94c",x"3ce9",x"37b9",x"0000",x"ba81",x"38a7",x"372b",x"3833"),
(x"b94c",x"3d04",x"37d8",x"0000",x"3b36",x"36eb",x"378a",x"3833",x"3a1b",x"3d04",x"37d8",x"0000",x"3b60",x"3632",x"378a",x"3575",x"b94c",x"3d01",x"3801",x"8000",x"3b45",x"36ac",x"377a",x"3833"),
(x"b94c",x"3ce9",x"37b9",x"0000",x"ba81",x"38a7",x"372b",x"3833",x"3a1b",x"3ce9",x"37b9",x"0000",x"ba3c",x"3903",x"372b",x"3574",x"b94c",x"3cdf",x"378c",x"0000",x"b9ec",x"3960",x"371b",x"3833"),
(x"b94c",x"3d17",x"3770",x"0000",x"3765",x"3b17",x"37b9",x"3833",x"3a1b",x"3d17",x"3770",x"0000",x"3916",x"3a2c",x"37b9",x"3576",x"b94c",x"3d12",x"3789",x"0000",x"39ed",x"395f",x"37a9",x"3833"),
(x"b94c",x"3cdf",x"378c",x"0000",x"b9ec",x"3960",x"371b",x"3833",x"3a1b",x"3cdf",x"378c",x"0000",x"b9d9",x"3975",x"371b",x"3574",x"b94c",x"3cd6",x"3765",x"068d",x"ba59",x"38de",x"370b",x"3833"),
(x"b94c",x"3d1b",x"376e",x"0000",x"3032",x"3bee",x"37c9",x"3833",x"3a1b",x"3d1b",x"376e",x"0000",x"3032",x"3bee",x"37c9",x"3576",x"b94c",x"3d17",x"3770",x"8000",x"3766",x"3b17",x"37b9",x"3833"),
(x"b94c",x"3cd6",x"3765",x"068d",x"ba59",x"38de",x"370b",x"3833",x"3a1b",x"3cd6",x"3765",x"8000",x"bb2c",x"3715",x"370b",x"3574",x"b94c",x"3cd5",x"374e",x"0000",x"bbf9",x"2d34",x"36fb",x"3832"),
(x"b94c",x"3d1c",x"374a",x"0000",x"3bfc",x"2b80",x"391b",x"3833",x"3a1b",x"3d1c",x"374a",x"0000",x"3bfc",x"2b80",x"391b",x"3578",x"b94c",x"3d1b",x"376e",x"0000",x"3bfc",x"2b80",x"3914",x"3833"),
(x"b94c",x"3d25",x"374a",x"0000",x"2fec",x"3bf0",x"37de",x"3833",x"3a1b",x"3d25",x"374a",x"0000",x"2907",x"3bfe",x"37de",x"34a1",x"b94c",x"3d1c",x"374a",x"0000",x"9e3f",x"3c00",x"37c9",x"3833"),
(x"b94c",x"3cfd",x"3807",x"0000",x"3838",x"3acb",x"376a",x"3833",x"3a1b",x"3cfd",x"3807",x"8000",x"3564",x"3b88",x"376a",x"3575",x"b94c",x"3cf9",x"3808",x"8000",x"b15f",x"3be2",x"375a",x"3833"),
(x"b94c",x"3d12",x"3789",x"0000",x"39ed",x"395f",x"37a9",x"3833",x"3a1b",x"3d12",x"3789",x"0000",x"39ff",x"394a",x"37a9",x"3575",x"b94c",x"3d0b",x"37aa",x"0000",x"3a78",x"38b4",x"3799",x"3833"),
(x"b94c",x"3d28",x"3746",x"8000",x"38ab",x"3a7e",x"37f2",x"3833",x"3a1b",x"3d28",x"3746",x"0000",x"3816",x"3ae0",x"37f2",x"34a1",x"b94c",x"3d25",x"374a",x"0000",x"2fec",x"3bf0",x"37de",x"3833"),
(x"b94c",x"3cf9",x"3808",x"8000",x"b15f",x"3be2",x"375a",x"3833",x"3a1b",x"3cf9",x"3808",x"0000",x"b636",x"3b5f",x"375a",x"3575",x"b94c",x"3cf5",x"3803",x"0000",x"b9d5",x"3979",x"374a",x"3833"),
(x"b94c",x"3d0b",x"37aa",x"0000",x"3a78",x"38b4",x"3799",x"3833",x"3a1b",x"3d0b",x"37aa",x"0000",x"3acc",x"3837",x"3799",x"3575",x"b94c",x"3d04",x"37d8",x"0000",x"3b36",x"36eb",x"378a",x"3833"),
(x"b94c",x"3d2f",x"3730",x"868d",x"3bfc",x"2baa",x"3803",x"3833",x"3a1b",x"3d2f",x"3730",x"0000",x"3bd6",x"3272",x"3803",x"34a2",x"b94c",x"3d28",x"3746",x"8000",x"38ab",x"3a7e",x"37f2",x"3833"),
(x"b94c",x"3cf5",x"3803",x"0000",x"b9d5",x"3979",x"374a",x"3833",x"3a1b",x"3cf5",x"3803",x"8000",x"ba74",x"38b9",x"374a",x"3574",x"b94c",x"3cef",x"37de",x"8000",x"baca",x"383b",x"373b",x"3833"),
(x"b94c",x"3d01",x"3801",x"8000",x"3b45",x"36ac",x"377a",x"3833",x"3a1b",x"3d01",x"3801",x"0000",x"3ab5",x"385c",x"377a",x"3575",x"b94c",x"3cfd",x"3807",x"0000",x"3838",x"3acb",x"376a",x"3833"),
(x"3af2",x"3d1b",x"3791",x"3bd8",x"324a",x"8000",x"38d5",x"381d",x"3af2",x"3d1b",x"b69c",x"3be0",x"3193",x"868d",x"38d4",x"3614",x"3af3",x"3d17",x"3793",x"3ab4",x"385d",x"0000",x"38d0",x"381e"),
(x"3aed",x"3cd6",x"3788",x"3099",x"bbea",x"1e0a",x"382d",x"35ae",x"3aee",x"3cd6",x"b693",x"312a",x"bbe5",x"8000",x"382f",x"3345",x"3ae0",x"3cd5",x"374e",x"30c7",x"bbe9",x"1da1",x"3831",x"359e"),
(x"3af2",x"3d1b",x"3791",x"2dff",x"3bf6",x"1c32",x"381b",x"35ee",x"3ade",x"3d1c",x"3751",x"2e0a",x"3bf6",x"1b93",x"3820",x"35de",x"3af2",x"3d1b",x"b69c",x"2e6e",x"3bf5",x"8000",x"381b",x"3359"),
(x"3b42",x"3cfd",x"3819",x"3a34",x"390d",x"8e8d",x"38b3",x"3833",x"3b41",x"3cfe",x"b739",x"3b04",x"37ae",x"0a8d",x"38b3",x"35ea",x"3b42",x"3cf9",x"381a",x"3b62",x"b628",x"8cea",x"38ad",x"3833"),
(x"3b3c",x"3d01",x"3812",x"37d0",x"3afb",x"8e8d",x"38b9",x"382f",x"3b35",x"3d02",x"b720",x"374f",x"3b1d",x"8000",x"38b9",x"35f3",x"3b42",x"3cfd",x"3819",x"3a34",x"390d",x"8e8d",x"38b3",x"3833"),
(x"3b3c",x"3cf5",x"3814",x"38f1",x"ba4a",x"8a8d",x"38a7",x"3831",x"3b42",x"3cf9",x"381a",x"3b62",x"b628",x"8cea",x"38ad",x"3833",x"3b38",x"3cf4",x"b72a",x"3902",x"ba3c",x"8000",x"38a7",x"35ee"),
(x"3b3c",x"3d01",x"3812",x"37d0",x"3afb",x"8e8d",x"38b9",x"382f",x"3b28",x"3d04",x"37fb",x"362b",x"3b61",x"868d",x"38bf",x"382a",x"3b35",x"3d02",x"b720",x"374f",x"3b1d",x"8000",x"38b9",x"35f3"),
(x"3b3c",x"3cf5",x"3814",x"38f1",x"ba4a",x"8a8d",x"38a7",x"3831",x"3b38",x"3cf4",x"b72a",x"3902",x"ba3c",x"8000",x"38a7",x"35ee",x"3b28",x"3cef",x"3800",x"3852",x"babb",x"0a8d",x"38a1",x"382c"),
(x"3b28",x"3d04",x"37fb",x"362b",x"3b61",x"868d",x"38bf",x"382a",x"3b0f",x"3d0b",x"37cd",x"382f",x"3ad1",x"8000",x"38c5",x"3826",x"3b20",x"3d06",x"b6f9",x"36de",x"3b39",x"8000",x"38bf",x"35fb"),
(x"3b28",x"3cef",x"3800",x"3852",x"babb",x"0a8d",x"38a1",x"382c",x"3b27",x"3cee",x"b704",x"385c",x"bab4",x"0a8d",x"38a1",x"35f8",x"3b17",x"3ce9",x"37dc",x"38b4",x"ba78",x"8000",x"389b",x"3828"),
(x"3b0f",x"3d0b",x"37cd",x"382f",x"3ad1",x"8000",x"38c5",x"3826",x"3afe",x"3d12",x"37ac",x"396f",x"39de",x"0a8d",x"38ca",x"3822",x"3b0d",x"3d0b",x"b6d2",x"38d1",x"3a62",x"0a8d",x"38c5",x"3604"),
(x"3b17",x"3ce9",x"37dc",x"38b4",x"ba78",x"8000",x"389b",x"3828",x"3b14",x"3ce8",x"b6e1",x"38fd",x"ba40",x"8000",x"389b",x"3600",x"3b00",x"3cdf",x"37af",x"396d",x"b9e0",x"068d",x"3896",x"3824"),
(x"3afe",x"3d12",x"37ac",x"396f",x"39de",x"0a8d",x"38ca",x"3822",x"3af3",x"3d17",x"3793",x"3ab4",x"385d",x"0000",x"38d0",x"381e",x"3aff",x"3d12",x"b6b5",x"3995",x"39ba",x"0a8d",x"38ca",x"360c"),
(x"3b00",x"3cdf",x"37af",x"396d",x"b9e0",x"068d",x"3896",x"3824",x"3b00",x"3cdf",x"b6b8",x"39a0",x"b9b0",x"0a8d",x"3896",x"3608",x"3aed",x"3cd6",x"3788",x"39be",x"b991",x"0a8d",x"3890",x"3820"),
(x"3ae0",x"3cd5",x"b68e",x"a724",x"b9b4",x"b99a",x"38d5",x"3513",x"3aee",x"3cd6",x"b693",x"a0c2",x"b9a8",x"b9a7",x"38d4",x"350c",x"3ae2",x"3cdf",x"b6b8",x"9da1",x"b9ce",x"b980",x"38cd",x"3512"),
(x"3b42",x"3cfa",x"b73d",x"8000",x"b59f",x"bb7d",x"38b6",x"34e0",x"3b41",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b3",x"34e1",x"3ae2",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b5",x"3512"),
(x"3b41",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b3",x"34e1",x"3b35",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38af",x"34e7",x"3ae2",x"3cfe",x"b739",x"0000",x"39e5",x"b967",x"38b3",x"3511"),
(x"3b42",x"3cfa",x"b73d",x"8000",x"b59f",x"bb7d",x"38b6",x"34e0",x"3ae2",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b5",x"3512",x"3b38",x"3cf4",x"b72a",x"8000",x"b9ed",x"b95e",x"38ba",x"34e6"),
(x"3b35",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38af",x"34e7",x"3b20",x"3d06",x"b6f9",x"8000",x"3b4f",x"b67e",x"38a9",x"34f1",x"3ae2",x"3d02",x"b720",x"0000",x"3b4b",x"b690",x"38ae",x"3511"),
(x"3b38",x"3cf4",x"b72a",x"8000",x"b9ed",x"b95e",x"38ba",x"34e6",x"3ae2",x"3cf4",x"b72a",x"8000",x"ba78",x"b8b4",x"38b9",x"3512",x"3b27",x"3cee",x"b704",x"8000",x"bacf",x"b832",x"38c0",x"34ef"),
(x"3b20",x"3d06",x"b6f9",x"8000",x"3b4f",x"b67e",x"38a9",x"34f1",x"3b0d",x"3d0b",x"b6d2",x"8000",x"3ab8",x"b856",x"38a3",x"34fb",x"3ae2",x"3d06",x"b6f9",x"8000",x"3b21",x"b73f",x"38a9",x"3511"),
(x"3b27",x"3cee",x"b704",x"8000",x"bacf",x"b832",x"38c0",x"34ef",x"3ae2",x"3cee",x"b704",x"0000",x"baba",x"b853",x"38bf",x"3512",x"3b14",x"3ce8",x"b6e1",x"0000",x"ba6e",x"b8c1",x"38c6",x"34f8"),
(x"3b0d",x"3d0b",x"b6d2",x"8000",x"3ab8",x"b856",x"38a3",x"34fb",x"3aff",x"3d12",x"b6b5",x"0000",x"39f0",x"b95c",x"389d",x"3502",x"3ae2",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bc",x"38a2",x"3511"),
(x"3b14",x"3ce8",x"b6e1",x"0000",x"ba6e",x"b8c1",x"38c6",x"34f8",x"3ae2",x"3ce8",x"b6e1",x"0000",x"ba3b",x"b904",x"38c5",x"3512",x"3b00",x"3cdf",x"b6b8",x"8000",x"b9ea",x"b962",x"38cd",x"3503"),
(x"3aff",x"3d12",x"b6b5",x"0000",x"39f0",x"b95c",x"389d",x"3502",x"3af3",x"3d17",x"b69f",x"0000",x"38fc",x"ba41",x"3899",x"3508",x"3ae2",x"3d12",x"b6b5",x"8000",x"39c4",x"b98b",x"389d",x"3511"),
(x"3af3",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cc",x"3545",x"3aa2",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38ca",x"3570",x"3af2",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38ce",x"3546"),
(x"3aed",x"3cd6",x"3788",x"3099",x"bbea",x"1e0a",x"382d",x"35ae",x"3ae0",x"3cd5",x"374e",x"30c7",x"bbe9",x"1da1",x"3831",x"359e",x"3aa2",x"3cd6",x"3788",x"0000",x"bbfa",x"2ca7",x"383d",x"35b3"),
(x"3af2",x"3d1b",x"3791",x"2dff",x"3bf6",x"1c32",x"381b",x"35ee",x"3aa2",x"3d1b",x"3791",x"0000",x"3bfc",x"2bc8",x"382e",x"35ef",x"3ade",x"3d1c",x"3751",x"2e0a",x"3bf6",x"1b93",x"3820",x"35de"),
(x"3b42",x"3cfd",x"3819",x"8000",x"3707",x"3b2f",x"38b4",x"351a",x"3b42",x"3cf9",x"381a",x"8000",x"b15d",x"3be2",x"38b2",x"351a",x"3aa2",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38af",x"356e"),
(x"3b42",x"3cfd",x"3819",x"8000",x"3707",x"3b2f",x"38b4",x"351a",x"3aa2",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38af",x"356e",x"3b3c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b7",x"351e"),
(x"3b42",x"3cf9",x"381a",x"8000",x"b15d",x"3be2",x"38b2",x"351a",x"3b3c",x"3cf5",x"3814",x"0000",x"b9d2",x"397c",x"38af",x"351d",x"3aa2",x"3cf9",x"381a",x"0000",x"b62d",x"3b61",x"38ad",x"356e"),
(x"3b3c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b7",x"351e",x"3aa2",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b2",x"356e",x"3b28",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38bc",x"3528"),
(x"3b3c",x"3cf5",x"3814",x"0000",x"b9d2",x"397c",x"38af",x"351d",x"3b28",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38a8",x"3527",x"3aa2",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38ab",x"356e"),
(x"3b28",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38bc",x"3528",x"3aa2",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38b8",x"356f",x"3b0f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c2",x"3536"),
(x"3b28",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38a8",x"3527",x"3b17",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a2",x"3530",x"3aa2",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38a4",x"356d"),
(x"3b0f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c2",x"3536",x"3aa2",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38bf",x"356f",x"3afe",x"3d12",x"37ac",x"8000",x"3a00",x"394a",x"38c8",x"353f"),
(x"3b17",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a2",x"3530",x"3b00",x"3cdf",x"37af",x"0000",x"b9ee",x"395e",x"3899",x"353b",x"3aa2",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"389f",x"356d"),
(x"3afe",x"3d12",x"37ac",x"8000",x"3a00",x"394a",x"38c8",x"353f",x"3aa2",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38c5",x"356f",x"3af3",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cc",x"3545"),
(x"3b00",x"3cdf",x"37af",x"0000",x"b9ee",x"395e",x"3899",x"353b",x"3aed",x"3cd6",x"3788",x"0000",x"b9c4",x"398b",x"3891",x"3544",x"3aa2",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"3897",x"356d"),
(x"3a1b",x"3cd5",x"374e",x"0000",x"0000",x"3c00",x"38fa",x"3381",x"3a1b",x"3cbf",x"374e",x"0000",x"0000",x"3c00",x"38ee",x"3381",x"b94c",x"3cd5",x"374e",x"0000",x"0000",x"3c00",x"38fa",x"3833"),
(x"3a1b",x"3cbf",x"374e",x"0000",x"bc00",x"0000",x"3907",x"33aa",x"3a1b",x"3cbf",x"36f7",x"0000",x"bc00",x"0000",x"38fa",x"33aa",x"b94c",x"3cbf",x"374e",x"0000",x"bc00",x"0000",x"3907",x"3833"),
(x"3a1b",x"3cbf",x"36f7",x"0000",x"8000",x"bc00",x"3913",x"33ac",x"3a1b",x"3cd5",x"36f7",x"0000",x"8000",x"bc00",x"3907",x"33ac",x"b94c",x"3cbf",x"36f7",x"0000",x"8000",x"bc00",x"3913",x"3833"),
(x"3a1b",x"3cd5",x"36f7",x"0000",x"bc00",x"0000",x"38ed",x"32f2",x"3a1b",x"3cd5",x"364d",x"0000",x"bc00",x"0000",x"38d7",x"32f2",x"b94c",x"3cd5",x"36f7",x"0000",x"bc00",x"0000",x"38ed",x"3833"),
(x"3a1b",x"3cd5",x"364d",x"0000",x"8000",x"bc00",x"388e",x"32f2",x"3a1b",x"3d1f",x"364d",x"0000",x"8000",x"bc00",x"3867",x"32f2",x"b94c",x"3cd5",x"364d",x"0000",x"8000",x"bc00",x"388e",x"3833"),
(x"ba24",x"3d17",x"b69f",x"0000",x"38fa",x"ba43",x"3899",x"357c",x"ba11",x"3d17",x"b69f",x"9c81",x"36c8",x"bb3e",x"3899",x"3574",x"ba22",x"3d1b",x"b69c",x"9ffc",x"30d9",x"bbe8",x"3897",x"357b"),
(x"3af3",x"3d17",x"b69f",x"0000",x"38fc",x"ba41",x"3899",x"3508",x"3af2",x"3d1b",x"b69c",x"2025",x"30de",x"bbe8",x"3896",x"3508",x"3ae2",x"3d17",x"b69f",x"1cb5",x"36b4",x"bb43",x"3899",x"3511"),
(x"ba22",x"3d1b",x"b69c",x"bbe0",x"3192",x"868d",x"381a",x"360e",x"ba22",x"3d1b",x"3791",x"bbd8",x"324a",x"8000",x"381a",x"381a",x"ba24",x"3d17",x"3793",x"bab4",x"385d",x"0000",x"3820",x"381b"),
(x"ba22",x"3d1b",x"b69c",x"ae6e",x"3bf5",x"8000",x"3823",x"3361",x"ba0f",x"3d1c",x"b69c",x"ae6e",x"3bf5",x"8000",x"3828",x"3361",x"ba0f",x"3d1c",x"3751",x"ae0a",x"3bf6",x"1b93",x"3826",x"35cd"),
(x"ba72",x"3cfe",x"b739",x"bb04",x"37ae",x"0a8d",x"3840",x"35e1",x"ba73",x"3cfd",x"3819",x"ba34",x"390d",x"8e8d",x"3840",x"3833",x"ba73",x"3cf9",x"381a",x"bb62",x"b628",x"8cea",x"3846",x"3833"),
(x"ba66",x"3d02",x"b720",x"b74f",x"3b1d",x"8000",x"3839",x"35eb",x"ba6c",x"3d01",x"3812",x"b7d0",x"3afb",x"8e8d",x"3839",x"382f",x"ba73",x"3cfd",x"3819",x"ba34",x"390d",x"8e8d",x"3840",x"3833"),
(x"ba69",x"3cf4",x"b72a",x"b902",x"ba3c",x"8000",x"384e",x"35e5",x"ba73",x"3cfa",x"b73d",x"bb54",x"b669",x"068d",x"3847",x"35de",x"ba73",x"3cf9",x"381a",x"bb62",x"b628",x"8cea",x"3846",x"3833"),
(x"ba66",x"3d02",x"b720",x"b74f",x"3b1d",x"8000",x"3839",x"35eb",x"ba51",x"3d06",x"b6f9",x"b6de",x"3b39",x"8000",x"3833",x"35f5",x"ba59",x"3d04",x"37fb",x"b62b",x"3b61",x"868d",x"3832",x"3829"),
(x"ba69",x"3cf4",x"b72a",x"b902",x"ba3c",x"8000",x"384e",x"35e5",x"ba6d",x"3cf5",x"3814",x"b8f1",x"ba4a",x"8a8d",x"384d",x"3830",x"ba59",x"3cef",x"3800",x"b852",x"babb",x"0a8d",x"3854",x"382c"),
(x"ba51",x"3d06",x"b6f9",x"b6de",x"3b39",x"8000",x"3833",x"35f5",x"ba3e",x"3d0b",x"b6d2",x"b8d1",x"3a62",x"0a8d",x"382c",x"35fe",x"ba3f",x"3d0b",x"37cd",x"b82f",x"3ad1",x"8000",x"382c",x"3824"),
(x"ba57",x"3cee",x"b704",x"b85c",x"bab4",x"0a8d",x"3854",x"35ee",x"ba59",x"3cef",x"3800",x"b852",x"babb",x"0a8d",x"3854",x"382c",x"ba48",x"3ce9",x"37dc",x"b8b5",x"ba78",x"8000",x"385a",x"3827"),
(x"ba3e",x"3d0b",x"b6d2",x"b8d1",x"3a62",x"0a8d",x"382c",x"35fe",x"ba30",x"3d12",x"b6b5",x"b995",x"39ba",x"0a8d",x"3826",x"3606",x"ba2f",x"3d12",x"37ac",x"b96f",x"39de",x"0a8d",x"3826",x"3820"),
(x"ba45",x"3ce8",x"b6e1",x"b8fd",x"ba41",x"8000",x"385a",x"35f7",x"ba48",x"3ce9",x"37dc",x"b8b5",x"ba78",x"8000",x"385a",x"3827",x"ba30",x"3cdf",x"37af",x"b96d",x"b9e0",x"068d",x"3861",x"3823"),
(x"ba30",x"3d12",x"b6b5",x"b995",x"39ba",x"0a8d",x"3826",x"3606",x"ba24",x"3d17",x"b69f",x"baa3",x"3877",x"8a8d",x"3820",x"360d",x"ba24",x"3d17",x"3793",x"bab4",x"385d",x"0000",x"3820",x"381b"),
(x"ba31",x"3cdf",x"b6b8",x"b9a0",x"b9b0",x"0a8d",x"3860",x"35ff",x"ba30",x"3cdf",x"37af",x"b96d",x"b9e0",x"068d",x"3861",x"3823",x"ba1e",x"3cd6",x"3788",x"b9be",x"b991",x"0a8d",x"3867",x"381f"),
(x"ba11",x"3cd5",x"374e",x"aca7",x"bbfa",x"1d04",x"382b",x"35b5",x"ba11",x"3cd6",x"b693",x"0000",x"bc00",x"9553",x"382e",x"337f",x"ba1f",x"3cd6",x"b693",x"ad09",x"bbf9",x"91bc",x"382a",x"3380"),
(x"ba11",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b4",x"3573",x"ba11",x"3cfe",x"b739",x"0000",x"39e6",x"b967",x"38b1",x"3573",x"ba72",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b2",x"359d"),
(x"ba11",x"3cfe",x"b739",x"0000",x"39e6",x"b967",x"38b1",x"3573",x"ba11",x"3d02",x"b720",x"8000",x"3b4b",x"b68f",x"38ad",x"3573",x"ba66",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38ae",x"3598"),
(x"ba11",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b4",x"3573",x"ba73",x"3cfa",x"b73d",x"8000",x"b59f",x"bb7d",x"38b4",x"359e",x"ba69",x"3cf4",x"b72a",x"0000",x"b9ee",x"b95e",x"38b8",x"3599"),
(x"ba11",x"3d02",x"b720",x"8000",x"3b4b",x"b68f",x"38ad",x"3573",x"ba11",x"3d06",x"b6f9",x"0000",x"3b21",x"b73f",x"38a8",x"3573",x"ba51",x"3d06",x"b6f9",x"0000",x"3b4f",x"b67f",x"38a8",x"358f"),
(x"ba11",x"3cf4",x"b72a",x"0000",x"ba78",x"b8b3",x"38b8",x"3573",x"ba69",x"3cf4",x"b72a",x"0000",x"b9ee",x"b95e",x"38b8",x"3599",x"ba57",x"3cee",x"b704",x"0000",x"bacf",x"b832",x"38be",x"3592"),
(x"ba11",x"3d06",x"b6f9",x"0000",x"3b21",x"b73f",x"38a8",x"3573",x"ba11",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bd",x"38a2",x"3573",x"ba3e",x"3d0b",x"b6d2",x"0000",x"3ab8",x"b856",x"38a2",x"3587"),
(x"ba11",x"3cee",x"b704",x"8000",x"baba",x"b853",x"38bd",x"3573",x"ba57",x"3cee",x"b704",x"0000",x"bacf",x"b832",x"38be",x"3592",x"ba45",x"3ce8",x"b6e1",x"8000",x"ba6e",x"b8c2",x"38c3",x"3589"),
(x"ba11",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bd",x"38a2",x"3573",x"ba11",x"3d12",x"b6b5",x"0000",x"39c3",x"b98b",x"389d",x"3574",x"ba30",x"3d12",x"b6b5",x"8000",x"39f0",x"b95c",x"389d",x"3581"),
(x"ba11",x"3ce8",x"b6e1",x"8000",x"ba3a",x"b904",x"38c3",x"3573",x"ba45",x"3ce8",x"b6e1",x"8000",x"ba6e",x"b8c2",x"38c3",x"3589",x"ba31",x"3cdf",x"b6b8",x"0000",x"b9ea",x"b962",x"38ca",x"3581"),
(x"ba11",x"3d12",x"b6b5",x"0000",x"39c3",x"b98b",x"389d",x"3574",x"ba11",x"3d17",x"b69f",x"9c81",x"36c8",x"bb3e",x"3899",x"3574",x"ba24",x"3d17",x"b69f",x"0000",x"38fa",x"ba43",x"3899",x"357c"),
(x"ba11",x"3cdf",x"b6b8",x"0000",x"b9cc",x"b983",x"38ca",x"3573",x"ba31",x"3cdf",x"b6b8",x"0000",x"b9ea",x"b962",x"38ca",x"3581",x"ba1f",x"3cd6",x"b693",x"0000",x"b9a2",x"b9ad",x"38d1",x"3579"),
(x"b9d3",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38cf",x"359f",x"ba24",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cf",x"35c2",x"ba22",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38d1",x"35c1"),
(x"b9d3",x"3cd6",x"3788",x"0000",x"bbfa",x"2ca7",x"383d",x"35c7",x"b9d3",x"3cd5",x"374e",x"0000",x"bbfa",x"2ca7",x"383d",x"35b4",x"ba11",x"3cd5",x"374e",x"aca7",x"bbfa",x"1d04",x"382b",x"35b5"),
(x"b9d3",x"3d1b",x"3791",x"0000",x"3bfc",x"2bc8",x"3831",x"35dd",x"ba22",x"3d1b",x"3791",x"adff",x"3bf6",x"1c32",x"3821",x"35db",x"ba0f",x"3d1c",x"3751",x"ae0a",x"3bf6",x"1b93",x"3826",x"35cd"),
(x"b9d3",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38b5",x"359f",x"b9d3",x"3cf9",x"381a",x"868d",x"b62d",x"3b61",x"38b4",x"359f",x"ba73",x"3cf9",x"381a",x"0000",x"b15c",x"3be2",x"38b4",x"35e4"),
(x"b9d3",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38b5",x"359f",x"ba73",x"3cfd",x"3819",x"8000",x"3707",x"3b2f",x"38b5",x"35e4",x"ba6c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b8",x"35e1"),
(x"b9d3",x"3cf9",x"381a",x"868d",x"b62d",x"3b61",x"38b4",x"359f",x"b9d3",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38b1",x"359f",x"ba6d",x"3cf5",x"3814",x"0000",x"b9d2",x"397b",x"38b1",x"35e1"),
(x"b9d3",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b8",x"359f",x"ba6c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b8",x"35e1",x"ba59",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38be",x"35d9"),
(x"b9d3",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38b1",x"359f",x"b9d3",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38ab",x"359f",x"ba59",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38ab",x"35d9"),
(x"b9d3",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38be",x"359f",x"ba59",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38be",x"35d9",x"ba3f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c5",x"35ce"),
(x"b9d3",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38ab",x"359f",x"b9d3",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"38a5",x"359f",x"ba48",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a5",x"35d1"),
(x"b9d3",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38c5",x"359f",x"ba3f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c5",x"35ce",x"ba2f",x"3d12",x"37ac",x"8000",x"3a00",x"3949",x"38ca",x"35c6"),
(x"b9d3",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"38a5",x"359f",x"b9d3",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"389e",x"359f",x"ba30",x"3cdf",x"37af",x"0000",x"b9ed",x"395f",x"389e",x"35c7"),
(x"b9d3",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38ca",x"359f",x"ba2f",x"3d12",x"37ac",x"8000",x"3a00",x"3949",x"38ca",x"35c6",x"ba24",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cf",x"35c2"),
(x"b9d3",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"389e",x"359f",x"b9d3",x"3cd6",x"3788",x"0000",x"b9c4",x"398b",x"3896",x"359f",x"ba1e",x"3cd6",x"3788",x"0000",x"b9c4",x"398a",x"3896",x"35bf"),
(x"3a1b",x"3d2f",x"364c",x"0000",x"3c00",x"1818",x"3819",x"34a2",x"3a1b",x"3d2f",x"3730",x"0000",x"3bd6",x"3272",x"3803",x"34a2",x"b94c",x"3d2f",x"3730",x"868d",x"3bfc",x"2baa",x"3803",x"3833"),
(x"3a1b",x"3cef",x"37de",x"0000",x"bacd",x"3836",x"373b",x"3574",x"3a1b",x"3ce9",x"37b9",x"0000",x"ba3c",x"3903",x"372b",x"3574",x"b94c",x"3ce9",x"37b9",x"0000",x"ba81",x"38a7",x"372b",x"3833"),
(x"3a1b",x"3d04",x"37d8",x"0000",x"3b60",x"3632",x"378a",x"3575",x"3a1b",x"3d01",x"3801",x"0000",x"3ab5",x"385c",x"377a",x"3575",x"b94c",x"3d01",x"3801",x"8000",x"3b45",x"36ac",x"377a",x"3833"),
(x"3a1b",x"3ce9",x"37b9",x"0000",x"ba3c",x"3903",x"372b",x"3574",x"3a1b",x"3cdf",x"378c",x"0000",x"b9d9",x"3975",x"371b",x"3574",x"b94c",x"3cdf",x"378c",x"0000",x"b9ec",x"3960",x"371b",x"3833"),
(x"3a1b",x"3d17",x"3770",x"0000",x"3916",x"3a2c",x"37b9",x"3576",x"3a1b",x"3d12",x"3789",x"0000",x"39ff",x"394a",x"37a9",x"3575",x"b94c",x"3d12",x"3789",x"0000",x"39ed",x"395f",x"37a9",x"3833"),
(x"3a1b",x"3cdf",x"378c",x"0000",x"b9d9",x"3975",x"371b",x"3574",x"3a1b",x"3cd6",x"3765",x"8000",x"bb2c",x"3715",x"370b",x"3574",x"b94c",x"3cd6",x"3765",x"068d",x"ba59",x"38de",x"370b",x"3833"),
(x"3a1b",x"3d1b",x"376e",x"0000",x"3032",x"3bee",x"37c9",x"3576",x"3a1b",x"3d17",x"3770",x"0000",x"3916",x"3a2c",x"37b9",x"3576",x"b94c",x"3d17",x"3770",x"0000",x"3765",x"3b17",x"37b9",x"3833"),
(x"3a1b",x"3cd6",x"3765",x"8000",x"bb2c",x"3716",x"370b",x"3574",x"3a1b",x"3cd5",x"374e",x"0000",x"bbf9",x"2d35",x"36fb",x"3574",x"b94c",x"3cd5",x"374e",x"0000",x"bbf9",x"2d35",x"36fb",x"3832"),
(x"3a1b",x"3d1c",x"374a",x"0000",x"3bfc",x"2b80",x"391b",x"3578",x"3a1b",x"3d1b",x"376e",x"0000",x"3bfc",x"2b80",x"3914",x"3578",x"b94c",x"3d1b",x"376e",x"0000",x"3bfc",x"2b80",x"3914",x"3833"),
(x"3a1b",x"3d25",x"374a",x"8000",x"290b",x"3bfe",x"37de",x"34a1",x"3a1b",x"3d1c",x"374a",x"0000",x"9e3f",x"3c00",x"37c9",x"34a1",x"b94c",x"3d1c",x"374a",x"0000",x"9e3f",x"3c00",x"37c9",x"3833"),
(x"3a1b",x"3cfd",x"3807",x"8000",x"3564",x"3b88",x"376a",x"3575",x"3a1b",x"3cf9",x"3808",x"0000",x"b636",x"3b5f",x"375a",x"3575",x"b94c",x"3cf9",x"3808",x"8000",x"b15f",x"3be2",x"375a",x"3833"),
(x"3a1b",x"3d12",x"3789",x"0000",x"39ff",x"394a",x"37a9",x"3575",x"3a1b",x"3d0b",x"37aa",x"0000",x"3acc",x"3837",x"3799",x"3575",x"b94c",x"3d0b",x"37aa",x"0000",x"3a78",x"38b4",x"3799",x"3833"),
(x"3a1b",x"3d28",x"3746",x"0000",x"3816",x"3ae0",x"37f2",x"34a1",x"3a1b",x"3d25",x"374a",x"0000",x"2907",x"3bfe",x"37de",x"34a1",x"b94c",x"3d25",x"374a",x"0000",x"2fec",x"3bf0",x"37de",x"3833"),
(x"3a1b",x"3cf9",x"3808",x"0000",x"b636",x"3b5f",x"375a",x"3575",x"3a1b",x"3cf5",x"3803",x"8000",x"ba74",x"38b9",x"374a",x"3574",x"b94c",x"3cf5",x"3803",x"0000",x"b9d5",x"3979",x"374a",x"3833"),
(x"3a1b",x"3d0b",x"37aa",x"0000",x"3acc",x"3837",x"3799",x"3575",x"3a1b",x"3d04",x"37d8",x"0000",x"3b60",x"3632",x"378a",x"3575",x"b94c",x"3d04",x"37d8",x"0000",x"3b36",x"36eb",x"378a",x"3833"),
(x"3a1b",x"3d2f",x"3730",x"0000",x"3bd6",x"3272",x"3803",x"34a2",x"3a1b",x"3d28",x"3746",x"0000",x"3816",x"3ae0",x"37f2",x"34a1",x"b94c",x"3d28",x"3746",x"8000",x"38ab",x"3a7e",x"37f2",x"3833"),
(x"3a1b",x"3cf5",x"3803",x"8000",x"ba74",x"38b9",x"374a",x"3574",x"3a1b",x"3cef",x"37de",x"0000",x"bacd",x"3836",x"373b",x"3574",x"b94c",x"3cef",x"37de",x"8000",x"baca",x"383b",x"373b",x"3833"),
(x"3a1b",x"3d01",x"3801",x"0000",x"3ab5",x"385c",x"377a",x"3575",x"3a1b",x"3cfd",x"3807",x"8000",x"3564",x"3b88",x"376a",x"3575",x"b94c",x"3cfd",x"3807",x"0000",x"3838",x"3acb",x"376a",x"3833"),
(x"3af2",x"3d1b",x"b69c",x"3be0",x"3193",x"868d",x"38d4",x"3614",x"3af3",x"3d17",x"b69f",x"3aa3",x"3877",x"8a8d",x"38cf",x"3612",x"3af3",x"3d17",x"3793",x"3ab4",x"385d",x"0000",x"38d0",x"381e"),
(x"3aee",x"3cd6",x"b693",x"312a",x"bbe5",x"8000",x"382f",x"3345",x"3ae0",x"3cd5",x"b68e",x"3151",x"bbe3",x"0000",x"3833",x"3349",x"3ae0",x"3cd5",x"374e",x"30c7",x"bbe9",x"1da1",x"3831",x"359e"),
(x"3ade",x"3d1c",x"3751",x"2e0a",x"3bf6",x"1b93",x"3820",x"35de",x"3ade",x"3d1c",x"b69c",x"2e6e",x"3bf5",x"8000",x"3820",x"3359",x"3af2",x"3d1b",x"b69c",x"2e6e",x"3bf5",x"8000",x"381b",x"3359"),
(x"3b41",x"3cfe",x"b739",x"3b04",x"37ae",x"0a8d",x"38b3",x"35ea",x"3b42",x"3cfa",x"b73d",x"3b54",x"b66a",x"068d",x"38ad",x"35e7",x"3b42",x"3cf9",x"381a",x"3b62",x"b628",x"8cea",x"38ad",x"3833"),
(x"3b35",x"3d02",x"b720",x"374f",x"3b1d",x"8000",x"38b9",x"35f3",x"3b41",x"3cfe",x"b739",x"3b04",x"37ae",x"0a8d",x"38b3",x"35ea",x"3b42",x"3cfd",x"3819",x"3a34",x"390d",x"8e8d",x"38b3",x"3833"),
(x"3b42",x"3cf9",x"381a",x"3b62",x"b628",x"8cea",x"38ad",x"3833",x"3b42",x"3cfa",x"b73d",x"3b54",x"b66a",x"068d",x"38ad",x"35e7",x"3b38",x"3cf4",x"b72a",x"3902",x"ba3c",x"8000",x"38a7",x"35ee"),
(x"3b28",x"3d04",x"37fb",x"362b",x"3b61",x"868d",x"38bf",x"382a",x"3b20",x"3d06",x"b6f9",x"36de",x"3b39",x"8000",x"38bf",x"35fb",x"3b35",x"3d02",x"b720",x"374f",x"3b1d",x"8000",x"38b9",x"35f3"),
(x"3b38",x"3cf4",x"b72a",x"3902",x"ba3c",x"8000",x"38a7",x"35ee",x"3b27",x"3cee",x"b704",x"385c",x"bab4",x"0a8d",x"38a1",x"35f8",x"3b28",x"3cef",x"3800",x"3852",x"babb",x"0a8d",x"38a1",x"382c"),
(x"3b0f",x"3d0b",x"37cd",x"382f",x"3ad1",x"8000",x"38c5",x"3826",x"3b0d",x"3d0b",x"b6d2",x"38d1",x"3a62",x"0a8d",x"38c5",x"3604",x"3b20",x"3d06",x"b6f9",x"36de",x"3b39",x"8000",x"38bf",x"35fb"),
(x"3b27",x"3cee",x"b704",x"385c",x"bab4",x"0a8d",x"38a1",x"35f8",x"3b14",x"3ce8",x"b6e1",x"38fd",x"ba40",x"8000",x"389b",x"3600",x"3b17",x"3ce9",x"37dc",x"38b4",x"ba78",x"8000",x"389b",x"3828"),
(x"3afe",x"3d12",x"37ac",x"396f",x"39de",x"0a8d",x"38ca",x"3822",x"3aff",x"3d12",x"b6b5",x"3995",x"39ba",x"0a8d",x"38ca",x"360c",x"3b0d",x"3d0b",x"b6d2",x"38d1",x"3a62",x"0a8d",x"38c5",x"3604"),
(x"3b14",x"3ce8",x"b6e1",x"38fd",x"ba40",x"8000",x"389b",x"3600",x"3b00",x"3cdf",x"b6b8",x"39a0",x"b9b0",x"0a8d",x"3896",x"3608",x"3b00",x"3cdf",x"37af",x"396d",x"b9e0",x"068d",x"3896",x"3824"),
(x"3af3",x"3d17",x"3793",x"3ab4",x"385d",x"0000",x"38d0",x"381e",x"3af3",x"3d17",x"b69f",x"3aa3",x"3877",x"8a8d",x"38cf",x"3612",x"3aff",x"3d12",x"b6b5",x"3995",x"39ba",x"0a8d",x"38ca",x"360c"),
(x"3b00",x"3cdf",x"b6b8",x"39a0",x"b9b0",x"0a8d",x"3896",x"3608",x"3aee",x"3cd6",x"b693",x"39b2",x"b99d",x"0000",x"3890",x"360f",x"3aed",x"3cd6",x"3788",x"39be",x"b991",x"0a8d",x"3890",x"3820"),
(x"3aee",x"3cd6",x"b693",x"a0c2",x"b9a8",x"b9a7",x"38d4",x"350c",x"3b00",x"3cdf",x"b6b8",x"8000",x"b9ea",x"b962",x"38cd",x"3503",x"3ae2",x"3cdf",x"b6b8",x"9da1",x"b9ce",x"b980",x"38cd",x"3512"),
(x"3b41",x"3cfe",x"b739",x"8000",x"385f",x"bab2",x"38b3",x"34e1",x"3ae2",x"3cfe",x"b739",x"0000",x"39e5",x"b967",x"38b3",x"3511",x"3ae2",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b5",x"3512"),
(x"3b35",x"3d02",x"b720",x"0000",x"3b16",x"b76b",x"38af",x"34e7",x"3ae2",x"3d02",x"b720",x"0000",x"3b4b",x"b690",x"38ae",x"3511",x"3ae2",x"3cfe",x"b739",x"0000",x"39e5",x"b967",x"38b3",x"3511"),
(x"3ae2",x"3cfa",x"b73d",x"0000",x"b575",x"bb85",x"38b5",x"3512",x"3ae2",x"3cf4",x"b72a",x"8000",x"ba78",x"b8b4",x"38b9",x"3512",x"3b38",x"3cf4",x"b72a",x"8000",x"b9ed",x"b95e",x"38ba",x"34e6"),
(x"3b20",x"3d06",x"b6f9",x"8000",x"3b4f",x"b67e",x"38a9",x"34f1",x"3ae2",x"3d06",x"b6f9",x"8000",x"3b21",x"b73f",x"38a9",x"3511",x"3ae2",x"3d02",x"b720",x"0000",x"3b4b",x"b690",x"38ae",x"3511"),
(x"3ae2",x"3cf4",x"b72a",x"8000",x"ba78",x"b8b4",x"38b9",x"3512",x"3ae2",x"3cee",x"b704",x"0000",x"baba",x"b853",x"38bf",x"3512",x"3b27",x"3cee",x"b704",x"8000",x"bacf",x"b832",x"38c0",x"34ef"),
(x"3b0d",x"3d0b",x"b6d2",x"8000",x"3ab8",x"b856",x"38a3",x"34fb",x"3ae2",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bc",x"38a2",x"3511",x"3ae2",x"3d06",x"b6f9",x"8000",x"3b21",x"b73f",x"38a9",x"3511"),
(x"3ae2",x"3cee",x"b704",x"0000",x"baba",x"b853",x"38bf",x"3512",x"3ae2",x"3ce8",x"b6e1",x"0000",x"ba3b",x"b904",x"38c5",x"3512",x"3b14",x"3ce8",x"b6e1",x"0000",x"ba6e",x"b8c1",x"38c6",x"34f8"),
(x"3aff",x"3d12",x"b6b5",x"0000",x"39f0",x"b95c",x"389d",x"3502",x"3ae2",x"3d12",x"b6b5",x"8000",x"39c4",x"b98b",x"389d",x"3511",x"3ae2",x"3d0b",x"b6d2",x"0000",x"3a72",x"b8bc",x"38a2",x"3511"),
(x"3ae2",x"3ce8",x"b6e1",x"0000",x"ba3b",x"b904",x"38c5",x"3512",x"3ae2",x"3cdf",x"b6b8",x"9da1",x"b9ce",x"b980",x"38cd",x"3512",x"3b00",x"3cdf",x"b6b8",x"8000",x"b9ea",x"b962",x"38cd",x"3503"),
(x"3af3",x"3d17",x"b69f",x"0000",x"38fc",x"ba41",x"3899",x"3508",x"3ae2",x"3d17",x"b69f",x"1cb5",x"36b4",x"bb43",x"3899",x"3511",x"3ae2",x"3d12",x"b6b5",x"8000",x"39c4",x"b98b",x"389d",x"3511"),
(x"3aa2",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38ca",x"3570",x"3aa2",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38cc",x"3570",x"3af2",x"3d1b",x"3791",x"0000",x"3031",x"3bee",x"38ce",x"3546"),
(x"3ae0",x"3cd5",x"374e",x"30c7",x"bbe9",x"1da1",x"3831",x"359e",x"3aa2",x"3cd5",x"374e",x"0000",x"bbfa",x"2ca7",x"383e",x"35a5",x"3aa2",x"3cd6",x"3788",x"0000",x"bbfa",x"2ca7",x"383d",x"35b3"),
(x"3aa2",x"3d1b",x"3791",x"0000",x"3bfc",x"2bc8",x"382e",x"35ef",x"3aa2",x"3d1c",x"3751",x"0000",x"3bfc",x"2bc8",x"382e",x"35de",x"3ade",x"3d1c",x"3751",x"2e0a",x"3bf6",x"1b93",x"3820",x"35de"),
(x"3b42",x"3cf9",x"381a",x"8000",x"b15d",x"3be2",x"38b2",x"351a",x"3aa2",x"3cf9",x"381a",x"0000",x"b62d",x"3b61",x"38ad",x"356e",x"3aa2",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38af",x"356e"),
(x"3aa2",x"3cfd",x"3819",x"0000",x"36fb",x"3b32",x"38af",x"356e",x"3aa2",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b2",x"356e",x"3b3c",x"3d01",x"3812",x"0000",x"3ab1",x"3860",x"38b7",x"351e"),
(x"3b3c",x"3cf5",x"3814",x"0000",x"b9d2",x"397c",x"38af",x"351d",x"3aa2",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38ab",x"356e",x"3aa2",x"3cf9",x"381a",x"0000",x"b62d",x"3b61",x"38ad",x"356e"),
(x"3aa2",x"3d01",x"3812",x"0000",x"3b41",x"36be",x"38b2",x"356e",x"3aa2",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38b8",x"356f",x"3b28",x"3d04",x"37fb",x"8000",x"3b62",x"3628",x"38bc",x"3528"),
(x"3b28",x"3cef",x"3800",x"0000",x"bac9",x"383b",x"38a8",x"3527",x"3aa2",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38a4",x"356d",x"3aa2",x"3cf5",x"3814",x"0000",x"ba6f",x"38c0",x"38ab",x"356e"),
(x"3aa2",x"3d04",x"37fb",x"0000",x"3b39",x"36df",x"38b8",x"356f",x"3aa2",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38bf",x"356f",x"3b0f",x"3d0b",x"37cd",x"8000",x"3ad1",x"382f",x"38c2",x"3536"),
(x"3b17",x"3ce9",x"37dc",x"8000",x"ba85",x"38a2",x"38a2",x"3530",x"3aa2",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"389f",x"356d",x"3aa2",x"3cef",x"3800",x"0000",x"bacd",x"3836",x"38a4",x"356d"),
(x"3aa2",x"3d0b",x"37cd",x"8000",x"3a7d",x"38ad",x"38bf",x"356f",x"3aa2",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38c5",x"356f",x"3afe",x"3d12",x"37ac",x"8000",x"3a00",x"394a",x"38c8",x"353f"),
(x"3b00",x"3cdf",x"37af",x"0000",x"b9ee",x"395e",x"3899",x"353b",x"3aa2",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"3897",x"356d",x"3aa2",x"3ce9",x"37dc",x"0000",x"ba40",x"38fd",x"389f",x"356d"),
(x"3aa2",x"3d12",x"37ac",x"0000",x"39ed",x"395e",x"38c5",x"356f",x"3aa2",x"3d17",x"3793",x"0000",x"376c",x"3b16",x"38ca",x"3570",x"3af3",x"3d17",x"3793",x"8000",x"3921",x"3a23",x"38cc",x"3545"),
(x"3aed",x"3cd6",x"3788",x"0000",x"b9c4",x"398b",x"3891",x"3544",x"3aa2",x"3cd6",x"3788",x"0000",x"b9c4",x"398b",x"388f",x"356c",x"3aa2",x"3cdf",x"37af",x"0000",x"b9da",x"3973",x"3897",x"356d"),
(x"3a1b",x"3cbf",x"374e",x"0000",x"0000",x"3c00",x"38ee",x"3381",x"b94c",x"3cbf",x"374e",x"0000",x"0000",x"3c00",x"38ee",x"3833",x"b94c",x"3cd5",x"374e",x"0000",x"0000",x"3c00",x"38fa",x"3833"),
(x"3a1b",x"3cbf",x"36f7",x"0000",x"bc00",x"0000",x"38fa",x"33aa",x"b94c",x"3cbf",x"36f7",x"0000",x"bc00",x"0000",x"38fa",x"3833",x"b94c",x"3cbf",x"374e",x"0000",x"bc00",x"0000",x"3907",x"3833"),
(x"3a1b",x"3cd5",x"36f7",x"0000",x"8000",x"bc00",x"3907",x"33ac",x"b94c",x"3cd5",x"36f7",x"0000",x"8000",x"bc00",x"3907",x"3833",x"b94c",x"3cbf",x"36f7",x"0000",x"8000",x"bc00",x"3913",x"3833"),
(x"3a1b",x"3cd5",x"364d",x"0000",x"bc00",x"0000",x"38d7",x"32f2",x"b94c",x"3cd5",x"364d",x"0000",x"bc00",x"0000",x"38d7",x"3833",x"b94c",x"3cd5",x"36f7",x"0000",x"bc00",x"0000",x"38ed",x"3833"),
(x"3a1b",x"3d1f",x"364d",x"0000",x"8000",x"bc00",x"3867",x"32f2",x"b94c",x"3d1f",x"364d",x"0000",x"8000",x"bc00",x"3867",x"3833",x"b94c",x"3cd5",x"364d",x"0000",x"8000",x"bc00",x"388e",x"3833"),
(x"ba11",x"3d17",x"b69f",x"9c81",x"36c8",x"bb3e",x"3899",x"3574",x"ba0f",x"3d1c",x"b69c",x"a32b",x"306c",x"bbec",x"3896",x"3573",x"ba22",x"3d1b",x"b69c",x"9ffc",x"30d9",x"bbe8",x"3897",x"357b"),
(x"3af2",x"3d1b",x"b69c",x"2025",x"30de",x"bbe8",x"3896",x"3508",x"3ade",x"3d1c",x"b69c",x"2345",x"307d",x"bbeb",x"3896",x"3512",x"3ae2",x"3d17",x"b69f",x"1cb5",x"36b4",x"bb43",x"3899",x"3511"),
(x"b9f6",x"4000",x"377d",x"b5fa",x"3ae9",x"3563",x"3641",x"34e8",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5",x"b9f7",x"3ffd",x"3794",x"b663",x"3a38",x"37c6",x"363b",x"34f0"),
(x"b9f6",x"4000",x"377d",x"b5fa",x"3ae9",x"3563",x"3641",x"34e8",x"ba00",x"3ffd",x"377a",x"b865",x"3a42",x"34ab",x"3647",x"34ee",x"b9fc",x"4001",x"3752",x"b24e",x"3bb3",x"31e9",x"364f",x"34df"),
(x"b9f5",x"3ff5",x"377c",x"b068",x"a815",x"3beb",x"35f4",x"1e8d",x"ba00",x"3ffd",x"377a",x"b068",x"a815",x"3beb",x"35ed",x"20c2",x"b9f6",x"4000",x"377d",x"b068",x"a815",x"3beb",x"35f4",x"2148"),
(x"b9f6",x"4000",x"377d",x"bbe8",x"aaec",x"b08c",x"35fb",x"3073",x"b9f7",x"3ffd",x"3794",x"bbe8",x"aaec",x"b08c",x"35fb",x"305f",x"b9f5",x"3ff5",x"377c",x"bbe8",x"aaec",x"b08c",x"35ed",x"3063"),
(x"ba07",x"3ffe",x"3752",x"ba94",x"b7fc",x"345d",x"365a",x"31b1",x"ba00",x"3ffd",x"377a",x"ba72",x"b86b",x"32c9",x"3669",x"31b3",x"b9f5",x"3ff5",x"377c",x"b9d9",x"b836",x"36f1",x"366f",x"3198"),
(x"b9e5",x"3ffc",x"37b2",x"b8ae",x"b826",x"38fc",x"3686",x"31ae",x"b9c9",x"3fdf",x"3787",x"b8c1",x"b811",x"38fb",x"3686",x"3146",x"b9ed",x"3fec",x"376e",x"b8f8",x"b816",x"38c1",x"366f",x"3179"),
(x"b9c9",x"3fdf",x"3787",x"3776",x"b053",x"3afe",x"3632",x"2c6d",x"b9e5",x"3ffc",x"37b2",x"3422",x"b30f",x"3b86",x"3632",x"2b49",x"b9db",x"3ffd",x"37ae",x"3776",x"b053",x"3afe",x"362b",x"2b5e"),
(x"b9e5",x"3ffc",x"37b2",x"b48b",x"3a04",x"38c2",x"362a",x"34ed",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5",x"b9db",x"3ffd",x"37ae",x"335d",x"39d9",x"3923",x"3626",x"34e7"),
(x"b9c9",x"3fdf",x"3787",x"3776",x"b053",x"3afe",x"3632",x"2c6d",x"b9db",x"3ffd",x"37ae",x"3776",x"b053",x"3afe",x"362b",x"2b5e",x"b9d2",x"3ffe",x"379f",x"38fe",x"ab38",x"3a3b",x"3623",x"2b7a"),
(x"b9c5",x"4000",x"3780",x"2cbf",x"3bc6",x"3329",x"3626",x"34ce",x"b9d2",x"3ffe",x"379f",x"354f",x"39c9",x"38d8",x"3624",x"34df",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"b9fc",x"4001",x"3752",x"b24e",x"3bb3",x"31e9",x"364f",x"34df",x"b9de",x"4001",x"3752",x"9d87",x"3bf5",x"2e87",x"3640",x"34ce",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"b9fc",x"4001",x"3752",x"b24e",x"3bb3",x"31e9",x"364f",x"34df",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5",x"b9f6",x"4000",x"377d",x"b5fa",x"3ae9",x"3563",x"3641",x"34e8"),
(x"b9b2",x"3fff",x"37ca",x"a393",x"3b79",x"35b2",x"362a",x"2f26",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e",x"b9a9",x"3ffc",x"37d9",x"3146",x"3a67",x"389c",x"3623",x"2f40"),
(x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b9b2",x"3fff",x"37ca",x"a393",x"3b79",x"35b2",x"362a",x"2f26",x"b9cc",x"3ffd",x"37d0",x"b1ec",x"3b16",x"36cd",x"363e",x"2f34"),
(x"b9b2",x"3ff6",x"37ca",x"3950",x"a0ea",x"39fa",x"35fe",x"1e8d",x"b9bb",x"3ffd",x"37d9",x"3950",x"a0ea",x"39fa",x"35f6",x"208e",x"b9b2",x"3fff",x"37ca",x"3950",x"a0ea",x"39fa",x"35fe",x"210b"),
(x"b9b2",x"3fff",x"37ca",x"b93c",x"95bc",x"3a0c",x"35e8",x"2d07",x"b9a9",x"3ffc",x"37d9",x"b93c",x"95bc",x"3a0c",x"35df",x"2d1a",x"b9b2",x"3ff6",x"37ca",x"b93c",x"95bc",x"3a0c",x"35e8",x"2d3f"),
(x"b9cc",x"3ffd",x"37d0",x"b33b",x"b811",x"3aa5",x"367e",x"322f",x"b9bb",x"3ffd",x"37d9",x"b325",x"b878",x"3a63",x"3671",x"322e",x"b9b2",x"3ff6",x"37ca",x"1e0a",x"b823",x"3ad8",x"366b",x"3246"),
(x"b994",x"3ffc",x"37cd",x"31e7",x"b81a",x"3ab5",x"3654",x"3237",x"b996",x"3fe3",x"3791",x"3252",x"b816",x"3ab1",x"3657",x"328b",x"b9b3",x"3fe8",x"37ad",x"a3bb",x"b81b",x"3add",x"366c",x"3272"),
(x"b996",x"3fe3",x"3791",x"3ae1",x"b415",x"370f",x"35b4",x"2fb8",x"b994",x"3ffc",x"37cd",x"3af6",x"b475",x"367c",x"35a3",x"3029",x"b98f",x"3ffc",x"37ba",x"3b3a",x"b41e",x"357a",x"35ab",x"3028"),
(x"b994",x"3ffc",x"37cd",x"358a",x"3a1b",x"385c",x"3613",x"2f2b",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e",x"b98f",x"3ffc",x"37ba",x"3925",x"39b7",x"3465",x"360f",x"2f0f"),
(x"b996",x"3fe3",x"3791",x"3ae1",x"b415",x"370f",x"35b4",x"2fb8",x"b98f",x"3ffc",x"37ba",x"3b3a",x"b41e",x"357a",x"35ab",x"3028",x"b98a",x"3ffc",x"379b",x"3ad4",x"b3bd",x"3760",x"35b7",x"3027"),
(x"b997",x"3fff",x"3781",x"31af",x"3bdf",x"1c18",x"3615",x"2eb7",x"b98a",x"3ffc",x"379b",x"3825",x"3acf",x"2d30",x"360b",x"2ee1",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b9c5",x"4000",x"3780",x"96f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e",x"b9b2",x"3fff",x"37ca",x"a393",x"3b79",x"35b2",x"362a",x"2f26"),
(x"b9c5",x"4000",x"3780",x"96f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b9d2",x"3ffe",x"379f",x"b94b",x"39eb",x"af9c",x"3644",x"2eeb"),
(x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b9cc",x"3ffd",x"37d0",x"b1ec",x"3b16",x"36cd",x"363e",x"2f34",x"b9d4",x"3ffd",x"37ba",x"b92f",x"39d8",x"32de",x"3644",x"2f14"),
(x"b9d4",x"3ffd",x"37ba",x"bb76",x"b463",x"3373",x"35ff",x"3145",x"b9cc",x"3ffd",x"37d0",x"b9f1",x"b5fe",x"3870",x"3609",x"314d",x"b9c9",x"3fdf",x"3787",x"bb76",x"b463",x"3373",x"3609",x"30e6"),
(x"b9c9",x"3fdf",x"3787",x"bb76",x"b463",x"3373",x"3609",x"30e6",x"b9d2",x"3ffe",x"379f",x"bbda",x"afe2",x"b0aa",x"35f6",x"313b",x"b9d4",x"3ffd",x"37ba",x"bb76",x"b463",x"3373",x"35ff",x"3145"),
(x"b98a",x"3ffc",x"379b",x"3ad4",x"b3bd",x"3760",x"35b7",x"3027",x"b992",x"3fe3",x"378f",x"345c",x"b0de",x"3b99",x"35b7",x"2fb9",x"b996",x"3fe3",x"3791",x"3ae1",x"b415",x"370f",x"35b4",x"2fb8"),
(x"b992",x"3fe3",x"378f",x"a8e0",x"aefd",x"3bf2",x"369d",x"30c9",x"b98a",x"3ffc",x"379b",x"b66b",x"ac20",x"3b4f",x"369d",x"307f",x"b990",x"3fdf",x"378e",x"3496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"b975",x"3ffc",x"37af",x"35ad",x"b6ed",x"3aa0",x"368c",x"3079",x"b96d",x"3fec",x"376e",x"3931",x"b7c9",x"38ad",x"367c",x"30b4",x"b990",x"3fdf",x"378e",x"3496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"b964",x"3ff5",x"377b",x"39d9",x"b840",x"36d9",x"3678",x"3096",x"b975",x"3ffc",x"37af",x"35ad",x"b6ed",x"3aa0",x"368c",x"3079",x"b962",x"3ffb",x"378b",x"3815",x"b8b5",x"3904",x"3679",x"3081"),
(x"b964",x"3ff5",x"377b",x"39d9",x"b840",x"36d9",x"3678",x"3096",x"b95a",x"3ffd",x"3775",x"3a73",x"b85c",x"3351",x"366e",x"3082",x"b953",x"3ffe",x"3752",x"3a86",x"b81f",x"3433",x"3660",x"3089"),
(x"b964",x"3ffd",x"3797",x"3b81",x"34c0",x"31b9",x"35cc",x"214e",x"b964",x"4000",x"3780",x"3bd2",x"3047",x"b134",x"35cc",x"200a",x"b962",x"3ffb",x"378b",x"3bd2",x"3047",x"b133",x"35c7",x"210d"),
(x"b964",x"3ff5",x"377b",x"3612",x"af46",x"3b58",x"35d6",x"214e",x"b964",x"4000",x"3780",x"366b",x"ad14",x"3b4c",x"35d6",x"1e80",x"b95a",x"3ffd",x"3775",x"366c",x"ad14",x"3b4c",x"35cd",x"1ffb"),
(x"b975",x"3ffc",x"37af",x"1fae",x"3964",x"39e8",x"35ca",x"32fc",x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec",x"b964",x"3ffd",x"3797",x"3553",x"3a2a",x"3859",x"35bc",x"3307"),
(x"b992",x"4001",x"3777",x"b179",x"3b46",x"3611",x"35c7",x"32bf",x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec",x"b98a",x"3ffc",x"379b",x"b5ee",x"392f",x"3951",x"35d0",x"32dc"),
(x"b992",x"4001",x"3777",x"b179",x"3b46",x"3611",x"35c7",x"32bf",x"b98a",x"3ffc",x"379b",x"b5ee",x"392f",x"3951",x"35d0",x"32dc",x"b997",x"3fff",x"3781",x"b106",x"3a66",x"38a1",x"35cd",x"32bf"),
(x"b992",x"4001",x"3777",x"b179",x"3b46",x"3611",x"35c7",x"32bf",x"b987",x"4001",x"375e",x"28c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec"),
(x"b95c",x"3fff",x"3777",x"391d",x"39e9",x"32d4",x"35ae",x"32ff",x"b95c",x"4001",x"3752",x"3411",x"3b93",x"3249",x"35a3",x"32ec",x"b95a",x"3ffd",x"3775",x"39ba",x"391c",x"347b",x"35ab",x"3307"),
(x"b987",x"4001",x"375e",x"28c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"b982",x"4001",x"3752",x"24f0",x"3bea",x"309d",x"35b4",x"32bf",x"b964",x"4000",x"3780",x"2de0",x"3bd5",x"31bf",x"35b4",x"32f9"),
(x"b95c",x"3fff",x"3777",x"391d",x"39e9",x"32d4",x"35ae",x"32ff",x"b964",x"4000",x"3780",x"2de0",x"3bd5",x"31bf",x"35b4",x"32f9",x"b95c",x"4001",x"3752",x"3411",x"3b93",x"3249",x"35a3",x"32ec"),
(x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5",x"b9e5",x"3ffc",x"37b2",x"b48b",x"3a04",x"38c2",x"362a",x"34ed",x"b9f7",x"3ffd",x"3794",x"b663",x"3a38",x"37c6",x"363b",x"34f0"),
(x"ba00",x"3ffd",x"377a",x"b865",x"3a42",x"34ab",x"3647",x"34ee",x"ba07",x"3ffe",x"3752",x"b892",x"3a2a",x"347f",x"3655",x"34e7",x"b9fc",x"4001",x"3752",x"b24e",x"3bb3",x"31e9",x"364f",x"34df"),
(x"b9f5",x"3ff5",x"377c",x"b9d9",x"b836",x"36f1",x"366f",x"3198",x"b9f4",x"3fee",x"3752",x"ba96",x"b7a7",x"34e2",x"3663",x"317c",x"ba07",x"3ffe",x"3752",x"ba94",x"b7fc",x"345d",x"365a",x"31b1"),
(x"b9f5",x"3ff5",x"377c",x"b9d9",x"b836",x"36f1",x"366f",x"3198",x"b9ed",x"3fec",x"376e",x"b8f8",x"b816",x"38c1",x"366f",x"3179",x"b9f4",x"3fee",x"3752",x"ba96",x"b7a7",x"34e2",x"3663",x"317c"),
(x"b9e5",x"3ffc",x"37b2",x"b8ae",x"b826",x"38fc",x"3686",x"31ae",x"b9f5",x"3ff5",x"377c",x"b9d9",x"b836",x"36f1",x"366f",x"3198",x"b9f7",x"3ffd",x"3794",x"b839",x"b89f",x"38fa",x"3675",x"31b3"),
(x"b9e5",x"3ffc",x"37b2",x"b8ae",x"b826",x"38fc",x"3686",x"31ae",x"b9ed",x"3fec",x"376e",x"b8f8",x"b816",x"38c1",x"366f",x"3179",x"b9f5",x"3ff5",x"377c",x"b9d9",x"b836",x"36f1",x"366f",x"3198"),
(x"b9d2",x"3ffe",x"379f",x"354f",x"39c9",x"38d8",x"3624",x"34df",x"b9db",x"3ffd",x"37ae",x"335d",x"39d9",x"3923",x"3626",x"34e7",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"b9de",x"4001",x"3752",x"9d87",x"3bf5",x"2e87",x"3640",x"34ce",x"b9c5",x"4000",x"3780",x"2cbf",x"3bc6",x"3329",x"3626",x"34ce",x"b9e1",x"4000",x"37a1",x"ab52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e",x"b994",x"3ffc",x"37cd",x"358a",x"3a1b",x"385c",x"3613",x"2f2b",x"b9a9",x"3ffc",x"37d9",x"3146",x"3a67",x"389c",x"3623",x"2f40"),
(x"b9b2",x"3fff",x"37ca",x"a393",x"3b79",x"35b2",x"362a",x"2f26",x"b9bb",x"3ffd",x"37d9",x"ae09",x"3b05",x"3784",x"3631",x"2f41",x"b9cc",x"3ffd",x"37d0",x"b1ec",x"3b16",x"36cd",x"363e",x"2f34"),
(x"b9b3",x"3fe8",x"37ad",x"a3bb",x"b81b",x"3add",x"366c",x"3272",x"b9c9",x"3fdf",x"3787",x"b409",x"b819",x"3a90",x"367e",x"3296",x"b9cc",x"3ffd",x"37d0",x"b33b",x"b811",x"3aa5",x"367e",x"322f"),
(x"b9cc",x"3ffd",x"37d0",x"b33b",x"b811",x"3aa5",x"367e",x"322f",x"b9b2",x"3ff6",x"37ca",x"1e0a",x"b823",x"3ad8",x"366b",x"3246",x"b9b3",x"3fe8",x"37ad",x"a3bb",x"b81b",x"3add",x"366c",x"3272"),
(x"b994",x"3ffc",x"37cd",x"31e7",x"b81a",x"3ab5",x"3654",x"3237",x"b9b2",x"3ff6",x"37ca",x"1e0a",x"b823",x"3ad8",x"366b",x"3246",x"b9a9",x"3ffc",x"37d9",x"324d",x"b8ad",x"3a4b",x"3664",x"3230"),
(x"b994",x"3ffc",x"37cd",x"31e7",x"b81a",x"3ab5",x"3654",x"3237",x"b9b3",x"3fe8",x"37ad",x"a3bb",x"b81b",x"3add",x"366c",x"3272",x"b9b2",x"3ff6",x"37ca",x"1e0a",x"b823",x"3ad8",x"366b",x"3246"),
(x"b98a",x"3ffc",x"379b",x"3825",x"3acf",x"2d30",x"360b",x"2ee1",x"b98f",x"3ffc",x"37ba",x"3925",x"39b7",x"3465",x"360f",x"2f0f",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"b9c5",x"4000",x"3780",x"96f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"b997",x"3fff",x"3781",x"31af",x"3bdf",x"1c18",x"3615",x"2eb7",x"b998",x"4000",x"37bc",x"30a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"b9ce",x"4000",x"37b1",x"af93",x"3bda",x"30c0",x"363e",x"2f02",x"b9d4",x"3ffd",x"37ba",x"b92f",x"39d8",x"32de",x"3644",x"2f14",x"b9d2",x"3ffe",x"379f",x"b94b",x"39eb",x"af9c",x"3644",x"2eeb"),
(x"b98a",x"3ffc",x"379b",x"b66b",x"ac20",x"3b4f",x"369d",x"307f",x"b975",x"3ffc",x"37af",x"35ad",x"b6ed",x"3aa0",x"368c",x"3079",x"b990",x"3fdf",x"378e",x"3496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"b96d",x"3fec",x"376e",x"3931",x"b7c9",x"38ad",x"367c",x"30b4",x"b98a",x"3fdf",x"377f",x"392b",x"b842",x"385f",x"3694",x"30d7",x"b990",x"3fdf",x"378e",x"3496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"b962",x"3ffb",x"378b",x"3815",x"b8b5",x"3904",x"3679",x"3081",x"b975",x"3ffc",x"37af",x"35ad",x"b6ed",x"3aa0",x"368c",x"3079",x"b964",x"3ffd",x"3797",x"3810",x"b8bd",x"3900",x"367c",x"3079"),
(x"b964",x"3ff5",x"377b",x"39d9",x"b840",x"36d9",x"3678",x"3096",x"b96d",x"3fec",x"376e",x"3931",x"b7c9",x"38ad",x"367c",x"30b4",x"b975",x"3ffc",x"37af",x"35ad",x"b6ed",x"3aa0",x"368c",x"3079"),
(x"b964",x"3ff5",x"377b",x"39d9",x"b840",x"36d9",x"3678",x"3096",x"b967",x"3fee",x"3752",x"3a94",x"b7fd",x"3459",x"3671",x"30b8",x"b96d",x"3fec",x"376e",x"3931",x"b7c9",x"38ad",x"367c",x"30b4"),
(x"b964",x"3ff5",x"377b",x"39d9",x"b840",x"36d9",x"3678",x"3096",x"b953",x"3ffe",x"3752",x"3a86",x"b81f",x"3433",x"3660",x"3089",x"b967",x"3fee",x"3752",x"3a94",x"b7fd",x"3459",x"3671",x"30b8"),
(x"b964",x"4000",x"3780",x"3bd2",x"3047",x"b134",x"35cc",x"200a",x"b964",x"3ff5",x"377b",x"3b82",x"286d",x"b57a",x"35bc",x"20d5",x"b962",x"3ffb",x"378b",x"3bd2",x"3047",x"b133",x"35c7",x"210d"),
(x"b964",x"4000",x"3780",x"366b",x"ad14",x"3b4c",x"35d6",x"1e80",x"b95c",x"3fff",x"3777",x"3827",x"3037",x"3ac1",x"35cf",x"1efe",x"b95a",x"3ffd",x"3775",x"366c",x"ad14",x"3b4c",x"35cd",x"1ffb"),
(x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec",x"b964",x"4000",x"3780",x"2de0",x"3bd5",x"31bf",x"35b4",x"32f9",x"b964",x"3ffd",x"3797",x"3553",x"3a2a",x"3859",x"35bc",x"3307"),
(x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec",x"b975",x"3ffc",x"37af",x"1fae",x"3964",x"39e8",x"35ca",x"32fc",x"b98a",x"3ffc",x"379b",x"b5ee",x"392f",x"3951",x"35d0",x"32dc"),
(x"b987",x"4001",x"375e",x"28c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"b964",x"4000",x"3780",x"2de0",x"3bd5",x"31bf",x"35b4",x"32f9",x"b97a",x"4000",x"37a0",x"10ea",x"3b79",x"35b5",x"35c6",x"32ec"),
(x"b95c",x"4001",x"3752",x"3411",x"3b93",x"3249",x"35a3",x"32ec",x"b953",x"3ffe",x"3752",x"38cb",x"39c5",x"358d",x"359e",x"32fc",x"b95a",x"3ffd",x"3775",x"39ba",x"391c",x"347b",x"35ab",x"3307"),
(x"b982",x"4001",x"3752",x"24f0",x"3bea",x"309d",x"35b4",x"32bf",x"b95c",x"4001",x"3752",x"3411",x"3b93",x"3249",x"35a3",x"32ec",x"b964",x"4000",x"3780",x"2de0",x"3bd5",x"31bf",x"35b4",x"32f9"),
(x"b9df",x"1ef5",x"376e",x"bb33",x"0000",x"b6f8",x"3276",x"21dd",x"b9df",x"3ce9",x"376e",x"bbb7",x"0000",x"b435",x"3277",x"3554",x"b9e1",x"22af",x"3794",x"bbff",x"0000",x"a460",x"32a3",x"2363"),
(x"b9e1",x"22af",x"3794",x"bbff",x"0000",x"a460",x"32a3",x"2363",x"b9e1",x"3ce9",x"3794",x"bbfe",x"0000",x"27ef",x"32a6",x"3554",x"b9de",x"2680",x"37e5",x"bbe2",x"0000",x"315e",x"32d0",x"2479"),
(x"b9de",x"2680",x"37e5",x"bbe2",x"0000",x"315e",x"32d0",x"2479",x"b9de",x"3ce9",x"37e5",x"bb99",x"0000",x"34ff",x"32d4",x"3554",x"b9d2",x"2805",x"3807",x"ba4b",x"8000",x"38f0",x"3301",x"253c"),
(x"b9d2",x"2805",x"3807",x"ba4b",x"8000",x"38f0",x"3301",x"253c",x"b9d2",x"3ce9",x"3807",x"b970",x"0000",x"39dd",x"3302",x"3554",x"b9c1",x"2869",x"3813",x"b68f",x"0000",x"3b4b",x"332f",x"25a6"),
(x"b9c1",x"2869",x"3813",x"b68f",x"0000",x"3b4b",x"332f",x"25a6",x"b9c1",x"3ce9",x"3813",x"b4a7",x"0000",x"3ba7",x"3330",x"3555",x"b9a7",x"28ad",x"3818",x"2495",x"0000",x"3bff",x"335d",x"25cb"),
(x"b9a7",x"3ce9",x"3818",x"2495",x"0000",x"3bff",x"335e",x"3555",x"b98f",x"3ce9",x"3812",x"361b",x"0000",x"3b64",x"338c",x"3555",x"b9a7",x"28ad",x"3818",x"2495",x"0000",x"3bff",x"335d",x"25cb"),
(x"b98f",x"3ce9",x"3812",x"361b",x"0000",x"3b64",x"338c",x"3555",x"b97c",x"3ce9",x"3802",x"39c4",x"0000",x"398b",x"33ba",x"3554",x"b98f",x"2870",x"3812",x"381e",x"0000",x"3adb",x"338b",x"2594"),
(x"b97c",x"3ce9",x"3802",x"39c4",x"0000",x"398b",x"33ba",x"3554",x"b975",x"3ce9",x"37e4",x"3b9c",x"0000",x"34ef",x"33e9",x"3554",x"b97c",x"27a4",x"3802",x"3a87",x"8000",x"389f",x"33b9",x"2503"),
(x"b975",x"3ce9",x"37e4",x"3b9c",x"0000",x"34ef",x"33e9",x"3554",x"b972",x"3ce9",x"37ba",x"3bfc",x"0000",x"2be2",x"340b",x"3554",x"b975",x"2661",x"37e4",x"3bd4",x"8000",x"328e",x"33e7",x"2438"),
(x"b972",x"3ce9",x"37ba",x"3bfc",x"0000",x"2be2",x"340b",x"3554",x"b972",x"3ce9",x"3775",x"3bfd",x"0000",x"aac8",x"3423",x"3554",x"b972",x"24c7",x"37ba",x"3bff",x"0000",x"26a1",x"340b",x"22bc"),
(x"b972",x"3ce9",x"3775",x"3bfd",x"0000",x"aac8",x"3423",x"3554",x"b976",x"3ce9",x"3764",x"3aa9",x"8000",x"b86d",x"343b",x"3554",x"b972",x"2065",x"3775",x"3be7",x"0000",x"b0fd",x"3423",x"2104"),
(x"b976",x"3ce9",x"3764",x"3aa9",x"8000",x"b86d",x"343b",x"3554",x"b97f",x"3ce9",x"3752",x"398d",x"8000",x"b9c2",x"3453",x"3554",x"b976",x"1d1b",x"3764",x"3a17",x"0000",x"b92f",x"343b",x"1d79"),
(x"b9d5",x"1a08",x"3752",x"ba65",x"8000",x"b8cd",x"3245",x"207d",x"b9d5",x"3ce9",x"3752",x"ba65",x"8000",x"b8cd",x"3248",x"3554",x"b9df",x"1ef5",x"376e",x"bb33",x"0000",x"b6f8",x"3276",x"21dd"),
(x"b98f",x"2870",x"3812",x"99bc",x"bac2",x"3846",x"35ed",x"3482",x"b97c",x"27a4",x"3802",x"2352",x"bab1",x"3860",x"35fb",x"3474",x"b9a7",x"28ad",x"3818",x"2495",x"ba9b",x"3881",x"35db",x"3487"),
(x"b9df",x"1ef5",x"376e",x"1c81",x"baa0",x"387b",x"35af",x"3433",x"b976",x"1d1b",x"3764",x"8a8d",x"baca",x"383a",x"35fd",x"342e",x"b9d5",x"1a08",x"3752",x"9a24",x"bb18",x"3761",x"35b6",x"3427"),
(x"b976",x"1d1b",x"3764",x"8a8d",x"baca",x"383a",x"35fd",x"342e",x"b9df",x"1ef5",x"376e",x"1c81",x"baa0",x"387b",x"35af",x"3433",x"b972",x"2065",x"3775",x"1da1",x"bab0",x"3862",x"3600",x"3436"),
(x"b972",x"2065",x"3775",x"1da1",x"bab0",x"3862",x"3600",x"3436",x"b9e1",x"22af",x"3794",x"1953",x"bac8",x"383d",x"35ae",x"3444",x"b972",x"24c7",x"37ba",x"928d",x"bad3",x"382c",x"3601",x"3454"),
(x"b972",x"24c7",x"37ba",x"928d",x"bad3",x"382c",x"3601",x"3454",x"b9de",x"2680",x"37e5",x"9af6",x"bad3",x"382b",x"35b1",x"3467",x"b975",x"2661",x"37e4",x"9b5f",x"badf",x"3817",x"3600",x"3466"),
(x"b97c",x"27a4",x"3802",x"2352",x"bab1",x"3860",x"35fb",x"3474",x"b975",x"2661",x"37e4",x"9b5f",x"badf",x"3817",x"3600",x"3466",x"b9c1",x"2869",x"3813",x"1e3f",x"bacb",x"3838",x"35c8",x"3482"),
(x"b9df",x"3ce9",x"376e",x"bbb7",x"0000",x"b435",x"3277",x"3554",x"b9e1",x"3ce9",x"3794",x"bbfe",x"0000",x"27ef",x"32a6",x"3554",x"b9e1",x"22af",x"3794",x"bbff",x"0000",x"a460",x"32a3",x"2363"),
(x"b9e1",x"3ce9",x"3794",x"bbfe",x"0000",x"27ef",x"32a6",x"3554",x"b9de",x"3ce9",x"37e5",x"bb99",x"0000",x"34ff",x"32d4",x"3554",x"b9de",x"2680",x"37e5",x"bbe2",x"0000",x"315e",x"32d0",x"2479"),
(x"b9de",x"3ce9",x"37e5",x"bb99",x"0000",x"34ff",x"32d4",x"3554",x"b9d2",x"3ce9",x"3807",x"b970",x"0000",x"39dd",x"3302",x"3554",x"b9d2",x"2805",x"3807",x"ba4b",x"8000",x"38f0",x"3301",x"253c"),
(x"b9d2",x"3ce9",x"3807",x"b970",x"0000",x"39dd",x"3302",x"3554",x"b9c1",x"3ce9",x"3813",x"b4a7",x"0000",x"3ba7",x"3330",x"3555",x"b9c1",x"2869",x"3813",x"b68f",x"0000",x"3b4b",x"332f",x"25a6"),
(x"b9c1",x"3ce9",x"3813",x"b4a7",x"0000",x"3ba7",x"3330",x"3555",x"b9a7",x"3ce9",x"3818",x"2495",x"0000",x"3bff",x"335e",x"3555",x"b9a7",x"28ad",x"3818",x"2495",x"0000",x"3bff",x"335d",x"25cb"),
(x"b98f",x"3ce9",x"3812",x"361b",x"0000",x"3b64",x"338c",x"3555",x"b98f",x"2870",x"3812",x"381e",x"0000",x"3adb",x"338b",x"2594",x"b9a7",x"28ad",x"3818",x"2495",x"0000",x"3bff",x"335d",x"25cb"),
(x"b97c",x"3ce9",x"3802",x"39c4",x"0000",x"398b",x"33ba",x"3554",x"b97c",x"27a4",x"3802",x"3a87",x"8000",x"389f",x"33b9",x"2503",x"b98f",x"2870",x"3812",x"381e",x"0000",x"3adb",x"338b",x"2594"),
(x"b975",x"3ce9",x"37e4",x"3b9c",x"0000",x"34ef",x"33e9",x"3554",x"b975",x"2661",x"37e4",x"3bd4",x"8000",x"328e",x"33e7",x"2438",x"b97c",x"27a4",x"3802",x"3a87",x"8000",x"389f",x"33b9",x"2503"),
(x"b972",x"3ce9",x"37ba",x"3bfc",x"0000",x"2be2",x"340b",x"3554",x"b972",x"24c7",x"37ba",x"3bff",x"0000",x"26a1",x"340b",x"22bc",x"b975",x"2661",x"37e4",x"3bd4",x"8000",x"328e",x"33e7",x"2438"),
(x"b972",x"3ce9",x"3775",x"3bfd",x"0000",x"aac8",x"3423",x"3554",x"b972",x"2065",x"3775",x"3be7",x"0000",x"b0fd",x"3423",x"2104",x"b972",x"24c7",x"37ba",x"3bff",x"0000",x"26a1",x"340b",x"22bc"),
(x"b976",x"3ce9",x"3764",x"3aa9",x"8000",x"b86d",x"343b",x"3554",x"b976",x"1d1b",x"3764",x"3a17",x"0000",x"b92f",x"343b",x"1d79",x"b972",x"2065",x"3775",x"3be7",x"0000",x"b0fd",x"3423",x"2104"),
(x"b97f",x"3ce9",x"3752",x"398d",x"8000",x"b9c2",x"3453",x"3554",x"b97f",x"1a6a",x"3752",x"398d",x"8000",x"b9c2",x"3453",x"1b5d",x"b976",x"1d1b",x"3764",x"3a17",x"0000",x"b92f",x"343b",x"1d79"),
(x"b9d5",x"3ce9",x"3752",x"ba65",x"8000",x"b8cd",x"3248",x"3554",x"b9df",x"3ce9",x"376e",x"bbb7",x"0000",x"b435",x"3277",x"3554",x"b9df",x"1ef5",x"376e",x"bb33",x"0000",x"b6f8",x"3276",x"21dd"),
(x"b97c",x"27a4",x"3802",x"2352",x"bab1",x"3860",x"35fb",x"3474",x"b9c1",x"2869",x"3813",x"1e3f",x"bacb",x"3838",x"35c8",x"3482",x"b9a7",x"28ad",x"3818",x"2495",x"ba9b",x"3881",x"35db",x"3487"),
(x"b976",x"1d1b",x"3764",x"8a8d",x"baca",x"383a",x"35fd",x"342e",x"b97f",x"1a6a",x"3752",x"1c32",x"bb56",x"3661",x"35f6",x"3427",x"b9d5",x"1a08",x"3752",x"9a24",x"bb18",x"3761",x"35b6",x"3427"),
(x"b9df",x"1ef5",x"376e",x"1c81",x"baa0",x"387b",x"35af",x"3433",x"b9e1",x"22af",x"3794",x"1953",x"bac8",x"383d",x"35ae",x"3444",x"b972",x"2065",x"3775",x"1da1",x"bab0",x"3862",x"3600",x"3436"),
(x"b9e1",x"22af",x"3794",x"1953",x"bac8",x"383d",x"35ae",x"3444",x"b9de",x"2680",x"37e5",x"9af6",x"bad3",x"382b",x"35b1",x"3467",x"b972",x"24c7",x"37ba",x"928d",x"bad3",x"382c",x"3601",x"3454"),
(x"b9de",x"2680",x"37e5",x"9af6",x"bad3",x"382b",x"35b1",x"3467",x"b9d2",x"2805",x"3807",x"9e59",x"bae9",x"3806",x"35bb",x"3479",x"b975",x"2661",x"37e4",x"9b5f",x"badf",x"3817",x"3600",x"3466"),
(x"b975",x"2661",x"37e4",x"9b5f",x"badf",x"3817",x"3600",x"3466",x"b9d2",x"2805",x"3807",x"9e59",x"bae9",x"3806",x"35bb",x"3479",x"b9c1",x"2869",x"3813",x"1e3f",x"bacb",x"3838",x"35c8",x"3482"),
(x"ba02",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"3620",x"334e",x"b9f6",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"3639",x"3346",x"ba0d",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"361f",x"3321"),
(x"b9fa",x"3ff0",x"3752",x"b8fd",x"390a",x"3765",x"3622",x"3363",x"b9f0",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"363a",x"3356",x"ba02",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"3620",x"334e"),
(x"b9e5",x"3fec",x"378f",x"28a8",x"3b7d",x"3597",x"363e",x"3365",x"b9f0",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"363a",x"3356",x"b9f2",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"3624",x"336f"),
(x"b9ed",x"3fa7",x"3777",x"bb1d",x"b0f4",x"36e3",x"3643",x"3291",x"b9f6",x"3fa8",x"3752",x"bafd",x"b17a",x"3748",x"3634",x"328d",x"b9fd",x"3fd8",x"3786",x"baf1",x"b050",x"37a7",x"3637",x"331f"),
(x"b9e6",x"3f8a",x"376d",x"baf9",x"af50",x"37a0",x"3649",x"323c",x"b9ee",x"3f8b",x"3752",x"bb0e",x"aeb1",x"3757",x"363e",x"323c",x"b9ed",x"3fa7",x"3777",x"bb1d",x"b0f4",x"36e3",x"3643",x"3291"),
(x"b9e5",x"3fec",x"378f",x"28a8",x"3b7d",x"3597",x"363e",x"3365",x"b9f2",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"3624",x"336f",x"b9da",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"3644",x"3373"),
(x"b9d1",x"3fe2",x"378c",x"39d1",x"382c",x"3722",x"364c",x"3387",x"b9da",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"3644",x"3373",x"b9d3",x"3fe5",x"3782",x"39d9",x"3972",x"a970",x"3645",x"3385"),
(x"b9e6",x"3f8a",x"376d",x"afaf",x"abf2",x"3bed",x"35ad",x"319a",x"b9ed",x"3fa7",x"3777",x"2b83",x"ac13",x"3bf8",x"35a9",x"31f0",x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"b9f5",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"35a5",x"327f",x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9fd",x"3fd8",x"3786",x"a82c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"b9f6",x"3fe5",x"378d",x"ae26",x"ac9e",x"3bf1",x"35a6",x"32a5",x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9fd",x"3fd8",x"3786",x"a82c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"b9f0",x"3fea",x"378e",x"ada8",x"257a",x"3bf7",x"35ab",x"32b3",x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9f6",x"3fe5",x"378d",x"ae26",x"ac9e",x"3bf1",x"35a6",x"32a5"),
(x"b9e3",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9e5",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"35b3",x"32b8"),
(x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9e3",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"b9da",x"3fea",x"378e",x"2e3a",x"2687",x"3bf5",x"35bc",x"32b1"),
(x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9d1",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"35c2",x"329a"),
(x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9cc",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"35c6",x"3293",x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274"),
(x"b9cd",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"35c4",x"323e",x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9cc",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"b9cc",x"3fa8",x"3777",x"abc1",x"ab62",x"3bf8",x"35c2",x"31f0",x"b9d5",x"3faa",x"3777",x"ac2f",x"accc",x"3bf5",x"35bc",x"31f5",x"b9cd",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"35c4",x"323e"),
(x"b9cb",x"3f83",x"3770",x"ae76",x"a7e2",x"3bf4",x"35c1",x"3184",x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9cc",x"3fa8",x"3777",x"abc1",x"ab62",x"3bf8",x"35c2",x"31f0"),
(x"b9da",x"3fab",x"3775",x"b235",x"abd2",x"3bd5",x"35b8",x"31f9",x"b9d5",x"3faa",x"3777",x"ac2f",x"accc",x"3bf5",x"35bc",x"31f5",x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c"),
(x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245",x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9da",x"3fab",x"3775",x"b235",x"abd2",x"3bd5",x"35b8",x"31f9"),
(x"b9d9",x"3fd5",x"3782",x"ae8f",x"aed5",x"3be9",x"35bb",x"3274",x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245"),
(x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293"),
(x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9e1",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"35b6",x"32a0"),
(x"b9e3",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9e5",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1",x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9e5",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298",x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d",x"b9f5",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"35a5",x"327f",x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298"),
(x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5",x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"b9da",x"3fab",x"3775",x"b235",x"abd2",x"3bd5",x"35b8",x"31f9",x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d",x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245",x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298",x"b9d9",x"3fd5",x"3782",x"ae8f",x"aed5",x"3be9",x"35bb",x"3274",x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1",x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293",x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298"),
(x"b9e5",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"35b3",x"32a3",x"b9e1",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"35b6",x"32a0",x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"b9c9",x"3fa7",x"378a",x"bbec",x"2581",x"3053",x"35e3",x"3284",x"b9cb",x"3f83",x"3770",x"bbe8",x"9d04",x"30d3",x"35e4",x"32f1",x"b9cb",x"3fa8",x"3783",x"bb1f",x"a907",x"3740",x"35e6",x"3285"),
(x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236",x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236",x"b9cb",x"3fa8",x"3783",x"bb1f",x"a907",x"3740",x"35e6",x"3285"),
(x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203",x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205",x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236"),
(x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5",x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec",x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203"),
(x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3",x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1",x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5"),
(x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc",x"b9c4",x"3fe1",x"37b6",x"ba64",x"b8cb",x"29c5",x"35e0",x"31dc",x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"b9c4",x"3fe1",x"37c1",x"badd",x"b464",x"b6f2",x"35dc",x"31dd",x"b9c4",x"3fe1",x"37b6",x"ba64",x"b8cb",x"29c5",x"35e0",x"31dc",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9c4",x"3fe1",x"37c1",x"badd",x"b464",x"b6f2",x"35dc",x"31dd",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9ca",x"3fc5",x"37c6",x"baf7",x"2fd7",x"b79c",x"35d2",x"322a"),
(x"b9c8",x"3fa9",x"379f",x"bbfa",x"2c56",x"a7a7",x"35dc",x"327e",x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"b9ca",x"3f8a",x"3790",x"bbff",x"25e3",x"1e73",x"35da",x"32db",x"b9c8",x"3fa9",x"379f",x"bbfa",x"2c56",x"a7a7",x"35dc",x"327e",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"b9ca",x"3f88",x"3798",x"bbe2",x"a70a",x"315a",x"35d6",x"32dd",x"b9ca",x"3f8a",x"3790",x"bbff",x"25e3",x"1e73",x"35da",x"32db",x"b9c9",x"3fa8",x"37b2",x"bbe6",x"a832",x"30eb",x"35d4",x"327f"),
(x"b9ca",x"3fc5",x"37c6",x"baf7",x"2fd7",x"b79c",x"35d2",x"322a",x"b9ca",x"3fc3",x"37d1",x"bbf3",x"a804",x"2ec7",x"35cd",x"322c",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"b9ca",x"3fd3",x"37de",x"bbe7",x"9cea",x"30f2",x"35cc",x"31fd",x"b9ca",x"3fc3",x"37d1",x"bbf3",x"a804",x"2ec7",x"35cd",x"322c",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"b9c9",x"3fdf",x"37dc",x"bbdc",x"28a8",x"31d9",x"35d0",x"31db",x"b9ca",x"3fd3",x"37de",x"bbe7",x"9cea",x"30f2",x"35cc",x"31fd",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"b9ca",x"3fe6",x"37cc",x"bbf2",x"2956",x"2ec5",x"35d9",x"31c8",x"b9c9",x"3fdf",x"37dc",x"bbdc",x"28a8",x"31d9",x"35d0",x"31db",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"b9cb",x"3fe8",x"37b8",x"bbfd",x"2581",x"2a45",x"35e1",x"31c5",x"b9ca",x"3fe6",x"37cc",x"bbf2",x"2956",x"2ec5",x"35d9",x"31c8",x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3",x"b9cb",x"3fe7",x"37a7",x"bbff",x"1ec2",x"2532",x"35e8",x"31ca",x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5",x"b9cb",x"3fe0",x"378e",x"bbf9",x"1818",x"2d46",x"35f0",x"31e1",x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"b9cc",x"3fe0",x"378b",x"baff",x"ad07",x"37a5",x"35f2",x"31e1",x"b9cb",x"3fe0",x"378e",x"bbf9",x"1818",x"2d46",x"35f0",x"31e1",x"b9cc",x"3fd4",x"3784",x"bbeb",x"a025",x"3082",x"35f2",x"3204"),
(x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203",x"b9cc",x"3fd4",x"3784",x"bbeb",x"a025",x"3082",x"35f2",x"3204",x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5"),
(x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236",x"b9cd",x"3fc3",x"377f",x"bbd2",x"a2f6",x"32b9",x"35f0",x"3237",x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203"),
(x"b9cd",x"3fc3",x"377f",x"bbd2",x"a2f6",x"32b9",x"35f0",x"3237",x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236",x"b9cc",x"3fa8",x"3777",x"bbc7",x"a659",x"336e",x"35eb",x"3285"),
(x"b9cc",x"3fa8",x"3777",x"bbc7",x"a659",x"336e",x"35eb",x"3285",x"b9cb",x"3fa8",x"3783",x"bb1f",x"a907",x"3740",x"35e6",x"3285",x"b9cb",x"3f83",x"3770",x"bbe8",x"9d04",x"30d3",x"35e4",x"32f1"),
(x"b9cb",x"3f83",x"3770",x"bbe8",x"9d04",x"30d3",x"35e4",x"32f1",x"b9c9",x"3fa7",x"378a",x"bbec",x"2581",x"3053",x"35e3",x"3284",x"b9ca",x"3f8a",x"3790",x"bbff",x"25e3",x"1e73",x"35da",x"32db"),
(x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9c8",x"3fa9",x"379f",x"bbfa",x"2c56",x"a7a7",x"35dc",x"327e",x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236"),
(x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205"),
(x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec"),
(x"b9c4",x"3fe1",x"37c1",x"badd",x"b464",x"b6f2",x"35dc",x"31dd",x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"b9c4",x"3fe1",x"37b6",x"ba64",x"b8cb",x"29c5",x"35e0",x"31dc",x"b9c4",x"3fe1",x"37c1",x"badd",x"b464",x"b6f2",x"35dc",x"31dd",x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"b9ca",x"3f88",x"3798",x"b86c",x"b134",x"3a89",x"35f5",x"3530",x"b9c9",x"3fa8",x"37b2",x"b870",x"b1f2",x"3a7c",x"35f5",x"3500",x"b9ab",x"3f87",x"37c0",x"248e",x"b255",x"3bd7",x"35d8",x"352f"),
(x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b9ca",x"3fc3",x"37d1",x"b885",x"b324",x"3a5a",x"35f4",x"34d4"),
(x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b9ca",x"3fd3",x"37de",x"b89a",x"ad78",x"3a82",x"35f2",x"34bc"),
(x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b9c9",x"3fdf",x"37dc",x"b869",x"323c",x"3a7d",x"35f0",x"34aa"),
(x"b9aa",x"3feb",x"37e2",x"1953",x"3ada",x"3821",x"35d7",x"349e",x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b9ca",x"3fe6",x"37cc",x"b783",x"398b",x"385f",x"35ef",x"349c"),
(x"b9cb",x"3fe8",x"37b8",x"b5d5",x"3b70",x"2a94",x"35f1",x"3494",x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495",x"b9ca",x"3fe6",x"37cc",x"b783",x"398b",x"385f",x"35ef",x"349c"),
(x"b9cb",x"3fe7",x"37a7",x"b572",x"3a96",x"b740",x"35f3",x"348e",x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e",x"b9cb",x"3fe8",x"37b8",x"b5d5",x"3b70",x"2a94",x"35f1",x"3494"),
(x"b9cb",x"3fe0",x"378e",x"b81d",x"395a",x"b849",x"35f9",x"3481",x"b9c2",x"3fe7",x"379c",x"b620",x"3a0a",x"b841",x"35ed",x"3488",x"b9cb",x"3fe7",x"37a7",x"b572",x"3a96",x"b740",x"35f3",x"348e"),
(x"b9c8",x"3fe1",x"378b",x"b994",x"399e",x"b082",x"35f6",x"3480",x"b9c2",x"3fe7",x"379c",x"b620",x"3a0a",x"b841",x"35ed",x"3488",x"b9cb",x"3fe0",x"378e",x"b81d",x"395a",x"b849",x"35f9",x"3481"),
(x"b9cc",x"3fe0",x"378b",x"388b",x"36b7",x"39a9",x"364e",x"338f",x"b9d1",x"3fe2",x"378c",x"39d1",x"382c",x"3722",x"364c",x"3387",x"b9cb",x"3fe1",x"3786",x"388d",x"3867",x"38e2",x"364c",x"3391"),
(x"b9cc",x"3fe0",x"378b",x"b8bf",x"3999",x"3659",x"35fa",x"3480",x"b9cb",x"3fe1",x"3786",x"b81c",x"39f5",x"36cf",x"35f8",x"347e",x"b9cb",x"3fe0",x"378e",x"b81e",x"395a",x"b84a",x"35f9",x"3481"),
(x"b953",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"35ab",x"2e39",x"b949",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"35ab",x"2e93",x"b960",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"35c4",x"2e47"),
(x"b95c",x"3ff0",x"3752",x"38fd",x"390a",x"3765",x"35ad",x"2e10",x"b953",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"35ab",x"2e39",x"b966",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"35c6",x"2e27"),
(x"b95c",x"3ff0",x"3752",x"38fd",x"390a",x"3765",x"35ad",x"2e10",x"b966",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"35c6",x"2e27",x"b964",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"35af",x"2df7"),
(x"b96a",x"3fa6",x"3775",x"3acd",x"b078",x"380f",x"35cf",x"2fb9",x"b959",x"3fd8",x"3786",x"3ad9",x"b071",x"37f4",x"35c2",x"2e97",x"b960",x"3fa8",x"3752",x"3adc",x"b152",x"37c7",x"35c0",x"2fbb"),
(x"b970",x"3f88",x"376d",x"3a64",x"ad63",x"38c3",x"35d7",x"3033",x"b96a",x"3fa6",x"3775",x"3acd",x"b078",x"380f",x"35cf",x"2fb9",x"b965",x"3f8b",x"3752",x"3ab6",x"ad4f",x"384c",x"35c9",x"302f"),
(x"b964",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"35af",x"2df7",x"b971",x"3fec",x"378f",x"a8a8",x"3b7d",x"3597",x"35ca",x"2e09",x"b97c",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"b985",x"3fe2",x"378c",x"b9bb",x"383c",x"3743",x"35d7",x"2dc5",x"b983",x"3fe5",x"3782",x"b9dc",x"3971",x"a62b",x"35d1",x"2dca",x"b97c",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"b970",x"3f88",x"376d",x"303d",x"a8e0",x"3bec",x"3614",x"3130",x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e",x"b96a",x"3fa6",x"3775",x"2b9a",x"acf0",x"3bf6",x"3611",x"30d8"),
(x"b96a",x"3fa6",x"3775",x"2b9a",x"acf0",x"3bf6",x"3611",x"30d8",x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2",x"b959",x"3fd8",x"3786",x"2e54",x"ae94",x"3beb",x"3607",x"3046"),
(x"b960",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"360d",x"3020",x"b959",x"3fd8",x"3786",x"2e54",x"ae94",x"3beb",x"3607",x"3046",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026"),
(x"b966",x"3fea",x"378e",x"2da8",x"257a",x"3bf7",x"3612",x"3012",x"b960",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"360d",x"3020",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"b966",x"3fea",x"378e",x"2da8",x"257a",x"3bf7",x"3612",x"3012",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a",x"b971",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"361b",x"300d"),
(x"b971",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"361b",x"300d",x"b972",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"361b",x"3016",x"b97c",x"3fea",x"378e",x"ae3a",x"2687",x"3bf5",x"3623",x"3014"),
(x"b97c",x"3fea",x"378e",x"ae3a",x"2687",x"3bf5",x"3623",x"3014",x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b985",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051",x"b989",x"3fe0",x"378b",x"af00",x"af3d",x"3be6",x"362d",x"3032",x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f"),
(x"b989",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"362b",x"3087",x"b98a",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"362d",x"3054",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082"),
(x"b989",x"3fa8",x"3777",x"26fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"b989",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"362b",x"3087",x"b981",x"3faa",x"3777",x"2c34",x"acb2",x"3bf5",x"3623",x"30d0"),
(x"b98b",x"3f89",x"3770",x"2987",x"a828",x"3bfc",x"3628",x"312f",x"b989",x"3fa8",x"3777",x"26fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"b981",x"3faa",x"3777",x"2c34",x"acb2",x"3bf5",x"3623",x"30d0",x"b97c",x"3fab",x"3775",x"3227",x"ab9d",x"3bd6",x"361f",x"30cb",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080",x"b97c",x"3fab",x"3775",x"3227",x"ab9d",x"3bd6",x"361f",x"30cb",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082"),
(x"b97d",x"3fd5",x"3782",x"2e8f",x"aed5",x"3be9",x"3623",x"3050",x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080",x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051"),
(x"b97d",x"3fd5",x"3782",x"2e8f",x"aed5",x"3be9",x"3623",x"3050",x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051",x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032",x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f",x"b975",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"361d",x"3025"),
(x"b975",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"361d",x"3025",x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b971",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"361a",x"3022"),
(x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b971",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"361a",x"3022",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026"),
(x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b961",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"360d",x"3046"),
(x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2"),
(x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2",x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e",x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0"),
(x"b97c",x"3fab",x"3775",x"3227",x"ab9d",x"3bd6",x"361f",x"30cb",x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080"),
(x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b97d",x"3fd5",x"3782",x"2e8f",x"aed5",x"3be9",x"3623",x"3050"),
(x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"b971",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"361a",x"3022",x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b975",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"361d",x"3025"),
(x"b98b",x"3f89",x"3770",x"3bf0",x"1d6d",x"2fcb",x"360f",x"3168",x"b98d",x"3fa8",x"378a",x"3be0",x"2467",x"319c",x"360d",x"31c3",x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4"),
(x"b98b",x"3fc2",x"378b",x"3a70",x"a9d2",x"38bb",x"3615",x"3211",x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4",x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b98b",x"3fc2",x"378b",x"3a70",x"a9d2",x"38bb",x"3615",x"3211",x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263",x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b"),
(x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268"),
(x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b",x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b991",x"3fe2",x"37b7",x"3a93",x"b88d",x"2474",x"360a",x"326f"),
(x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b",x"b991",x"3fe2",x"37b7",x"3a93",x"b88d",x"2474",x"360a",x"326f",x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277"),
(x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277",x"b991",x"3fe1",x"37c3",x"3b15",x"b384",x"b669",x"3606",x"326c",x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266",x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b98c",x"3fd3",x"37d2",x"3a75",x"2987",x"b8b5",x"35fc",x"3249"),
(x"b98c",x"3fd3",x"37d2",x"3a75",x"2987",x"b8b5",x"35fc",x"3249",x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e"),
(x"b98c",x"3fa9",x"37a5",x"3bef",x"2703",x"afec",x"3603",x"31c9",x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e",x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9"),
(x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9",x"b98b",x"3f85",x"378d",x"3bff",x"2504",x"1d6d",x"3604",x"3160",x"b98c",x"3fa9",x"37a5",x"3bef",x"2703",x"afec",x"3603",x"31c9"),
(x"b98c",x"3f84",x"3797",x"3be3",x"a752",x"313e",x"3600",x"315e",x"b98c",x"3fa8",x"37b0",x"3bfa",x"a217",x"2ca7",x"35ff",x"31c8",x"b98b",x"3f85",x"378d",x"3bff",x"2504",x"1d6d",x"3604",x"3160"),
(x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e",x"b98c",x"3fa9",x"37a5",x"3bef",x"2703",x"afec",x"3603",x"31c9",x"b98c",x"3fc3",x"37d0",x"3bff",x"a2f6",x"24f7",x"35f8",x"321b"),
(x"b98c",x"3fd3",x"37d2",x"3a75",x"2987",x"b8b5",x"35fc",x"3249",x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e",x"b98c",x"3fd3",x"37dc",x"3bff",x"15bc",x"a673",x"35f8",x"324b"),
(x"b98c",x"3fd3",x"37d2",x"3a75",x"2987",x"b8b5",x"35fc",x"3249",x"b98c",x"3fd3",x"37dc",x"3bff",x"15bc",x"a673",x"35f8",x"324b",x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266",x"b98c",x"3fde",x"37db",x"3bff",x"1953",x"2560",x"35fb",x"326b",x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277"),
(x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277",x"b98c",x"3fe6",x"37cd",x"3bf7",x"29c5",x"2d1b",x"3603",x"327f",x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b"),
(x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b",x"b98b",x"3fe7",x"37a7",x"3bff",x"0cea",x"269a",x"3612",x"327d"),
(x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263",x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b98a",x"3fe0",x"378e",x"3bf8",x"15bc",x"2d81",x"361b",x"3266"),
(x"b98a",x"3fe0",x"378e",x"3bf8",x"15bc",x"2d81",x"361b",x"3266",x"b989",x"3fe0",x"378b",x"3aff",x"ad07",x"37a5",x"361c",x"3266",x"b98a",x"3fd4",x"3784",x"3bea",x"a025",x"3095",x"361c",x"3243"),
(x"b98a",x"3fe0",x"378e",x"3bf8",x"15bc",x"2d81",x"361b",x"3266",x"b98a",x"3fd4",x"3784",x"3bea",x"a025",x"3095",x"361c",x"3243",x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263"),
(x"b98b",x"3fc2",x"378b",x"3a70",x"a9d2",x"38bb",x"3615",x"3211",x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b989",x"3fc3",x"377f",x"3bce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"b989",x"3fa8",x"3777",x"3bc5",x"a793",x"3389",x"3615",x"31c2",x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4",x"b989",x"3fc3",x"377f",x"3bce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4",x"b989",x"3fa8",x"3777",x"3bc5",x"a793",x"3389",x"3615",x"31c2",x"b98b",x"3f89",x"3770",x"3bf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"b98b",x"3f85",x"378d",x"3bff",x"2504",x"1d6d",x"3604",x"3160",x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9",x"b98b",x"3f89",x"3770",x"3bf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"b98d",x"3fa8",x"378a",x"3be0",x"2467",x"319c",x"360d",x"31c3",x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9",x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211",x"b991",x"3fc5",x"37be",x"3beb",x"2c4d",x"b006",x"3601",x"321f",x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242",x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b"),
(x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b",x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268"),
(x"b991",x"3fe1",x"37c3",x"3b15",x"b384",x"b669",x"3606",x"326c",x"b991",x"3fe2",x"37b7",x"3a93",x"b88d",x"2474",x"360a",x"326f",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268"),
(x"b98c",x"3f84",x"3797",x"382d",x"b0b5",x"3ab8",x"35bc",x"3537",x"b9ab",x"3f87",x"37c0",x"248e",x"b255",x"3bd7",x"35d8",x"352f",x"b98c",x"3fa8",x"37b0",x"387f",x"b1e6",x"3a73",x"35ba",x"3500"),
(x"b98c",x"3fa8",x"37b0",x"387f",x"b1e6",x"3a73",x"35ba",x"3500",x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b98c",x"3fc3",x"37d0",x"3896",x"b2c0",x"3a54",x"35bb",x"34d5"),
(x"b98c",x"3fc3",x"37d0",x"3896",x"b2c0",x"3a54",x"35bb",x"34d5",x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b98c",x"3fd3",x"37dc",x"3892",x"ade1",x"3a86",x"35bc",x"34bc"),
(x"b98c",x"3fd3",x"37dc",x"3892",x"ade1",x"3a86",x"35bc",x"34bc",x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b98c",x"3fde",x"37db",x"3885",x"3126",x"3a79",x"35be",x"34ab"),
(x"b98c",x"3fde",x"37db",x"3885",x"3126",x"3a79",x"35be",x"34ab",x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b98c",x"3fe6",x"37cd",x"37e6",x"396d",x"3859",x"35bf",x"349d"),
(x"b98b",x"3fe8",x"37b8",x"361b",x"3b60",x"2bbe",x"35be",x"3495",x"b98c",x"3fe6",x"37cd",x"37e6",x"396d",x"3859",x"35bf",x"349d",x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495"),
(x"b98b",x"3fe7",x"37a7",x"3619",x"3a76",x"b730",x"35bb",x"348f",x"b98b",x"3fe8",x"37b8",x"361b",x"3b60",x"2bbe",x"35be",x"3495",x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e"),
(x"b98a",x"3fe0",x"378e",x"3967",x"383c",x"b81a",x"35b4",x"3483",x"b98b",x"3fe7",x"37a7",x"3619",x"3a76",x"b730",x"35bb",x"348f",x"b993",x"3fe4",x"3789",x"3646",x"3a25",x"b80b",x"35bd",x"3481"),
(x"b993",x"3fe4",x"3789",x"3646",x"3a25",x"b80b",x"35bd",x"3481",x"b98e",x"3fe1",x"378b",x"38bd",x"3a6d",x"2bf2",x"35b7",x"3482",x"b98a",x"3fe0",x"378e",x"3967",x"383c",x"b81a",x"35b4",x"3483"),
(x"b989",x"3fe0",x"378b",x"b8ee",x"37c0",x"38f6",x"35d9",x"2db4",x"b98c",x"3fe1",x"3782",x"b8d3",x"3873",x"3892",x"35d6",x"2daa",x"b985",x"3fe2",x"378c",x"b9bb",x"383c",x"3743",x"35d7",x"2dc5"),
(x"b98a",x"3fe0",x"378e",x"3967",x"383c",x"b81a",x"35b4",x"3483",x"b98e",x"3fe1",x"378b",x"38bd",x"3a6d",x"2bf2",x"35b7",x"3482",x"b989",x"3fe0",x"378b",x"3862",x"3a94",x"30e6",x"35b3",x"3481"),
(x"b970",x"3f88",x"376d",x"3a64",x"ad63",x"38c3",x"35d7",x"3033",x"b965",x"3f8b",x"3752",x"3ab6",x"ad4f",x"384c",x"35c9",x"302f",x"b970",x"3f7e",x"376e",x"3abb",x"aad9",x"384d",x"35d9",x"3052"),
(x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e",x"b970",x"3f88",x"376d",x"303d",x"a8e0",x"3bec",x"3614",x"3130",x"b979",x"3f83",x"3770",x"2e2b",x"280b",x"3bf5",x"361a",x"3141"),
(x"b979",x"3f83",x"3770",x"2e2b",x"280b",x"3bf5",x"361a",x"3141",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e",x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e"),
(x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e",x"b979",x"3f83",x"3770",x"2e2b",x"280b",x"3bf5",x"361a",x"3141",x"b98b",x"3f89",x"3770",x"2987",x"a828",x"3bfc",x"3628",x"312f"),
(x"b9e6",x"3f8a",x"376d",x"baf9",x"af50",x"37a0",x"3649",x"323c",x"b9e4",x"3f7a",x"376e",x"bb00",x"aaa4",x"37b3",x"364e",x"320e",x"b9ee",x"3f8b",x"3752",x"bb0e",x"aeb1",x"3757",x"363e",x"323c"),
(x"b9e4",x"3f7a",x"376e",x"ad21",x"068d",x"3bf9",x"35ad",x"316b",x"b9e6",x"3f8a",x"376d",x"afaf",x"abf2",x"3bed",x"35ad",x"319a",x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"b9e4",x"3f7a",x"376e",x"ad21",x"068d",x"3bf9",x"35ad",x"316b",x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"b9d3",x"3f7f",x"3770",x"a93f",x"1af6",x"3bfe",x"35ba",x"3179"),
(x"b9d3",x"3f7f",x"3770",x"a93f",x"1af6",x"3bfe",x"35ba",x"3179",x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9cb",x"3f83",x"3770",x"ae76",x"a7e2",x"3bf4",x"35c1",x"3184"),
(x"b9f7",x"4032",x"377d",x"b601",x"3ae5",x"3571",x"3629",x"2fc2",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9",x"b9f8",x"4030",x"3794",x"b663",x"3a38",x"37c6",x"3623",x"2fe3"),
(x"b9f7",x"4032",x"377d",x"b601",x"3ae5",x"3571",x"3629",x"2fc2",x"ba01",x"4030",x"377a",x"b864",x"3a40",x"34bc",x"3630",x"2fdb",x"b9fd",x"4033",x"3752",x"b24d",x"3bb2",x"31fb",x"3638",x"2fa0"),
(x"b9f6",x"402c",x"377c",x"b068",x"a815",x"3beb",x"362f",x"3221",x"ba01",x"4030",x"377a",x"b068",x"a815",x"3beb",x"362f",x"3205",x"b9f7",x"4032",x"377d",x"b068",x"a815",x"3beb",x"3626",x"3206"),
(x"b9f7",x"4032",x"377d",x"bbe8",x"aaf0",x"b08c",x"35e0",x"1e8d",x"b9f8",x"4030",x"3794",x"bbe8",x"aaf0",x"b08c",x"35d7",x"1fd1",x"b9f6",x"402c",x"377c",x"bbe8",x"aaf0",x"b08c",x"35e0",x"214e"),
(x"ba08",x"4031",x"3752",x"ba9b",x"b7a9",x"34c2",x"3635",x"3436",x"ba01",x"4030",x"377a",x"ba71",x"b86a",x"32e5",x"3645",x"3436",x"b9f6",x"402c",x"377c",x"b9ed",x"b7fd",x"372e",x"364a",x"3429"),
(x"b9e5",x"4030",x"37b3",x"b89d",x"b810",x"391d",x"3662",x"3434",x"b9c9",x"4021",x"3787",x"b88f",x"b80c",x"392d",x"3662",x"3401",x"b9ed",x"4027",x"376e",x"b8ec",x"b7ef",x"38e6",x"364a",x"3418"),
(x"b9c9",x"4021",x"3787",x"3776",x"b053",x"3afe",x"359c",x"3429",x"b9e5",x"4030",x"37b3",x"3422",x"b30f",x"3b86",x"359c",x"33ee",x"b9dc",x"4030",x"37ae",x"3777",x"b053",x"3afe",x"3595",x"33f3"),
(x"b9e5",x"4030",x"37b3",x"b48b",x"3a03",x"38c2",x"3611",x"2fda",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9",x"b9dc",x"4030",x"37ae",x"335d",x"39d9",x"3923",x"360d",x"2fc2"),
(x"b9c9",x"4021",x"3787",x"3776",x"b053",x"3afe",x"359c",x"3429",x"b9dc",x"4030",x"37ae",x"3777",x"b053",x"3afe",x"3595",x"33f3",x"b9d3",x"4031",x"379f",x"38fe",x"ab38",x"3a3b",x"358d",x"33fa"),
(x"b9c5",x"4033",x"3780",x"2cce",x"3bc5",x"3334",x"360d",x"2f61",x"b9d3",x"4031",x"379f",x"354f",x"39c9",x"38d8",x"360b",x"2fa1",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"b9fd",x"4033",x"3752",x"b24d",x"3bb2",x"31fb",x"3638",x"2fa0",x"b9df",x"4033",x"3752",x"9d04",x"3bf5",x"2e94",x"3627",x"2f61",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"b9fd",x"4033",x"3752",x"b24d",x"3bb2",x"31fb",x"3638",x"2fa0",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9",x"b9f7",x"4032",x"377d",x"b601",x"3ae5",x"3571",x"3629",x"2fc2"),
(x"b9b2",x"4031",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"3355",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349",x"b9a9",x"4030",x"37da",x"3146",x"3a67",x"389c",x"3659",x"3362"),
(x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b9b2",x"4031",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"3355",x"b9cc",x"4030",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"335c"),
(x"b9b2",x"402d",x"37cb",x"3950",x"a0dd",x"39fa",x"35e9",x"2d02",x"b9bb",x"4030",x"37da",x"3950",x"a0dd",x"39fa",x"35e9",x"2ccc",x"b9b2",x"4031",x"37cb",x"3950",x"a0dd",x"39fa",x"35df",x"2cd5"),
(x"b9b2",x"4031",x"37cb",x"b93c",x"95bc",x"3a0c",x"35ec",x"2cc6",x"b9a9",x"4030",x"37da",x"b93c",x"95bc",x"3a0c",x"35ec",x"2c9f",x"b9b2",x"402d",x"37cb",x"b93c",x"95bc",x"3a0c",x"35df",x"2cab"),
(x"b9cc",x"4030",x"37d1",x"b33b",x"b811",x"3aa5",x"3689",x"30d9",x"b9bb",x"4030",x"37da",x"b325",x"b878",x"3a63",x"367b",x"30d7",x"b9b2",x"402d",x"37cb",x"1e0a",x"b823",x"3ad8",x"3676",x"30ef"),
(x"b994",x"4030",x"37cd",x"31e7",x"b81a",x"3ab5",x"365e",x"30e1",x"b996",x"4023",x"3791",x"3252",x"b816",x"3ab1",x"3661",x"3135",x"b9b3",x"4026",x"37ad",x"a3bb",x"b81b",x"3add",x"3677",x"311b"),
(x"b996",x"4023",x"3791",x"3ad4",x"b414",x"3743",x"35b5",x"3046",x"b994",x"4030",x"37cd",x"3af6",x"b475",x"367c",x"35a4",x"3094",x"b98f",x"4030",x"37ba",x"3b3a",x"b41e",x"357a",x"35ac",x"3093"),
(x"b994",x"4030",x"37cd",x"358a",x"3a1b",x"385c",x"3649",x"3358",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349",x"b98f",x"4030",x"37ba",x"3926",x"39b7",x"3465",x"3645",x"334a"),
(x"b996",x"4023",x"3791",x"3ad4",x"b414",x"3743",x"35b5",x"3046",x"b98f",x"4030",x"37ba",x"3b3a",x"b41e",x"357a",x"35ac",x"3093",x"b98a",x"4030",x"379b",x"3abf",x"b3b7",x"37ae",x"35b9",x"3091"),
(x"b997",x"4032",x"3781",x"31af",x"3bdf",x"1c18",x"364b",x"331d",x"b98a",x"4030",x"379b",x"3825",x"3acf",x"2d30",x"3640",x"3332",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b9c5",x"4033",x"3780",x"96f6",x"3bfe",x"27c1",x"366e",x"331d",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349",x"b9b2",x"4031",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"3355"),
(x"b9c5",x"4033",x"3780",x"96f6",x"3bfe",x"27c1",x"366e",x"331d",x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b9d3",x"4031",x"379f",x"b94c",x"39eb",x"af9a",x"367a",x"3337"),
(x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b9cc",x"4030",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"335c",x"b9d5",x"4030",x"37ba",x"b92f",x"39d8",x"32de",x"367a",x"334c"),
(x"b9d5",x"4030",x"37ba",x"bb76",x"b463",x"3373",x"3640",x"2ea4",x"b9cc",x"4030",x"37d1",x"b9f1",x"b5fe",x"3870",x"3649",x"2eb4",x"b9c9",x"4021",x"3787",x"bb76",x"b463",x"3373",x"3649",x"2de4"),
(x"b9c9",x"4021",x"3787",x"bb76",x"b463",x"3373",x"3649",x"2de4",x"b9d3",x"4031",x"379f",x"bbda",x"afe2",x"b0aa",x"3637",x"2e90",x"b9d5",x"4030",x"37ba",x"bb76",x"b463",x"3373",x"3640",x"2ea4"),
(x"b98a",x"4030",x"379b",x"3abf",x"b3b7",x"37ae",x"35b9",x"3091",x"b992",x"4023",x"378f",x"32ea",x"b07f",x"3bba",x"35b9",x"3044",x"b996",x"4023",x"3791",x"3ad4",x"b414",x"3743",x"35b5",x"3046"),
(x"b992",x"4023",x"378f",x"2822",x"af6e",x"3bf1",x"366b",x"352d",x"b98a",x"4030",x"379b",x"b65b",x"ac2a",x"3b52",x"366b",x"3506",x"b990",x"4021",x"378e",x"34a7",x"b630",x"3b00",x"3668",x"3531"),
(x"b975",x"4030",x"37b0",x"35ad",x"b6ed",x"3aa0",x"3659",x"3502",x"b96c",x"4028",x"376e",x"392f",x"b7c9",x"38af",x"3649",x"3520",x"b990",x"4021",x"378e",x"34a7",x"b630",x"3b00",x"3668",x"3531"),
(x"b964",x"402c",x"377a",x"39d4",x"b83f",x"36e9",x"3645",x"3511",x"b975",x"4030",x"37b0",x"35ad",x"b6ed",x"3aa0",x"3659",x"3502",x"b961",x"402f",x"378b",x"3815",x"b8b5",x"3904",x"3646",x"3507"),
(x"b964",x"402c",x"377a",x"39d5",x"b83f",x"36e9",x"3645",x"3511",x"b959",x"4030",x"3775",x"3a72",x"b85a",x"3373",x"363b",x"3507",x"b952",x"4031",x"3752",x"3a84",x"b81e",x"3444",x"362e",x"350b"),
(x"b963",x"4030",x"3797",x"3b81",x"34c0",x"31b9",x"35bb",x"214e",x"b963",x"4032",x"3780",x"3bd2",x"3047",x"b134",x"35bb",x"2006",x"b961",x"402f",x"378b",x"3bd2",x"3047",x"b133",x"35b6",x"210c"),
(x"b964",x"402c",x"377a",x"3612",x"af46",x"3b58",x"362f",x"3202",x"b963",x"4032",x"3780",x"366c",x"ad14",x"3b4c",x"362f",x"31e1",x"b959",x"4030",x"3775",x"366c",x"ad14",x"3b4c",x"3626",x"31ed"),
(x"b975",x"4030",x"37b0",x"1fc8",x"3964",x"39e8",x"360f",x"2e1f",x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f",x"b963",x"4030",x"3797",x"3553",x"3a2a",x"3859",x"361e",x"2e0a"),
(x"b991",x"4033",x"3777",x"b179",x"3b46",x"3611",x"3613",x"2e9a",x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f",x"b98a",x"4030",x"379b",x"b5ee",x"392f",x"3951",x"3609",x"2e60"),
(x"b991",x"4033",x"3777",x"b179",x"3b46",x"3611",x"3613",x"2e9a",x"b98a",x"4030",x"379b",x"b5ee",x"392f",x"3951",x"3609",x"2e60",x"b997",x"4032",x"3781",x"b106",x"3a66",x"38a1",x"360c",x"2e9b"),
(x"b991",x"4033",x"3777",x"b179",x"3b46",x"3611",x"3613",x"2e9a",x"b986",x"4033",x"375d",x"28bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f"),
(x"b95b",x"4032",x"3777",x"391e",x"39e5",x"32f0",x"362c",x"2e19",x"b95b",x"4033",x"3752",x"3410",x"3b92",x"3261",x"3637",x"2e3f",x"b959",x"4030",x"3775",x"39b9",x"391a",x"348e",x"362e",x"2e0a"),
(x"b986",x"4033",x"375d",x"28bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"b981",x"4033",x"3752",x"24c2",x"3be9",x"30b5",x"3625",x"2e99",x"b963",x"4032",x"3780",x"2de3",x"3bd5",x"31ce",x"3625",x"2e26"),
(x"b95b",x"4032",x"3777",x"391e",x"39e5",x"32f0",x"362c",x"2e19",x"b963",x"4032",x"3780",x"2de3",x"3bd5",x"31ce",x"3625",x"2e26",x"b95b",x"4033",x"3752",x"3410",x"3b92",x"3261",x"3637",x"2e3f"),
(x"b9f7",x"405d",x"377d",x"b601",x"3ae5",x"3571",x"365f",x"33e0",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db",x"b9f8",x"405b",x"3794",x"b663",x"3a38",x"37c6",x"3659",x"33f1"),
(x"b9f7",x"405d",x"377d",x"b601",x"3ae5",x"3571",x"365f",x"33e0",x"ba01",x"405b",x"377a",x"b865",x"3a40",x"34bc",x"3665",x"33ed",x"b9fd",x"405e",x"3752",x"b24d",x"3bb2",x"31fb",x"366d",x"33ce"),
(x"b9f6",x"4057",x"377c",x"b068",x"a815",x"3beb",x"362f",x"3241",x"ba01",x"405b",x"377a",x"b068",x"a815",x"3beb",x"362f",x"3224",x"b9f7",x"405d",x"377d",x"b068",x"a815",x"3beb",x"3626",x"3226"),
(x"b9f7",x"405d",x"377d",x"bbe8",x"aaf0",x"b08c",x"35e1",x"20e0",x"b9f8",x"405b",x"3794",x"bbe8",x"aaf0",x"b08c",x"35eb",x"210c",x"b9f6",x"4057",x"377c",x"bbe8",x"aaf0",x"b08c",x"35eb",x"1e8d"),
(x"ba08",x"405c",x"3752",x"ba92",x"b7f9",x"346d",x"3646",x"3307",x"ba01",x"405b",x"377a",x"ba71",x"b86a",x"32e5",x"3655",x"3309",x"b9f6",x"4057",x"377c",x"b9d5",x"b835",x"3700",x"365a",x"32ee"),
(x"b9e5",x"405b",x"37b3",x"b8ae",x"b826",x"38fc",x"3671",x"3303",x"b9c9",x"404c",x"3787",x"b8c1",x"b811",x"38fc",x"3671",x"329b",x"b9ed",x"4053",x"376e",x"b8f6",x"b815",x"38c2",x"365a",x"32ce"),
(x"b9c9",x"404c",x"3787",x"3776",x"b054",x"3afe",x"359b",x"33e2",x"b9e5",x"405b",x"37b3",x"3422",x"b30f",x"3b86",x"359b",x"337d",x"b9dc",x"405b",x"37ae",x"3776",x"b053",x"3afe",x"3594",x"3382"),
(x"b9e5",x"405b",x"37b3",x"b48b",x"3a04",x"38c2",x"3648",x"33ec",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db",x"b9dc",x"405b",x"37ae",x"335d",x"39d9",x"3923",x"3644",x"33e0"),
(x"b9c9",x"404c",x"3787",x"3776",x"b054",x"3afe",x"359b",x"33e2",x"b9dc",x"405b",x"37ae",x"3776",x"b053",x"3afe",x"3594",x"3382",x"b9d3",x"405b",x"379f",x"38fe",x"ab38",x"3a3b",x"358c",x"3389"),
(x"b9c5",x"405d",x"3780",x"2cce",x"3bc5",x"3335",x"3644",x"33ae",x"b9d3",x"405b",x"379f",x"354f",x"39c9",x"38d8",x"3642",x"33cf",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db"),
(x"b9fd",x"405e",x"3752",x"b24d",x"3bb2",x"31fb",x"366d",x"33ce",x"b9df",x"405e",x"3752",x"9d04",x"3bf5",x"2e94",x"365d",x"33ae",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db"),
(x"b9fd",x"405e",x"3752",x"b24d",x"3bb2",x"31fb",x"366d",x"33ce",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db",x"b9f7",x"405d",x"377d",x"b601",x"3ae5",x"3571",x"365f",x"33e0"),
(x"b9b2",x"405c",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"252a",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9",x"b9a9",x"405b",x"37da",x"3146",x"3a67",x"389c",x"3659",x"2595"),
(x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b9b2",x"405c",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"252a",x"b9cc",x"405b",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"2563"),
(x"b9b2",x"4057",x"37cb",x"3950",x"a0dd",x"39fa",x"35bc",x"1ee4",x"b9bb",x"405b",x"37da",x"3950",x"a0dd",x"39fa",x"35c9",x"1fba",x"b9b2",x"405c",x"37cb",x"3950",x"a0dd",x"39fa",x"35c9",x"1d62"),
(x"b9b2",x"405c",x"37cb",x"b93c",x"95bc",x"3a0c",x"35eb",x"305f",x"b9a9",x"405b",x"37da",x"b93c",x"95bc",x"3a0c",x"35e3",x"3069",x"b9b2",x"4057",x"37cb",x"b93c",x"95bc",x"3a0c",x"35eb",x"307c"),
(x"b9cc",x"405b",x"37d1",x"b33b",x"b811",x"3aa5",x"3600",x"28cc",x"b9bb",x"405b",x"37da",x"b325",x"b878",x"3a63",x"35f3",x"28c6",x"b9b2",x"4057",x"37cb",x"1e0a",x"b823",x"3ad8",x"35ed",x"2927"),
(x"b994",x"405a",x"37cd",x"31e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"b996",x"404e",x"3791",x"3252",x"b816",x"3ab1",x"35d8",x"2a3e",x"b9b3",x"4051",x"37ad",x"a3bb",x"b81b",x"3add",x"35ee",x"29d8"),
(x"b996",x"404e",x"3791",x"3af1",x"b416",x"36d1",x"362a",x"31a9",x"b994",x"405a",x"37cd",x"3af6",x"b475",x"367c",x"362a",x"3154",x"b98f",x"405a",x"37ba",x"3b3a",x"b41e",x"357a",x"3622",x"315a"),
(x"b994",x"405a",x"37cd",x"358a",x"3a1b",x"385c",x"3649",x"253f",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9",x"b98f",x"405a",x"37ba",x"3926",x"39b7",x"3464",x"3645",x"24cf"),
(x"b996",x"404e",x"3791",x"3af1",x"b416",x"36d1",x"362a",x"31a9",x"b98f",x"405a",x"37ba",x"3b3a",x"b41e",x"357a",x"3622",x"315a",x"b98a",x"405b",x"379b",x"3aed",x"b3c2",x"3700",x"3617",x"3165"),
(x"b997",x"405c",x"3781",x"31af",x"3bdf",x"1c18",x"364b",x"22d3",x"b98a",x"405b",x"379b",x"3825",x"3acf",x"2d30",x"3640",x"2413",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b9c5",x"405d",x"3780",x"975f",x"3bfe",x"27c1",x"366e",x"22d4",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9",x"b9b2",x"405c",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"252a"),
(x"b9c5",x"405d",x"3780",x"975f",x"3bfe",x"27c1",x"366e",x"22d4",x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b9d3",x"405b",x"379f",x"b94b",x"39eb",x"af9d",x"367a",x"243b"),
(x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b9cc",x"405b",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"2563",x"b9d5",x"405b",x"37ba",x"b92f",x"39d8",x"32de",x"367a",x"24e0"),
(x"b9d5",x"405b",x"37ba",x"bb76",x"b463",x"3373",x"3596",x"345c",x"b9cc",x"405b",x"37d1",x"b9f1",x"b5fe",x"3870",x"35a0",x"3460",x"b9c9",x"404c",x"3787",x"bb76",x"b463",x"3373",x"35a0",x"342c"),
(x"b9c9",x"404c",x"3787",x"bb76",x"b463",x"3373",x"35a0",x"342c",x"b9d3",x"405b",x"379f",x"bbda",x"afe2",x"b0aa",x"358d",x"3457",x"b9d5",x"405b",x"37ba",x"bb76",x"b463",x"3373",x"3596",x"345c"),
(x"b98a",x"405b",x"379b",x"3aed",x"b3c2",x"3700",x"3617",x"3165",x"b992",x"404e",x"378f",x"35a5",x"b161",x"3b5d",x"3626",x"31a8",x"b996",x"404e",x"3791",x"3af1",x"b416",x"36d1",x"362a",x"31a9"),
(x"b990",x"404c",x"378e",x"3850",x"b763",x"39a2",x"3686",x"3221",x"b992",x"404e",x"378f",x"b67e",x"ac15",x"3b4a",x"3689",x"3214",x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5",x"b96c",x"4052",x"376e",x"392f",x"b7c9",x"38af",x"3668",x"3200",x"b990",x"404c",x"378e",x"3850",x"b763",x"39a2",x"3686",x"3221"),
(x"b964",x"4057",x"377a",x"39d4",x"b83f",x"36e9",x"3663",x"31e2",x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5",x"b961",x"405a",x"378b",x"3815",x"b8b5",x"3904",x"3664",x"31ce"),
(x"b964",x"4057",x"377a",x"39d4",x"b83f",x"36e9",x"3663",x"31e2",x"b959",x"405b",x"3775",x"3a72",x"b85a",x"3374",x"365a",x"31ce",x"b952",x"405c",x"3752",x"3a84",x"b81e",x"3444",x"364c",x"31d5"),
(x"b963",x"405b",x"3797",x"3b81",x"34c0",x"31b9",x"35aa",x"1ea6",x"b963",x"405d",x"3780",x"3bd2",x"3047",x"b134",x"35a0",x"1f3a",x"b961",x"405a",x"378b",x"3bd2",x"3047",x"b133",x"35aa",x"2000"),
(x"b964",x"4057",x"377a",x"3612",x"af46",x"3b58",x"362f",x"31de",x"b963",x"405d",x"3780",x"366b",x"ad14",x"3b4c",x"362f",x"31bd",x"b959",x"405b",x"3775",x"366b",x"ad14",x"3b4c",x"3626",x"31c9"),
(x"b975",x"405a",x"37b0",x"1fc8",x"3964",x"39e8",x"3641",x"2b5a",x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b",x"b963",x"405b",x"3797",x"3553",x"3a2a",x"3858",x"3650",x"2b30"),
(x"b991",x"405d",x"3777",x"b179",x"3b46",x"3611",x"3645",x"2c28",x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b",x"b98a",x"405b",x"379b",x"b5ee",x"392f",x"3951",x"363c",x"2bdc"),
(x"b991",x"405d",x"3777",x"b179",x"3b46",x"3611",x"3645",x"2c28",x"b98a",x"405b",x"379b",x"b5ee",x"392f",x"3951",x"363c",x"2bdc",x"b997",x"405c",x"3781",x"b106",x"3a66",x"38a1",x"363f",x"2c29"),
(x"b991",x"405d",x"3777",x"b179",x"3b46",x"3611",x"3645",x"2c28",x"b986",x"405d",x"375d",x"28bc",x"3bf3",x"2e92",x"3652",x"2c29",x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b"),
(x"b95b",x"405c",x"3777",x"391e",x"39e5",x"32f0",x"365f",x"2b4f",x"b95b",x"405d",x"3752",x"3410",x"3b92",x"3261",x"3669",x"2b9b",x"b959",x"405b",x"3775",x"39b9",x"391a",x"348e",x"3661",x"2b30"),
(x"b986",x"405d",x"375d",x"28bc",x"3bf3",x"2e92",x"3652",x"2c29",x"b981",x"405e",x"3752",x"24c2",x"3be9",x"30b5",x"3658",x"2c27",x"b963",x"405d",x"3780",x"2de3",x"3bd5",x"31ce",x"3658",x"2b68"),
(x"b95b",x"405c",x"3777",x"391e",x"39e5",x"32f0",x"365f",x"2b4f",x"b963",x"405d",x"3780",x"2de3",x"3bd5",x"31ce",x"3658",x"2b68",x"b95b",x"405d",x"3752",x"3410",x"3b92",x"3261",x"3669",x"2b9b"),
(x"b9f6",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"3639",x"3346",x"b9fd",x"3fd8",x"3786",x"baf1",x"b050",x"37a7",x"3637",x"331f",x"ba0d",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"361f",x"3321"),
(x"b9f0",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"363a",x"3356",x"b9f6",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"3639",x"3346",x"ba02",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"3620",x"334e"),
(x"b9f0",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"363a",x"3356",x"b9fa",x"3ff0",x"3752",x"b8fd",x"390a",x"3765",x"3622",x"3363",x"b9f2",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"3624",x"336f"),
(x"b9f6",x"3fa8",x"3752",x"bafd",x"b17a",x"3748",x"3634",x"328d",x"ba0d",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"361f",x"3321",x"b9fd",x"3fd8",x"3786",x"baf1",x"b050",x"37a7",x"3637",x"331f"),
(x"b9ee",x"3f8b",x"3752",x"bb0e",x"aeb1",x"3757",x"363e",x"323c",x"b9f6",x"3fa8",x"3752",x"bafd",x"b17a",x"3748",x"3634",x"328d",x"b9ed",x"3fa7",x"3777",x"bb1d",x"b0f4",x"36e3",x"3643",x"3291"),
(x"b9da",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"3644",x"3373",x"b9f2",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"3624",x"336f",x"b9d3",x"3fe5",x"3782",x"39d9",x"3972",x"a970",x"3645",x"3385"),
(x"b9ed",x"3fa7",x"3777",x"2b83",x"ac13",x"3bf8",x"35a9",x"31f0",x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9ed",x"3fa7",x"3777",x"2b83",x"ac13",x"3bf8",x"35a9",x"31f0",x"b9fd",x"3fd8",x"3786",x"a82c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9f5",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"35a5",x"327f",x"b9fd",x"3fd8",x"3786",x"a82c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9f6",x"3fe5",x"378d",x"ae26",x"ac9e",x"3bf1",x"35a6",x"32a5"),
(x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9f0",x"3fea",x"378e",x"ada8",x"257a",x"3bf7",x"35ab",x"32b3",x"b9e5",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"35b3",x"32b8"),
(x"b9e3",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"b9e5",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"35b3",x"32b8",x"b9da",x"3fea",x"378e",x"2e3a",x"2687",x"3bf5",x"35bc",x"32b1"),
(x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9da",x"3fea",x"378e",x"2e3a",x"2687",x"3bf5",x"35bc",x"32b1",x"b9d1",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"35c2",x"329a"),
(x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9cc",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"35c6",x"3293",x"b9cc",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9d1",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"35c2",x"329a",x"b9cc",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"35c6",x"3293"),
(x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9cc",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"b9d5",x"3faa",x"3777",x"ac2f",x"accc",x"3bf5",x"35bc",x"31f5",x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9cd",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"35c4",x"323e"),
(x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9d5",x"3faa",x"3777",x"ac2f",x"accc",x"3bf5",x"35bc",x"31f5",x"b9cc",x"3fa8",x"3777",x"abc1",x"ab62",x"3bf8",x"35c2",x"31f0"),
(x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9d5",x"3faa",x"3777",x"ac2f",x"accc",x"3bf5",x"35bc",x"31f5",x"b9da",x"3fab",x"3775",x"b235",x"abd2",x"3bd5",x"35b8",x"31f9"),
(x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9d7",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"35bd",x"3243",x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245"),
(x"b9d5",x"3fd5",x"3788",x"b21b",x"aee2",x"3bce",x"35bf",x"3274",x"b9d9",x"3fd5",x"3782",x"ae8f",x"aed5",x"3be9",x"35bb",x"3274",x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293"),
(x"b9d7",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"35be",x"3295",x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293",x"b9e1",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"35b6",x"32a0"),
(x"b9de",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"35b9",x"32a9",x"b9e1",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"35b6",x"32a0",x"b9e5",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9e3",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"b9e5",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9ec",x"3fe8",x"378f",x"2c49",x"b2ca",x"3bcc",x"35ad",x"32ab",x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"b9f5",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"35a5",x"327f",x"b9f1",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"35a9",x"329f",x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298"),
(x"b9e6",x"3fa9",x"3776",x"31d8",x"aa80",x"3bda",x"35af",x"31f3",x"b9f5",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"35a5",x"327f",x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245",x"b9da",x"3fab",x"3775",x"b235",x"abd2",x"3bd5",x"35b8",x"31f9",x"b9e3",x"3fa9",x"3773",x"2c3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"b9d9",x"3fd5",x"3782",x"ae8f",x"aed5",x"3be9",x"35bb",x"3274",x"b9dd",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"35b8",x"3245",x"b9f1",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293",x"b9d9",x"3fd5",x"3782",x"ae8f",x"aed5",x"3be9",x"35bb",x"3274",x"b9ee",x"3fe1",x"3785",x"2e7b",x"afea",x"3be5",x"35ac",x"3298"),
(x"b9e1",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"35b6",x"32a0",x"b9db",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"35ba",x"3293",x"b9ea",x"3fe5",x"3787",x"309e",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236",x"b9c9",x"3fa7",x"378a",x"bbec",x"2581",x"3053",x"35e3",x"3284",x"b9cb",x"3fa8",x"3783",x"bb1f",x"a907",x"3740",x"35e6",x"3285"),
(x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205",x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236",x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236"),
(x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec",x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205",x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203"),
(x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1",x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec",x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5"),
(x"b9c4",x"3fe1",x"37b6",x"ba64",x"b8cb",x"29c5",x"35e0",x"31dc",x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1",x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"b9c4",x"3fe1",x"37b6",x"ba64",x"b8cb",x"29c5",x"35e0",x"31dc",x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"b9c4",x"3fe1",x"37c1",x"badd",x"b464",x"b6f2",x"35dc",x"31dd",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe",x"b9ca",x"3fc5",x"37c6",x"baf7",x"2fd7",x"b79c",x"35d2",x"322a"),
(x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9ca",x"3fc5",x"37c6",x"baf7",x"2fd7",x"b79c",x"35d2",x"322a",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"b9ca",x"3f8a",x"3790",x"bbff",x"25e3",x"1e73",x"35da",x"32db",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e",x"b9c9",x"3fa8",x"37b2",x"bbe6",x"a832",x"30eb",x"35d4",x"327f"),
(x"b9ca",x"3fc3",x"37d1",x"bbf3",x"a804",x"2ec7",x"35cd",x"322c",x"b9c9",x"3fa8",x"37b2",x"bbe6",x"a832",x"30eb",x"35d4",x"327f",x"b9ca",x"3fa8",x"37a7",x"bbb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"b9ca",x"3fc3",x"37d1",x"bbf3",x"a804",x"2ec7",x"35cd",x"322c",x"b9ca",x"3fc5",x"37c6",x"baf7",x"2fd7",x"b79c",x"35d2",x"322a",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"b9ca",x"3fd3",x"37de",x"bbe7",x"9cea",x"30f2",x"35cc",x"31fd",x"b9ca",x"3fd3",x"37d4",x"bb45",x"2659",x"b6aa",x"35d0",x"31fe",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"b9c9",x"3fdf",x"37dc",x"bbdc",x"28a8",x"31d9",x"35d0",x"31db",x"b9ca",x"3fde",x"37d2",x"bb61",x"add1",x"b5fd",x"35d3",x"31e0",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"b9ca",x"3fe6",x"37cc",x"bbf2",x"2956",x"2ec5",x"35d9",x"31c8",x"b9cb",x"3fe3",x"37c8",x"bb6f",x"b4b7",x"b314",x"35d9",x"31d1",x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"b9cb",x"3fe7",x"37a7",x"bbff",x"1ec2",x"2532",x"35e8",x"31ca",x"b9cb",x"3fe8",x"37b8",x"bbfd",x"2581",x"2a45",x"35e1",x"31c5",x"b9cb",x"3fe6",x"37b7",x"bb9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"b9cb",x"3fe0",x"378e",x"bbf9",x"1818",x"2d46",x"35f0",x"31e1",x"b9cb",x"3fe7",x"37a7",x"bbff",x"1ec2",x"2532",x"35e8",x"31ca",x"b9cb",x"3fe4",x"37aa",x"bb36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"b9cc",x"3fd4",x"3784",x"bbeb",x"a025",x"3082",x"35f2",x"3204",x"b9cb",x"3fe0",x"378e",x"bbf9",x"1818",x"2d46",x"35f0",x"31e1",x"b9cb",x"3fde",x"3799",x"bb18",x"b180",x"36da",x"35ec",x"31e5"),
(x"b9cd",x"3fc3",x"377f",x"bbd2",x"a2f6",x"32b9",x"35f0",x"3237",x"b9cc",x"3fd4",x"3784",x"bbeb",x"a025",x"3082",x"35f2",x"3204",x"b9cb",x"3fd4",x"3790",x"bada",x"acd9",x"3814",x"35ed",x"3203"),
(x"b9cb",x"3fc2",x"378b",x"bacd",x"a90b",x"3833",x"35eb",x"3236",x"b9cb",x"3fa8",x"3783",x"bb1f",x"a907",x"3740",x"35e6",x"3285",x"b9cc",x"3fa8",x"3777",x"bbc7",x"a659",x"336e",x"35eb",x"3285"),
(x"b9c9",x"3fa7",x"378a",x"bbec",x"2581",x"3053",x"35e3",x"3284",x"b9c8",x"3fa9",x"379f",x"bbfa",x"2c56",x"a7a7",x"35dc",x"327e",x"b9ca",x"3f8a",x"3790",x"bbff",x"25e3",x"1e73",x"35da",x"32db"),
(x"b9c8",x"3fa9",x"379f",x"bbfa",x"2c56",x"a7a7",x"35dc",x"327e",x"b9c9",x"3fa7",x"378a",x"bbec",x"2581",x"3053",x"35e3",x"3284",x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236"),
(x"b9c4",x"3fc5",x"37ba",x"bbe1",x"2c8e",x"b0f7",x"35d8",x"3228",x"b9c6",x"3fc2",x"3794",x"bbb1",x"2446",x"345f",x"35e6",x"3236",x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205"),
(x"b9c4",x"3fd3",x"37c9",x"bbcf",x"29e6",x"b2c7",x"35d6",x"3200",x"b9c6",x"3fd3",x"3798",x"bbae",x"a64c",x"3470",x"35e8",x"3205",x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec"),
(x"b9c4",x"3fdd",x"37c7",x"bb8c",x"a66c",x"b548",x"35d9",x"31e6",x"b9c4",x"3fdc",x"37a3",x"bbad",x"a9fd",x"346f",x"35e5",x"31ec",x"b9c4",x"3fe0",x"37ac",x"bb37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"b9c9",x"3fa8",x"37b2",x"b870",x"b1f2",x"3a7c",x"35f5",x"3500",x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b9ab",x"3f87",x"37c0",x"248e",x"b255",x"3bd7",x"35d8",x"352f"),
(x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b9c9",x"3fa8",x"37b2",x"b870",x"b1f2",x"3a7c",x"35f5",x"3500",x"b9ca",x"3fc3",x"37d1",x"b885",x"b324",x"3a5a",x"35f4",x"34d4"),
(x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b9ca",x"3fc3",x"37d1",x"b885",x"b324",x"3a5a",x"35f4",x"34d4",x"b9ca",x"3fd3",x"37de",x"b89a",x"ad78",x"3a82",x"35f2",x"34bc"),
(x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b9ca",x"3fd3",x"37de",x"b89a",x"ad78",x"3a82",x"35f2",x"34bc",x"b9c9",x"3fdf",x"37dc",x"b869",x"323c",x"3a7d",x"35f0",x"34aa"),
(x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b9c9",x"3fdf",x"37dc",x"b869",x"323c",x"3a7d",x"35f0",x"34aa",x"b9ca",x"3fe6",x"37cc",x"b783",x"398b",x"385f",x"35ef",x"349c"),
(x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495",x"b9aa",x"3feb",x"37e2",x"1953",x"3ada",x"3821",x"35d7",x"349e",x"b9ca",x"3fe6",x"37cc",x"b783",x"398b",x"385f",x"35ef",x"349c"),
(x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e",x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495",x"b9cb",x"3fe8",x"37b8",x"b5d5",x"3b70",x"2a94",x"35f1",x"3494"),
(x"b9c2",x"3fe7",x"379c",x"b620",x"3a0a",x"b841",x"35ed",x"3488",x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e",x"b9cb",x"3fe7",x"37a7",x"b572",x"3a96",x"b740",x"35f3",x"348e"),
(x"b9d1",x"3fe2",x"378c",x"39d1",x"382c",x"3722",x"364c",x"3387",x"b9d3",x"3fe5",x"3782",x"39d9",x"3972",x"a970",x"3645",x"3385",x"b9cb",x"3fe1",x"3786",x"388d",x"3867",x"38e2",x"364c",x"3391"),
(x"b9cb",x"3fe1",x"3786",x"b81b",x"39f5",x"36d0",x"35f8",x"347e",x"b9c8",x"3fe1",x"378b",x"b994",x"399e",x"b082",x"35f6",x"3480",x"b9cb",x"3fe0",x"378e",x"b81d",x"395a",x"b849",x"35f9",x"3481"),
(x"b949",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"35ab",x"2e93",x"b959",x"3fd8",x"3786",x"3ad9",x"b071",x"37f4",x"35c2",x"2e97",x"b960",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"35c4",x"2e47"),
(x"b953",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"35ab",x"2e39",x"b960",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"35c4",x"2e47",x"b966",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"35c6",x"2e27"),
(x"b966",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"35c6",x"2e27",x"b971",x"3fec",x"378f",x"a8a8",x"3b7d",x"3597",x"35ca",x"2e09",x"b964",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"35af",x"2df7"),
(x"b959",x"3fd8",x"3786",x"3ad9",x"b071",x"37f4",x"35c2",x"2e97",x"b949",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"35ab",x"2e93",x"b960",x"3fa8",x"3752",x"3adc",x"b152",x"37c7",x"35c0",x"2fbb"),
(x"b96a",x"3fa6",x"3775",x"3acd",x"b078",x"380f",x"35cf",x"2fb9",x"b960",x"3fa8",x"3752",x"3adc",x"b152",x"37c7",x"35c0",x"2fbb",x"b965",x"3f8b",x"3752",x"3ab6",x"ad4f",x"384c",x"35c9",x"302f"),
(x"b983",x"3fe5",x"3782",x"b9dc",x"3971",x"a62b",x"35d1",x"2dca",x"b964",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"35af",x"2df7",x"b97c",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e",x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2",x"b96a",x"3fa6",x"3775",x"2b9a",x"acf0",x"3bf6",x"3611",x"30d8"),
(x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2",x"b961",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"360d",x"3046",x"b959",x"3fd8",x"3786",x"2e54",x"ae94",x"3beb",x"3607",x"3046"),
(x"b959",x"3fd8",x"3786",x"2e54",x"ae94",x"3beb",x"3607",x"3046",x"b961",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"360d",x"3046",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026"),
(x"b960",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"360d",x"3020",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a",x"b972",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"361b",x"3016",x"b971",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"361b",x"300d"),
(x"b972",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"361b",x"3016",x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b97c",x"3fea",x"378e",x"ae3a",x"2687",x"3bf5",x"3623",x"3014"),
(x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f",x"b985",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f",x"b989",x"3fe0",x"378b",x"af00",x"af3d",x"3be6",x"362d",x"3032",x"b985",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051",x"b98a",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"362d",x"3054",x"b989",x"3fe0",x"378b",x"af00",x"af3d",x"3be6",x"362d",x"3032"),
(x"b98a",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"362d",x"3054",x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082"),
(x"b989",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"362b",x"3087",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082",x"b981",x"3faa",x"3777",x"2c34",x"acb2",x"3bf5",x"3623",x"30d0"),
(x"b989",x"3fa8",x"3777",x"26fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"b981",x"3faa",x"3777",x"2c34",x"acb2",x"3bf5",x"3623",x"30d0",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"b97c",x"3fab",x"3775",x"3227",x"ab9d",x"3bd6",x"361f",x"30cb",x"b981",x"3faa",x"3777",x"2c34",x"acb2",x"3bf5",x"3623",x"30d0",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082"),
(x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080",x"b97f",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"3624",x"3082",x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051"),
(x"b981",x"3fd5",x"3788",x"321b",x"aee2",x"3bce",x"3626",x"3051",x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f",x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"b97f",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"3625",x"302f",x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b975",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"361d",x"3025"),
(x"b978",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"3620",x"301c",x"b972",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"361b",x"3016",x"b971",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"361a",x"3022"),
(x"b971",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"361a",x"3022",x"b972",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"361b",x"3016",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b96a",x"3fe8",x"378f",x"ac4b",x"b2ca",x"3bcc",x"3615",x"301a",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026"),
(x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b965",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"3611",x"3026",x"b961",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"360d",x"3046"),
(x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b961",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"360d",x"3046",x"b970",x"3fa9",x"3776",x"affb",x"abfc",x"3beb",x"3616",x"30d2"),
(x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"b977",x"3f89",x"376f",x"2217",x"a8a5",x"3bfe",x"3619",x"312e",x"b983",x"3f89",x"3770",x"2b4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"b973",x"3fa9",x"3773",x"ac2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"b97c",x"3fab",x"3775",x"3227",x"ab9d",x"3bd6",x"361f",x"30cb",x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080"),
(x"b964",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"3610",x"3048",x"b979",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"361f",x"3080",x"b97d",x"3fd5",x"3782",x"2e8f",x"aed5",x"3be9",x"3623",x"3050"),
(x"b968",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"3614",x"302d",x"b97d",x"3fd5",x"3782",x"2e8f",x"aed5",x"3be9",x"3623",x"3050",x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"b96c",x"3fe5",x"3787",x"b09e",x"b24e",x"3bc1",x"3616",x"3024",x"b97b",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"3621",x"3032",x"b975",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"361d",x"3025"),
(x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4",x"b98d",x"3fa8",x"378a",x"3be0",x"2467",x"319c",x"360d",x"31c3",x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"b98b",x"3fc2",x"378b",x"3a70",x"a9d2",x"38bb",x"3615",x"3211",x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211",x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242",x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b"),
(x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263",x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268"),
(x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268",x"b991",x"3fe2",x"37b7",x"3a93",x"b88d",x"2474",x"360a",x"326f"),
(x"b991",x"3fe2",x"37b7",x"3a93",x"b88d",x"2474",x"360a",x"326f",x"b991",x"3fe1",x"37c3",x"3b15",x"b384",x"b669",x"3606",x"326c",x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277"),
(x"b991",x"3fe1",x"37c3",x"3b15",x"b384",x"b669",x"3606",x"326c",x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b98c",x"3fd3",x"37d2",x"3a75",x"2987",x"b8b5",x"35fc",x"3249"),
(x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b991",x"3fc5",x"37be",x"3beb",x"2c4d",x"b006",x"3601",x"321f",x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e"),
(x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e",x"b991",x"3fc5",x"37be",x"3beb",x"2c4d",x"b006",x"3601",x"321f",x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9"),
(x"b98c",x"3fa8",x"37b0",x"3bfa",x"a217",x"2ca7",x"35ff",x"31c8",x"b98c",x"3fa9",x"37a5",x"3bef",x"2703",x"afec",x"3603",x"31c9",x"b98b",x"3f85",x"378d",x"3bff",x"2504",x"1d6d",x"3604",x"3160"),
(x"b98c",x"3fa9",x"37a5",x"3bef",x"2703",x"afec",x"3603",x"31c9",x"b98c",x"3fa8",x"37b0",x"3bfa",x"a217",x"2ca7",x"35ff",x"31c8",x"b98c",x"3fc3",x"37d0",x"3bff",x"a2f6",x"24f7",x"35f8",x"321b"),
(x"b98c",x"3fc4",x"37c6",x"3af8",x"2fc1",x"b79c",x"35fc",x"321e",x"b98c",x"3fc3",x"37d0",x"3bff",x"a2f6",x"24f7",x"35f8",x"321b",x"b98c",x"3fd3",x"37dc",x"3bff",x"15bc",x"a673",x"35f8",x"324b"),
(x"b98c",x"3fd3",x"37dc",x"3bff",x"15bc",x"a673",x"35f8",x"324b",x"b98c",x"3fde",x"37db",x"3bff",x"1953",x"2560",x"35fb",x"326b",x"b98c",x"3fdd",x"37d0",x"3b3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"b98c",x"3fde",x"37db",x"3bff",x"1953",x"2560",x"35fb",x"326b",x"b98c",x"3fe6",x"37cd",x"3bf7",x"29c5",x"2d1b",x"3603",x"327f",x"b98b",x"3fe3",x"37c9",x"3b72",x"b453",x"b3d7",x"3604",x"3277"),
(x"b98c",x"3fe6",x"37cd",x"3bf7",x"29c5",x"2d1b",x"3603",x"327f",x"b98b",x"3fe8",x"37b8",x"3bfd",x"1edc",x"29f0",x"360c",x"3283",x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b"),
(x"b98b",x"3fe5",x"37b7",x"3bb2",x"b454",x"25bc",x"360b",x"327b",x"b98b",x"3fe8",x"37b8",x"3bfd",x"1edc",x"29f0",x"360c",x"3283",x"b98b",x"3fe7",x"37a7",x"3bff",x"0cea",x"269a",x"3612",x"327d"),
(x"b98b",x"3fe4",x"37aa",x"3b50",x"b4c5",x"3465",x"3610",x"3274",x"b98b",x"3fe7",x"37a7",x"3bff",x"0cea",x"269a",x"3612",x"327d",x"b98a",x"3fe0",x"378e",x"3bf8",x"15bc",x"2d81",x"361b",x"3266"),
(x"b98a",x"3fd4",x"3784",x"3bea",x"a025",x"3095",x"361c",x"3243",x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b98a",x"3fde",x"3798",x"3b1d",x"b165",x"36cb",x"3617",x"3263"),
(x"b98b",x"3fd4",x"3790",x"3adf",x"ac91",x"380d",x"3618",x"3244",x"b98a",x"3fd4",x"3784",x"3bea",x"a025",x"3095",x"361c",x"3243",x"b989",x"3fc3",x"377f",x"3bce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"b98b",x"3fa8",x"3782",x"3b3c",x"a8f7",x"36cb",x"3611",x"31c4",x"b98b",x"3fc2",x"378b",x"3a70",x"a9d2",x"38bb",x"3615",x"3211",x"b989",x"3fc3",x"377f",x"3bce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9",x"b98d",x"3fa8",x"378a",x"3be0",x"2467",x"319c",x"360d",x"31c3",x"b98b",x"3f89",x"3770",x"3bf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"b98e",x"3fa9",x"37a1",x"3bf1",x"2c5d",x"ae42",x"3605",x"31c9",x"b991",x"3fc5",x"37be",x"3beb",x"2c4d",x"b006",x"3601",x"321f",x"b990",x"3fc2",x"3794",x"3bcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"b991",x"3fc5",x"37be",x"3beb",x"2c4d",x"b006",x"3601",x"321f",x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b990",x"3fd3",x"3798",x"3bbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"b992",x"3fd3",x"37c9",x"3bd1",x"2963",x"b2aa",x"3601",x"3246",x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b992",x"3fdc",x"37a3",x"3bc0",x"accc",x"3386",x"3610",x"325b"),
(x"b991",x"3fdd",x"37c9",x"3b95",x"ac0e",x"b4fe",x"3603",x"3262",x"b991",x"3fe1",x"37c3",x"3b15",x"b384",x"b669",x"3606",x"326c",x"b991",x"3fe0",x"37ac",x"3b6f",x"b421",x"3438",x"360e",x"3268"),
(x"b9ab",x"3f87",x"37c0",x"248e",x"b255",x"3bd7",x"35d8",x"352f",x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b98c",x"3fa8",x"37b0",x"387f",x"b1e6",x"3a73",x"35ba",x"3500"),
(x"b9aa",x"3fa8",x"37dc",x"2217",x"b41e",x"3bba",x"35d7",x"34fc",x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b98c",x"3fc3",x"37d0",x"3896",x"b2c0",x"3a54",x"35bb",x"34d5"),
(x"b9ac",x"3fc7",x"3800",x"231d",x"b311",x"3bcd",x"35d8",x"34cd",x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b98c",x"3fd3",x"37dc",x"3892",x"ade1",x"3a86",x"35bc",x"34bc"),
(x"b9ab",x"3fd7",x"3804",x"2194",x"28d6",x"3bfe",x"35d8",x"34b8",x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b98c",x"3fde",x"37db",x"3885",x"3126",x"3a79",x"35be",x"34ab"),
(x"b9aa",x"3fe6",x"37fd",x"212b",x"36f9",x"3b33",x"35d7",x"34a8",x"b9aa",x"3feb",x"37e2",x"1953",x"3ada",x"3821",x"35d7",x"349e",x"b98c",x"3fe6",x"37cd",x"37e6",x"396d",x"3859",x"35bf",x"349d"),
(x"b98c",x"3fe6",x"37cd",x"37e6",x"396d",x"3859",x"35bf",x"349d",x"b9aa",x"3feb",x"37e2",x"1953",x"3ada",x"3821",x"35d7",x"349e",x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495"),
(x"b98b",x"3fe8",x"37b8",x"361b",x"3b60",x"2bbe",x"35be",x"3495",x"b9aa",x"3fee",x"37c9",x"1b5f",x"3bbd",x"340d",x"35d7",x"3495",x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e"),
(x"b98b",x"3fe7",x"37a7",x"3619",x"3a76",x"b730",x"35bb",x"348f",x"b9aa",x"3fee",x"37b3",x"29ed",x"3baa",x"b482",x"35d7",x"348e",x"b993",x"3fe4",x"3789",x"3646",x"3a25",x"b80b",x"35bd",x"3481"),
(x"b98c",x"3fe1",x"3782",x"b8d3",x"3873",x"3892",x"35d6",x"2daa",x"b983",x"3fe5",x"3782",x"b9dc",x"3971",x"a62b",x"35d1",x"2dca",x"b985",x"3fe2",x"378c",x"b9bb",x"383c",x"3743",x"35d7",x"2dc5"),
(x"b98e",x"3fe1",x"378b",x"38bd",x"3a6d",x"2bf2",x"35b7",x"3482",x"b98c",x"3fe1",x"3782",x"3865",x"3aa9",x"2c27",x"35b6",x"347e",x"b989",x"3fe0",x"378b",x"3862",x"3a94",x"30e6",x"35b3",x"3481"),
(x"b965",x"3f8b",x"3752",x"3ab6",x"ad4f",x"384c",x"35c9",x"302f",x"b96a",x"3f6f",x"3752",x"3ae4",x"ad23",x"3802",x"35d2",x"307e",x"b970",x"3f7e",x"376e",x"3abb",x"aad9",x"384d",x"35d9",x"3052"),
(x"b970",x"3f88",x"376d",x"303d",x"a8e0",x"3bec",x"3614",x"3130",x"b970",x"3f7e",x"376e",x"312d",x"203f",x"3be4",x"3613",x"314f",x"b979",x"3f83",x"3770",x"2e2b",x"280b",x"3bf5",x"361a",x"3141"),
(x"b9e4",x"3f7a",x"376e",x"bb00",x"aaa4",x"37b3",x"364e",x"320e",x"b9ea",x"3f6e",x"3752",x"bb03",x"aae6",x"37a4",x"3646",x"31e8",x"b9ee",x"3f8b",x"3752",x"bb0e",x"aeb1",x"3757",x"363e",x"323c"),
(x"b9df",x"3f8b",x"376f",x"8cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"b9d3",x"3f8b",x"3770",x"ac6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"b9d3",x"3f7f",x"3770",x"a93f",x"1af6",x"3bfe",x"35ba",x"3179"),
(x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9",x"b9e5",x"4030",x"37b3",x"b48b",x"3a03",x"38c2",x"3611",x"2fda",x"b9f8",x"4030",x"3794",x"b663",x"3a38",x"37c6",x"3623",x"2fe3"),
(x"ba01",x"4030",x"377a",x"b864",x"3a40",x"34bc",x"3630",x"2fdb",x"ba08",x"4031",x"3752",x"b890",x"3a28",x"3491",x"363e",x"2fc0",x"b9fd",x"4033",x"3752",x"b24d",x"3bb2",x"31fb",x"3638",x"2fa0"),
(x"b9f6",x"402c",x"377c",x"b9ed",x"b7fd",x"372e",x"364a",x"3429",x"b9f5",x"4028",x"3752",x"baa2",x"b726",x"355e",x"363e",x"341a",x"ba08",x"4031",x"3752",x"ba9b",x"b7a9",x"34c2",x"3635",x"3436"),
(x"b9f6",x"402c",x"377c",x"b9ed",x"b7fd",x"372e",x"364a",x"3429",x"b9ed",x"4027",x"376e",x"b8ec",x"b7ef",x"38e6",x"364a",x"3418",x"b9f5",x"4028",x"3752",x"baa2",x"b726",x"355e",x"363e",x"341a"),
(x"b9e5",x"4030",x"37b3",x"b89d",x"b810",x"391d",x"3662",x"3434",x"b9f6",x"402c",x"377c",x"b9ed",x"b7fd",x"372e",x"364a",x"3429",x"b9f8",x"4030",x"3794",x"b839",x"b89f",x"38fa",x"3650",x"3436"),
(x"b9e5",x"4030",x"37b3",x"b89d",x"b810",x"391d",x"3662",x"3434",x"b9ed",x"4027",x"376e",x"b8ec",x"b7ef",x"38e6",x"364a",x"3418",x"b9f6",x"402c",x"377c",x"b9ed",x"b7fd",x"372e",x"364a",x"3429"),
(x"b9d3",x"4031",x"379f",x"354f",x"39c9",x"38d8",x"360b",x"2fa1",x"b9dc",x"4030",x"37ae",x"335d",x"39d9",x"3923",x"360d",x"2fc2",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"b9df",x"4033",x"3752",x"9d04",x"3bf5",x"2e94",x"3627",x"2f61",x"b9c5",x"4033",x"3780",x"2cce",x"3bc5",x"3334",x"360d",x"2f61",x"b9e1",x"4032",x"37a2",x"ab58",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349",x"b994",x"4030",x"37cd",x"358a",x"3a1b",x"385c",x"3649",x"3358",x"b9a9",x"4030",x"37da",x"3146",x"3a67",x"389c",x"3659",x"3362"),
(x"b9b2",x"4031",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"3355",x"b9bb",x"4030",x"37da",x"ae09",x"3b05",x"3784",x"3667",x"3363",x"b9cc",x"4030",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"335c"),
(x"b9b3",x"4026",x"37ad",x"a3bb",x"b81b",x"3add",x"3677",x"311b",x"b9c9",x"4021",x"3787",x"b409",x"b819",x"3a90",x"3689",x"3140",x"b9cc",x"4030",x"37d1",x"b33b",x"b811",x"3aa5",x"3689",x"30d9"),
(x"b9cc",x"4030",x"37d1",x"b33b",x"b811",x"3aa5",x"3689",x"30d9",x"b9b2",x"402d",x"37cb",x"1e0a",x"b823",x"3ad8",x"3676",x"30ef",x"b9b3",x"4026",x"37ad",x"a3bb",x"b81b",x"3add",x"3677",x"311b"),
(x"b994",x"4030",x"37cd",x"31e7",x"b81a",x"3ab5",x"365e",x"30e1",x"b9b2",x"402d",x"37cb",x"1e0a",x"b823",x"3ad8",x"3676",x"30ef",x"b9a9",x"4030",x"37da",x"324d",x"b8ad",x"3a4b",x"366f",x"30d9"),
(x"b994",x"4030",x"37cd",x"31e7",x"b81a",x"3ab5",x"365e",x"30e1",x"b9b3",x"4026",x"37ad",x"a3bb",x"b81b",x"3add",x"3677",x"311b",x"b9b2",x"402d",x"37cb",x"1e0a",x"b823",x"3ad8",x"3676",x"30ef"),
(x"b98a",x"4030",x"379b",x"3825",x"3acf",x"2d30",x"3640",x"3332",x"b98f",x"4030",x"37ba",x"3926",x"39b7",x"3465",x"3645",x"334a",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"b9c5",x"4033",x"3780",x"96f6",x"3bfe",x"27c1",x"366e",x"331d",x"b997",x"4032",x"3781",x"31af",x"3bdf",x"1c18",x"364b",x"331d",x"b998",x"4032",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"b9ce",x"4032",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"3343",x"b9d5",x"4030",x"37ba",x"b92f",x"39d8",x"32de",x"367a",x"334c",x"b9d3",x"4031",x"379f",x"b94c",x"39eb",x"af9a",x"367a",x"3337"),
(x"b98a",x"4030",x"379b",x"b65b",x"ac2a",x"3b52",x"366b",x"3506",x"b975",x"4030",x"37b0",x"35ad",x"b6ed",x"3aa0",x"3659",x"3502",x"b990",x"4021",x"378e",x"34a7",x"b630",x"3b00",x"3668",x"3531"),
(x"b96c",x"4028",x"376e",x"392f",x"b7c9",x"38af",x"3649",x"3520",x"b98a",x"4021",x"377f",x"392b",x"b843",x"385f",x"3662",x"3532",x"b990",x"4021",x"378e",x"34a7",x"b630",x"3b00",x"3668",x"3531"),
(x"b961",x"402f",x"378b",x"3815",x"b8b5",x"3904",x"3646",x"3507",x"b975",x"4030",x"37b0",x"35ad",x"b6ed",x"3aa0",x"3659",x"3502",x"b963",x"4030",x"3797",x"3810",x"b8bd",x"3900",x"3649",x"3503"),
(x"b964",x"402c",x"377a",x"39d4",x"b83f",x"36e9",x"3645",x"3511",x"b96c",x"4028",x"376e",x"392f",x"b7c9",x"38af",x"3649",x"3520",x"b975",x"4030",x"37b0",x"35ad",x"b6ed",x"3aa0",x"3659",x"3502"),
(x"b964",x"402c",x"377a",x"39d4",x"b83f",x"36e9",x"3645",x"3511",x"b966",x"4029",x"3752",x"3a92",x"b7fc",x"346b",x"363e",x"3522",x"b96c",x"4028",x"376e",x"392f",x"b7c9",x"38af",x"3649",x"3520"),
(x"b964",x"402c",x"377a",x"39d4",x"b83f",x"36e9",x"3645",x"3511",x"b952",x"4031",x"3752",x"3a84",x"b81e",x"3444",x"362e",x"350b",x"b966",x"4029",x"3752",x"3a92",x"b7fc",x"346b",x"363e",x"3522"),
(x"b963",x"4032",x"3780",x"3bd2",x"3047",x"b134",x"35bb",x"2006",x"b964",x"402c",x"377a",x"3b82",x"286a",x"b57a",x"35ac",x"20d4",x"b961",x"402f",x"378b",x"3bd2",x"3047",x"b133",x"35b6",x"210c"),
(x"b963",x"4032",x"3780",x"366c",x"ad14",x"3b4c",x"362f",x"31e1",x"b95b",x"4032",x"3777",x"3827",x"3037",x"3ac1",x"3628",x"31e5",x"b959",x"4030",x"3775",x"366c",x"ad14",x"3b4c",x"3626",x"31ed"),
(x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f",x"b963",x"4032",x"3780",x"2de3",x"3bd5",x"31ce",x"3625",x"2e26",x"b963",x"4030",x"3797",x"3553",x"3a2a",x"3859",x"361e",x"2e0a"),
(x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f",x"b975",x"4030",x"37b0",x"1fc8",x"3964",x"39e8",x"360f",x"2e1f",x"b98a",x"4030",x"379b",x"b5ee",x"392f",x"3951",x"3609",x"2e60"),
(x"b986",x"4033",x"375d",x"28bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"b963",x"4032",x"3780",x"2de3",x"3bd5",x"31ce",x"3625",x"2e26",x"b97a",x"4032",x"37a0",x"11bc",x"3b79",x"35b5",x"3613",x"2e3f"),
(x"b95b",x"4033",x"3752",x"3410",x"3b92",x"3261",x"3637",x"2e3f",x"b952",x"4031",x"3752",x"38c8",x"39c1",x"35a4",x"363b",x"2e1f",x"b959",x"4030",x"3775",x"39b9",x"391a",x"348e",x"362e",x"2e0a"),
(x"b981",x"4033",x"3752",x"24c2",x"3be9",x"30b5",x"3625",x"2e99",x"b95b",x"4033",x"3752",x"3410",x"3b92",x"3261",x"3637",x"2e3f",x"b963",x"4032",x"3780",x"2de3",x"3bd5",x"31ce",x"3625",x"2e26"),
(x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db",x"b9e5",x"405b",x"37b3",x"b48b",x"3a04",x"38c2",x"3648",x"33ec",x"b9f8",x"405b",x"3794",x"b663",x"3a38",x"37c6",x"3659",x"33f1"),
(x"ba01",x"405b",x"377a",x"b865",x"3a40",x"34bc",x"3665",x"33ed",x"ba08",x"405c",x"3752",x"b890",x"3a28",x"3491",x"3673",x"33df",x"b9fd",x"405e",x"3752",x"b24d",x"3bb2",x"31fb",x"366d",x"33ce"),
(x"b9f6",x"4057",x"377c",x"b9d5",x"b835",x"3700",x"365a",x"32ee",x"b9f5",x"4054",x"3752",x"ba92",x"b7a6",x"34f5",x"364e",x"32d1",x"ba08",x"405c",x"3752",x"ba92",x"b7f9",x"346d",x"3646",x"3307"),
(x"b9f6",x"4057",x"377c",x"b9d5",x"b835",x"3700",x"365a",x"32ee",x"b9ed",x"4053",x"376e",x"b8f6",x"b815",x"38c2",x"365a",x"32ce",x"b9f5",x"4054",x"3752",x"ba92",x"b7a6",x"34f5",x"364e",x"32d1"),
(x"b9e5",x"405b",x"37b3",x"b8ae",x"b826",x"38fc",x"3671",x"3303",x"b9f6",x"4057",x"377c",x"b9d5",x"b835",x"3700",x"365a",x"32ee",x"b9f8",x"405b",x"3794",x"b839",x"b89f",x"38fa",x"3660",x"3309"),
(x"b9e5",x"405b",x"37b3",x"b8ae",x"b826",x"38fc",x"3671",x"3303",x"b9ed",x"4053",x"376e",x"b8f6",x"b815",x"38c2",x"365a",x"32ce",x"b9f6",x"4057",x"377c",x"b9d5",x"b835",x"3700",x"365a",x"32ee"),
(x"b9d3",x"405b",x"379f",x"354f",x"39c9",x"38d8",x"3642",x"33cf",x"b9dc",x"405b",x"37ae",x"335d",x"39d9",x"3923",x"3644",x"33e0",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db"),
(x"b9df",x"405e",x"3752",x"9d04",x"3bf5",x"2e94",x"365d",x"33ae",x"b9c5",x"405d",x"3780",x"2cce",x"3bc5",x"3335",x"3644",x"33ae",x"b9e1",x"405d",x"37a2",x"ab58",x"3bb1",x"344b",x"364b",x"33db"),
(x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9",x"b994",x"405a",x"37cd",x"358a",x"3a1b",x"385c",x"3649",x"253f",x"b9a9",x"405b",x"37da",x"3146",x"3a67",x"389c",x"3659",x"2595"),
(x"b9b2",x"405c",x"37cb",x"a393",x"3b79",x"35b2",x"3660",x"252a",x"b9bb",x"405b",x"37da",x"ae09",x"3b05",x"3784",x"3667",x"2596",x"b9cc",x"405b",x"37d1",x"b1ec",x"3b16",x"36cd",x"3674",x"2563"),
(x"b9b3",x"4051",x"37ad",x"a3bb",x"b81b",x"3add",x"35ee",x"29d8",x"b9c9",x"404c",x"3787",x"b409",x"b819",x"3a90",x"3600",x"2a6b",x"b9cc",x"405b",x"37d1",x"b33b",x"b811",x"3aa5",x"3600",x"28cc"),
(x"b9cc",x"405b",x"37d1",x"b33b",x"b811",x"3aa5",x"3600",x"28cc",x"b9b2",x"4057",x"37cb",x"1e0a",x"b823",x"3ad8",x"35ed",x"2927",x"b9b3",x"4051",x"37ad",x"a3bb",x"b81b",x"3add",x"35ee",x"29d8"),
(x"b994",x"405a",x"37cd",x"31e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"b9b2",x"4057",x"37cb",x"1e0a",x"b823",x"3ad8",x"35ed",x"2927",x"b9a9",x"405b",x"37da",x"324d",x"b8ad",x"3a4b",x"35e6",x"28d0"),
(x"b994",x"405a",x"37cd",x"31e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"b9b3",x"4051",x"37ad",x"a3bb",x"b81b",x"3add",x"35ee",x"29d8",x"b9b2",x"4057",x"37cb",x"1e0a",x"b823",x"3ad8",x"35ed",x"2927"),
(x"b98a",x"405b",x"379b",x"3825",x"3acf",x"2d30",x"3640",x"2413",x"b98f",x"405a",x"37ba",x"3926",x"39b7",x"3464",x"3645",x"24cf",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"b9c5",x"405d",x"3780",x"96f6",x"3bfe",x"27c1",x"366e",x"22d4",x"b997",x"405c",x"3781",x"31af",x"3bdf",x"1c18",x"364b",x"22d3",x"b998",x"405c",x"37bd",x"30a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"b9ce",x"405d",x"37b1",x"af93",x"3bda",x"30c0",x"3674",x"249a",x"b9d5",x"405b",x"37ba",x"b92f",x"39d8",x"32de",x"367a",x"24e0",x"b9d3",x"405b",x"379f",x"b94b",x"39eb",x"af9d",x"367a",x"243b"),
(x"b992",x"404e",x"378f",x"b67e",x"ac15",x"3b4a",x"3689",x"3214",x"b98a",x"405b",x"379b",x"b713",x"a8bc",x"3b2b",x"3689",x"31cb",x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"b96c",x"4052",x"376e",x"392f",x"b7c9",x"38af",x"3668",x"3200",x"b98a",x"404c",x"377f",x"392b",x"b843",x"385f",x"3680",x"3225",x"b990",x"404c",x"378e",x"3850",x"b763",x"39a2",x"3686",x"3221"),
(x"b961",x"405a",x"378b",x"3815",x"b8b5",x"3904",x"3664",x"31ce",x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5",x"b963",x"405b",x"3797",x"3810",x"b8bd",x"3900",x"3668",x"31c5"),
(x"b964",x"4057",x"377a",x"39d4",x"b83f",x"36e9",x"3663",x"31e2",x"b96c",x"4052",x"376e",x"392f",x"b7c9",x"38af",x"3668",x"3200",x"b975",x"405a",x"37b0",x"3564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"b964",x"4057",x"377a",x"39d4",x"b83f",x"36e9",x"3663",x"31e2",x"b966",x"4053",x"3752",x"3a92",x"b7fc",x"346c",x"365c",x"3204",x"b96c",x"4052",x"376e",x"392f",x"b7c9",x"38af",x"3668",x"3200"),
(x"b964",x"4057",x"377a",x"39d4",x"b83f",x"36e9",x"3663",x"31e2",x"b952",x"405c",x"3752",x"3a84",x"b81e",x"3444",x"364c",x"31d5",x"b966",x"4053",x"3752",x"3a92",x"b7fc",x"346c",x"365c",x"3204"),
(x"b963",x"405d",x"3780",x"3bd2",x"3047",x"b134",x"35a0",x"1f3a",x"b964",x"4057",x"377a",x"3b82",x"286a",x"b57a",x"35aa",x"214e",x"b961",x"405a",x"378b",x"3bd2",x"3047",x"b133",x"35aa",x"2000"),
(x"b963",x"405d",x"3780",x"366b",x"ad14",x"3b4c",x"362f",x"31bd",x"b95b",x"405c",x"3777",x"3827",x"3037",x"3ac1",x"3628",x"31c1",x"b959",x"405b",x"3775",x"366b",x"ad14",x"3b4c",x"3626",x"31c9"),
(x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b",x"b963",x"405d",x"3780",x"2de3",x"3bd5",x"31ce",x"3658",x"2b68",x"b963",x"405b",x"3797",x"3553",x"3a2a",x"3858",x"3650",x"2b30"),
(x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b",x"b975",x"405a",x"37b0",x"1fc8",x"3964",x"39e8",x"3641",x"2b5a",x"b98a",x"405b",x"379b",x"b5ee",x"392f",x"3951",x"363c",x"2bdc"),
(x"b986",x"405d",x"375d",x"28bc",x"3bf3",x"2e92",x"3652",x"2c29",x"b963",x"405d",x"3780",x"2de3",x"3bd5",x"31ce",x"3658",x"2b68",x"b97a",x"405d",x"37a0",x"10ea",x"3b79",x"35b5",x"3646",x"2b9b"),
(x"b95b",x"405d",x"3752",x"3410",x"3b92",x"3261",x"3669",x"2b9b",x"b952",x"405c",x"3752",x"38c8",x"39c1",x"35a4",x"366e",x"2b5b",x"b959",x"405b",x"3775",x"39b9",x"391a",x"348e",x"3661",x"2b30"),
(x"b981",x"405e",x"3752",x"24c2",x"3be9",x"30b5",x"3658",x"2c27",x"b95b",x"405d",x"3752",x"3410",x"3b92",x"3261",x"3669",x"2b9b",x"b963",x"405d",x"3780",x"2de3",x"3bd5",x"31ce",x"3658",x"2b68"),
(x"b9d3",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"b9e2",x"3f95",x"37cf",x"bafd",x"36b2",x"b3e9",x"3562",x"3530",x"b9f7",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518"),
(x"b9d3",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"b9e2",x"3f95",x"37cf",x"b33d",x"35ad",x"3b41",x"3604",x"30cf"),
(x"b981",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4",x"b970",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce",x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"b963",x"3f47",x"3752",x"0000",x"0000",x"3c00",x"35b6",x"2b4f",x"b96e",x"3f46",x"3752",x"330f",x"b68f",x"3b14",x"35af",x"2b2d",x"b95a",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88"),
(x"b970",x"3f95",x"37ce",x"373e",x"b495",x"3ac1",x"358b",x"2d70",x"b94a",x"3f58",x"3752",x"374a",x"b488",x"3ac0",x"35c3",x"2c17",x"b985",x"3f77",x"37bd",x"367e",x"b50d",x"3adc",x"3585",x"2cb9"),
(x"b94a",x"3f58",x"3752",x"3b2b",x"3633",x"b2e4",x"35e5",x"2c0c",x"b970",x"3f95",x"37ce",x"3af6",x"36ac",x"b42c",x"359e",x"2d3c",x"b95d",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91"),
(x"b9ce",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"b9e7",x"3f46",x"3752",x"b179",x"b6cc",x"3b1c",x"350b",x"349a",x"b9f1",x"3f48",x"3752",x"b5a1",x"b590",x"3af3",x"3506",x"349f"),
(x"b9e2",x"3f95",x"37cf",x"ba59",x"b59a",x"37f3",x"353f",x"350c",x"b9ce",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"ba0b",x"3f58",x"3752",x"b6ba",x"b4d8",x"3ad7",x"34fb",x"34bd"),
(x"b9a7",x"3f4b",x"380b",x"3b6a",x"b5fa",x"a856",x"35e2",x"2e9e",x"b9a9",x"3f49",x"380d",x"3ac4",x"b843",x"a386",x"35e1",x"2e92",x"b9a6",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1"),
(x"b9a9",x"3f49",x"382e",x"b94c",x"b9fe",x"2025",x"3582",x"3498",x"b9a9",x"3f49",x"380d",x"ba6f",x"b8bf",x"a6fd",x"356a",x"3496",x"b9ad",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c"),
(x"b9a7",x"3f4b",x"380b",x"3b6a",x"b5fa",x"a856",x"35e2",x"2e9e",x"b9a6",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1",x"b985",x"3f77",x"37bd",x"3b7c",x"b5a3",x"a1ae",x"3602",x"2fb5"),
(x"b9a6",x"3f4b",x"382c",x"38c7",x"30be",x"3a4d",x"35d2",x"31ac",x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"b970",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce"),
(x"b9e2",x"3f95",x"37cf",x"ba59",x"b59a",x"37f3",x"353f",x"350c",x"b9ad",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c",x"b9ce",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd"),
(x"b9ad",x"3f4b",x"382c",x"b89c",x"310b",x"3a6a",x"35d7",x"31ad",x"b9e2",x"3f95",x"37cf",x"b33d",x"35ad",x"3b41",x"3604",x"30cf",x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad"),
(x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"b9a6",x"3f4b",x"382c",x"38c7",x"30be",x"3a4d",x"35d2",x"31ac",x"b9a9",x"3f49",x"382e",x"2467",x"b509",x"3b97",x"35d4",x"31b1"),
(x"b9ad",x"3f4b",x"382c",x"b89c",x"310b",x"3a6a",x"35d7",x"31ad",x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"b9a9",x"3f49",x"382e",x"2467",x"b509",x"3b97",x"35d4",x"31b1"),
(x"b9d3",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"b9a9",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"b981",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4",x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"b9a9",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1"),
(x"b9a9",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"b9d3",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"b9b6",x"3fa3",x"37a0",x"363d",x"3811",x"3a23",x"35e2",x"3096"),
(x"b9a9",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"b995",x"3fa2",x"379c",x"b829",x"38f7",x"38b1",x"35c6",x"3094",x"b981",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4"),
(x"b995",x"3fa2",x"379c",x"38d4",x"376b",x"b92f",x"35ad",x"2dca",x"b98b",x"3f82",x"3752",x"381e",x"3818",x"b980",x"35d8",x"2d45",x"b981",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a"),
(x"b9b6",x"3fa3",x"37a0",x"b70f",x"36eb",x"ba4a",x"3560",x"355b",x"b9d3",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"b9d2",x"3f71",x"3752",x"b43c",x"3773",x"bac1",x"3517",x"3533"),
(x"b9b2",x"407a",x"3802",x"b75e",x"39fd",x"37a1",x"34fe",x"334f",x"ba10",x"407a",x"3752",x"b75e",x"39fd",x"37a1",x"355f",x"334f",x"b9b2",x"4088",x"3752",x"b75e",x"39fd",x"37a1",x"352a",x"32d0"),
(x"b9b1",x"4072",x"37be",x"39fd",x"0000",x"394d",x"3625",x"2c04",x"b982",x"4072",x"3752",x"39fd",x"0000",x"394d",x"35ef",x"2c07",x"b9b1",x"405c",x"37be",x"39fd",x"0000",x"394d",x"3625",x"2d00"),
(x"b9b1",x"405c",x"37be",x"b9ee",x"068d",x"395e",x"3641",x"2d01",x"b9e2",x"405e",x"3752",x"b9ee",x"0a8d",x"395e",x"360a",x"2d16",x"b9b1",x"4072",x"37be",x"b9ee",x"0a8d",x"395e",x"3641",x"2dfd"),
(x"ba10",x"407a",x"3752",x"b7fd",x"b973",x"3847",x"3615",x"2aa4",x"b9b2",x"407a",x"3802",x"b837",x"b940",x"3851",x"35b4",x"2aa4",x"b9e2",x"4071",x"3752",x"b837",x"b940",x"3851",x"35fc",x"2bb2"),
(x"b955",x"407a",x"3752",x"380d",x"b969",x"3846",x"34fe",x"3480",x"b982",x"4072",x"3752",x"3854",x"b926",x"3853",x"3516",x"34a2",x"b9b2",x"407a",x"3802",x"3854",x"b926",x"3853",x"355f",x"3481"),
(x"b955",x"407a",x"3752",x"374c",x"3a02",x"37a3",x"3597",x"2c08",x"b9b2",x"407a",x"3802",x"374c",x"3a02",x"37a3",x"3537",x"2c1c",x"b9b2",x"4088",x"3752",x"374c",x"3a02",x"37a3",x"3566",x"2d0f"),
(x"b9e7",x"3dc2",x"3752",x"baa2",x"935f",x"3878",x"34ae",x"3122",x"b9e8",x"3f49",x"3754",x"bab7",x"9f2b",x"3858",x"34ae",x"259c",x"b9aa",x"3dc3",x"3804",x"bab6",x"9af6",x"385a",x"345b",x"311f"),
(x"b9a9",x"3f4b",x"380f",x"3ad7",x"a303",x"3824",x"3507",x"2563",x"b96c",x"3f46",x"3755",x"3abd",x"9ffc",x"384e",x"34af",x"25db",x"b9aa",x"3dc3",x"3804",x"3abc",x"9c9b",x"3850",x"3507",x"311e"),
(x"b9a9",x"3f4b",x"380f",x"3ad7",x"a303",x"3824",x"3507",x"2563",x"b985",x"3f7c",x"37bc",x"3ad1",x"ab2e",x"3828",x"34d9",x"1b5d",x"b96c",x"3f46",x"3755",x"3abd",x"9ffc",x"384e",x"34af",x"25db"),
(x"b9a9",x"3f4b",x"380f",x"bac7",x"a224",x"383e",x"3455",x"2566",x"b9e8",x"3f49",x"3754",x"bab7",x"9f2b",x"3858",x"34ae",x"259c",x"b9cf",x"3f7c",x"37bb",x"bac2",x"abcb",x"383f",x"3483",x"1b5d"),
(x"b9a9",x"3db1",x"3832",x"b904",x"38e5",x"37b5",x"350c",x"3524",x"ba0f",x"3db3",x"3752",x"b8d1",x"395c",x"36f1",x"348c",x"3524",x"b9aa",x"3dc3",x"3804",x"b8d1",x"395c",x"36f1",x"34f0",x"3544"),
(x"b9a9",x"3db1",x"3832",x"38f7",x"3907",x"377c",x"3477",x"3500",x"b9aa",x"3dc3",x"3804",x"38d0",x"395f",x"36e9",x"3493",x"3520",x"b945",x"3db3",x"3752",x"38d0",x"395f",x"36e9",x"34f7",x"3500"),
(x"b9a9",x"3d16",x"3834",x"ba6e",x"1cd0",x"38c1",x"358f",x"1ca0",x"ba10",x"3d4c",x"3752",x"ba6d",x"1c32",x"38c3",x"3512",x"263e",x"b9a9",x"3db1",x"3832",x"ba6c",x"1b93",x"38c3",x"358f",x"2bd9"),
(x"b9a9",x"3d16",x"3834",x"3a6b",x"191e",x"38c5",x"3587",x"3495",x"b9a9",x"3db1",x"3832",x"3a6f",x"1d6d",x"38c0",x"3587",x"3369",x"b942",x"3d4d",x"3752",x"3a6f",x"1d6d",x"38c0",x"3505",x"3446"),
(x"b9a9",x"3d16",x"3834",x"1c67",x"3a22",x"3922",x"35eb",x"26d8",x"ba0d",x"3cfb",x"3871",x"a581",x"3a1a",x"392b",x"359d",x"2239",x"ba10",x"3d4c",x"3752",x"a8f7",x"3a35",x"3909",x"359e",x"2b69"),
(x"b946",x"3cfa",x"3872",x"27ce",x"3a15",x"3930",x"3638",x"221d",x"b9a9",x"3d16",x"3834",x"1c67",x"3a22",x"3922",x"35eb",x"26d8",x"b942",x"3d4d",x"3752",x"29e6",x"3a2c",x"3912",x"3638",x"2b6a"),
(x"b9a9",x"3d16",x"3834",x"1c67",x"3a22",x"3922",x"35eb",x"26d8",x"b946",x"3cfa",x"3872",x"27ce",x"3a15",x"3930",x"3638",x"221d",x"ba0d",x"3cfb",x"3871",x"a581",x"3a1a",x"392b",x"359d",x"2239"),
(x"ba11",x"3ca2",x"3752",x"bbff",x"1b5f",x"2393",x"3514",x"323a",x"ba10",x"3d4c",x"3752",x"bbff",x"1b5f",x"2393",x"3514",x"304b",x"ba0d",x"3cfb",x"3871",x"bbff",x"1b5f",x"2393",x"35aa",x"3137"),
(x"ba0d",x"3cfb",x"3871",x"9ef6",x"b9f8",x"3952",x"345f",x"34f8",x"b946",x"3cfa",x"3872",x"9b5f",x"b9fc",x"394f",x"34fa",x"34f8",x"ba11",x"3ca2",x"3752",x"9ac2",x"b9fc",x"394e",x"345f",x"3435"),
(x"b946",x"3cfa",x"3872",x"3bff",x"928d",x"2425",x"350a",x"301f",x"b942",x"3d4d",x"3752",x"3bff",x"928d",x"2425",x"35a1",x"310e",x"b943",x"3ca2",x"3752",x"3bff",x"928d",x"2425",x"35a1",x"2e3b"),
(x"ba10",x"30ed",x"3752",x"bc00",x"168d",x"9a24",x"350e",x"2c14",x"ba0f",x"3520",x"3752",x"bc00",x"168d",x"9a24",x"350d",x"2ff1",x"ba10",x"3396",x"3874",x"bc00",x"168d",x"9a24",x"35a6",x"2e06"),
(x"ba0f",x"3520",x"3752",x"205a",x"3a22",x"3922",x"3460",x"32b2",x"b943",x"351b",x"3752",x"0e8d",x"3a2a",x"3918",x"34fa",x"32b2",x"ba10",x"3396",x"3874",x"0e8d",x"3a2a",x"3918",x"3461",x"3131"),
(x"ba10",x"30ed",x"3752",x"191e",x"ba22",x"3922",x"3464",x"32c1",x"ba10",x"3396",x"3874",x"96f6",x"ba26",x"391d",x"3465",x"3428",x"b943",x"30ef",x"3752",x"9624",x"ba26",x"391d",x"34f9",x"32bf"),
(x"b945",x"3397",x"3877",x"3c00",x"11bc",x"205a",x"34ff",x"3271",x"b943",x"351b",x"3752",x"3c00",x"11bc",x"205a",x"3593",x"317b",x"b943",x"30ef",x"3752",x"3c00",x"11bc",x"205a",x"359b",x"336c"),
(x"b9f8",x"4024",x"378d",x"ba5b",x"36b9",x"3703",x"3622",x"3459",x"b9ff",x"401f",x"3786",x"baf9",x"ae2b",x"37ae",x"3620",x"344a",x"ba05",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"360a",x"345b"),
(x"b9f2",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3624",x"3460",x"b9f8",x"4024",x"378d",x"ba5b",x"36b9",x"3703",x"3622",x"3459",x"b9fc",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"360c",x"3464"),
(x"b9e7",x"4027",x"378f",x"2731",x"3bb3",x"3450",x"3628",x"3467",x"b9f2",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3624",x"3460",x"b9f4",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"360e",x"346a"),
(x"b9f0",x"400d",x"3777",x"bb0c",x"b28a",x"36d3",x"362a",x"3414",x"b9f8",x"400d",x"3752",x"bae9",x"b336",x"3733",x"361b",x"3412",x"b9ff",x"401f",x"3786",x"baf9",x"ae2b",x"37ae",x"3620",x"344a"),
(x"b9e8",x"4002",x"376d",x"baf0",x"b0d8",x"3796",x"362f",x"33e9",x"b9f0",x"4002",x"3752",x"bb07",x"b070",x"374f",x"3623",x"33e8",x"b9f0",x"400d",x"3777",x"bb0c",x"b28a",x"36d3",x"362a",x"3414"),
(x"b9e7",x"4027",x"378f",x"2731",x"3bb3",x"3450",x"3628",x"3467",x"b9f4",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"360e",x"346a",x"b9dc",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"362c",x"346e"),
(x"b9d3",x"4023",x"378c",x"3949",x"390d",x"367c",x"3632",x"3477",x"b9dc",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"362c",x"346e",x"b9d5",x"4024",x"3782",x"3904",x"3a39",x"a8ac",x"362c",x"3476"),
(x"b9e8",x"4002",x"376d",x"afac",x"ad49",x"3bea",x"357c",x"34d1",x"b9f0",x"400d",x"3777",x"9d6d",x"aedf",x"3bf4",x"3578",x"34f2",x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"b9ff",x"401f",x"3786",x"b0fd",x"b014",x"3bd6",x"356f",x"3528",x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9f0",x"400d",x"3777",x"9d6d",x"aedf",x"3bf4",x"3578",x"34f2"),
(x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9f8",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3575",x"3536"),
(x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9f2",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"357a",x"353b"),
(x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9e7",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3582",x"353d"),
(x"b9e0",x"4025",x"378f",x"b17c",x"b4ab",x"3b87",x"3587",x"3537",x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9dc",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"b9d3",x"4023",x"378c",x"287a",x"ad2b",x"3bf8",x"3591",x"3531",x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9dc",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9cf",x"4022",x"378b",x"2ef6",x"b0cc",x"3bdc",x"3594",x"352f",x"b9d7",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"358e",x"3523"),
(x"b9cf",x"4017",x"377f",x"27d5",x"aef0",x"3bf2",x"3593",x"350f",x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9ce",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"b9cf",x"400d",x"3777",x"abbe",x"ace8",x"3bf6",x"3591",x"34f1",x"b9d7",x"400e",x"3777",x"ac2d",x"ae61",x"3bf1",x"358b",x"34f3",x"b9cf",x"4017",x"377f",x"27d5",x"aef0",x"3bf2",x"3593",x"350f"),
(x"b9cd",x"3fff",x"3770",x"ae76",x"a942",x"3bf3",x"3590",x"34c9",x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9cf",x"400d",x"3777",x"abbe",x"ace8",x"3bf6",x"3591",x"34f1"),
(x"b9dc",x"400e",x"3775",x"b232",x"ad32",x"3bd2",x"3587",x"34f5",x"b9d7",x"400e",x"3777",x"ac2d",x"ae61",x"3bf1",x"358b",x"34f3",x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2"),
(x"b9df",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3586",x"3512",x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9dc",x"400e",x"3775",x"b232",x"ad32",x"3bd2",x"3587",x"34f5"),
(x"b9d7",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"358e",x"3523",x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523"),
(x"b9dd",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3589",x"352f",x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523"),
(x"b9e0",x"4025",x"378f",x"b17c",x"b4ab",x"3b87",x"3587",x"3537",x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534"),
(x"b9e7",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3581",x"3535",x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534"),
(x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534",x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9e7",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3581",x"3535"),
(x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531",x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534"),
(x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527",x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3",x"b9e8",x"400d",x"3776",x"349f",x"a9d6",x"3ba6",x"357d",x"34f3",x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527"),
(x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"b9e8",x"400d",x"3776",x"349f",x"a9d6",x"3ba6",x"357d",x"34f3",x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"b9dc",x"400e",x"3775",x"b232",x"ad32",x"3bd2",x"3587",x"34f5",x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527",x"b9df",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3586",x"3512",x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523",x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527"),
(x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534",x"b9dd",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3589",x"352f",x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"b9e7",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3581",x"3535",x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534",x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534"),
(x"b9cb",x"400d",x"378a",x"bbec",x"2694",x"3049",x"3648",x"317b",x"b9cd",x"3fff",x"3770",x"bbe8",x"9e0a",x"30d2",x"3648",x"31cd",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b"),
(x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140",x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b"),
(x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a",x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b",x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140"),
(x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102",x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108",x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a"),
(x"b9cd",x"4024",x"37aa",x"ba49",x"b805",x"35c1",x"364a",x"30f4",x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff",x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee",x"b9c6",x"4023",x"37b6",x"b9d1",x"b94b",x"31cf",x"3644",x"30fb",x"b9cd",x"4024",x"37aa",x"ba49",x"b805",x"35c1",x"364a",x"30f4"),
(x"b9cd",x"4023",x"37c8",x"bb6a",x"b4dc",x"b301",x"363e",x"30f1",x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112"),
(x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133"),
(x"b9ca",x"400d",x"379f",x"bbf8",x"2d3a",x"a850",x"3640",x"3175",x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"b9cd",x"3fff",x"3790",x"bbfe",x"2874",x"9fc8",x"363d",x"31c9",x"b9ca",x"400d",x"379f",x"bbf8",x"2d3a",x"a850",x"3640",x"3175",x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"b9cd",x"3fff",x"3790",x"bbfe",x"2874",x"9fc8",x"363d",x"31c9",x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174",x"b9cc",x"3fff",x"3798",x"bbe2",x"a7a0",x"314e",x"363a",x"31c7"),
(x"b9cc",x"4017",x"37d1",x"bbf6",x"a89b",x"2d9b",x"3632",x"3134",x"b9cb",x"400d",x"37b2",x"bbee",x"a8fd",x"2fea",x"3638",x"3174",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133"),
(x"b9cc",x"401d",x"37de",x"bbe7",x"9e8d",x"30f2",x"3631",x"3110",x"b9cc",x"4017",x"37d1",x"bbf6",x"a89b",x"2d9b",x"3632",x"3134",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112"),
(x"b9cc",x"4022",x"37dc",x"bbdb",x"2a31",x"31d8",x"3635",x"30f7",x"b9cc",x"401d",x"37de",x"bbe7",x"9e8d",x"30f2",x"3631",x"3110",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"b9cc",x"4024",x"37cc",x"bbf1",x"2b1a",x"2ec3",x"363d",x"30ea",x"b9cc",x"4022",x"37dc",x"bbdb",x"2a31",x"31d8",x"3635",x"30f7",x"b9cd",x"4023",x"37c8",x"bb6a",x"b4dc",x"b301",x"363e",x"30f1"),
(x"b9cd",x"4025",x"37b8",x"bbfc",x"2752",x"2a48",x"3645",x"30e8",x"b9cc",x"4024",x"37cc",x"bbf1",x"2b1a",x"2ec3",x"363d",x"30ea",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9cd",x"4024",x"37aa",x"ba49",x"b805",x"35c1",x"364a",x"30f4",x"b9cd",x"4025",x"37a7",x"bbff",x"21bc",x"2518",x"364c",x"30ed",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9ce",x"4022",x"378e",x"bbf3",x"a2c2",x"2ede",x"3654",x"3100",x"b9cd",x"4025",x"37a7",x"bbff",x"21bc",x"2518",x"364c",x"30ed",x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"b9cf",x"4022",x"378b",x"bafb",x"aeae",x"37a0",x"3656",x"3100",x"b9ce",x"4022",x"378e",x"bbf3",x"a2c2",x"2ede",x"3654",x"3100",x"b9ce",x"401e",x"3784",x"bbd5",x"a432",x"3276",x"3656",x"311b"),
(x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102",x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a",x"b9ce",x"4022",x"378e",x"bbf3",x"a2c2",x"2ede",x"3654",x"3100"),
(x"b9cf",x"4017",x"377f",x"bbc6",x"a57a",x"337e",x"3654",x"3142",x"b9ce",x"401e",x"3784",x"bbd5",x"a432",x"3276",x"3656",x"311b",x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140"),
(x"b9cf",x"400d",x"3777",x"bbc7",x"a88b",x"3365",x"364f",x"317c",x"b9cf",x"4017",x"377f",x"bbc6",x"a57a",x"337e",x"3654",x"3142",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b"),
(x"b9cf",x"400d",x"3777",x"bbc7",x"a88b",x"3365",x"364f",x"317c",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b",x"b9cd",x"3fff",x"3770",x"bbe8",x"9e0a",x"30d2",x"3648",x"31cd"),
(x"b9cd",x"3fff",x"3770",x"bbe8",x"9e0a",x"30d2",x"3648",x"31cd",x"b9cb",x"400d",x"378a",x"bbec",x"2694",x"3049",x"3648",x"317b",x"b9cd",x"3fff",x"3790",x"bbfe",x"2874",x"9fc8",x"363d",x"31c9"),
(x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9ca",x"400d",x"379f",x"bbf8",x"2d3a",x"a850",x"3640",x"3175",x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f"),
(x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b"),
(x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108"),
(x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff"),
(x"b9c6",x"4023",x"37b6",x"b9d1",x"b94b",x"31cf",x"3644",x"30fb",x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff"),
(x"b9cc",x"3fff",x"3798",x"b864",x"b1fa",x"3a84",x"35df",x"341e",x"b9cb",x"400d",x"37b2",x"b866",x"b31b",x"3a70",x"35df",x"33e6",x"b9ae",x"3ffe",x"37c0",x"2418",x"b372",x"3bc7",x"35c2",x"341c"),
(x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b9cc",x"4017",x"37d1",x"b86f",x"b4aa",x"3a3c",x"35de",x"33a2"),
(x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b9cc",x"401d",x"37de",x"b896",x"af43",x"3a7d",x"35db",x"337c"),
(x"b9ac",x"4024",x"37fd",x"23bb",x"3849",x"3ac0",x"35c1",x"3362",x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b9cc",x"4022",x"37dc",x"b830",x"3619",x"3a17",x"35d9",x"3360"),
(x"b9cc",x"4024",x"37cc",x"b5be",x"3a7e",x"375e",x"35d9",x"334c",x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351",x"b9cc",x"4022",x"37dc",x"b830",x"3619",x"3a17",x"35d9",x"3360"),
(x"b9cd",x"4025",x"37b8",x"b483",x"3bab",x"291b",x"35da",x"333c",x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341",x"b9cc",x"4024",x"37cc",x"b5be",x"3a7e",x"375e",x"35d9",x"334c"),
(x"b9cd",x"4025",x"37a7",x"b469",x"3b1b",x"b5df",x"35db",x"332f",x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331",x"b9cd",x"4025",x"37b8",x"b483",x"3bab",x"291b",x"35da",x"333c"),
(x"b9ce",x"4022",x"378e",x"b717",x"3a25",x"b764",x"35e0",x"3319",x"b9c4",x"4025",x"379c",x"b51a",x"3ab3",x"b716",x"35d5",x"3325",x"b9cd",x"4025",x"37a7",x"b469",x"3b1b",x"b5df",x"35db",x"332f"),
(x"b9ca",x"4023",x"378b",x"b8bf",x"3a5d",x"afac",x"35dc",x"3317",x"b9c4",x"4025",x"379c",x"b51a",x"3ab3",x"b716",x"35d5",x"3325",x"b9ce",x"4022",x"378e",x"b717",x"3a25",x"b764",x"35e0",x"3319"),
(x"b9cf",x"4022",x"378b",x"3842",x"3832",x"3950",x"3633",x"347b",x"b9d3",x"4023",x"378c",x"3949",x"390d",x"367c",x"3632",x"3477",x"b9cd",x"4022",x"3786",x"3818",x"3947",x"3865",x"3631",x"347c"),
(x"b9cf",x"4022",x"378b",x"b80a",x"3a5a",x"3567",x"35e0",x"3316",x"b9cd",x"4022",x"3786",x"b6e0",x"3aa3",x"35b0",x"35df",x"3313",x"b9ce",x"4022",x"378e",x"b718",x"3a24",x"b765",x"35e0",x"3319"),
(x"b94b",x"4020",x"3752",x"3acd",x"aeb3",x"381f",x"363b",x"3478",x"b95b",x"401f",x"3786",x"3ae5",x"ae76",x"37f1",x"3652",x"3477",x"b956",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"363c",x"3466"),
(x"b956",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"363c",x"3466",x"b962",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3655",x"3468",x"b95e",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"363e",x"345e"),
(x"b95e",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"363e",x"345e",x"b968",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3656",x"3461",x"b966",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"3640",x"3458"),
(x"b96c",x"400d",x"3775",x"3abf",x"b1e9",x"3808",x"365d",x"34ae",x"b95b",x"401f",x"3786",x"3ae5",x"ae76",x"37f1",x"3652",x"3477",x"b962",x"400d",x"3752",x"3aca",x"b303",x"37b2",x"364e",x"34af"),
(x"b972",x"4001",x"376d",x"3a5f",x"af27",x"38c0",x"3663",x"34cf",x"b96c",x"400d",x"3775",x"3abf",x"b1e9",x"3808",x"365d",x"34ae",x"b967",x"4002",x"3752",x"3ab1",x"af0f",x"3849",x"3656",x"34ce"),
(x"b966",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"3640",x"3458",x"b973",x"4027",x"378f",x"a731",x"3bb3",x"3450",x"365a",x"345a",x"b97e",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"365e",x"3453"),
(x"b987",x"4023",x"378c",x"b932",x"391d",x"3694",x"3664",x"344a",x"b985",x"4024",x"3782",x"b907",x"3a38",x"a54c",x"365e",x"344b",x"b97e",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"365e",x"3453"),
(x"b972",x"4001",x"376d",x"303c",x"aa80",x"3beb",x"3641",x"30bf",x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0",x"b96c",x"400d",x"3775",x"2b97",x"ae90",x"3bf1",x"3642",x"307d"),
(x"b96c",x"400d",x"3775",x"2b97",x"ae90",x"3bf1",x"3642",x"307d",x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079",x"b95b",x"401f",x"3786",x"2e5c",x"b067",x"3be2",x"363e",x"300d"),
(x"b95b",x"401f",x"3786",x"2e5c",x"b067",x"3be2",x"363e",x"300d",x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e",x"b962",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3645",x"2fe4"),
(x"b962",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3645",x"2fe4",x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee",x"b968",x"4026",x"378e",x"2d5c",x"a067",x"3bf8",x"364b",x"2fd2"),
(x"b968",x"4026",x"378e",x"2d5c",x"a067",x"3bf8",x"364b",x"2fd2",x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf",x"b973",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3653",x"2fce"),
(x"b973",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3653",x"2fce",x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd",x"b97e",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"365b",x"2fdd"),
(x"b987",x"4023",x"378c",x"a87a",x"ad2b",x"3bf8",x"3661",x"3001",x"b97e",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"365b",x"2fdd",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003"),
(x"b983",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"365c",x"301d",x"b98c",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3664",x"3007",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003"),
(x"b98b",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"365f",x"3047",x"b98c",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3662",x"3020",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040"),
(x"b98c",x"400d",x"3777",x"296a",x"ace7",x"3bf8",x"365a",x"3081",x"b98b",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"365f",x"3047",x"b983",x"400e",x"3777",x"2c32",x"ae3d",x"3bf1",x"3654",x"307b"),
(x"b98d",x"4000",x"3770",x"2c3e",x"a8a5",x"3bfa",x"3655",x"30cc",x"b98c",x"400d",x"3777",x"296a",x"ace7",x"3bf8",x"365a",x"3081",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"b983",x"400e",x"3777",x"2c32",x"ae3d",x"3bf1",x"3654",x"307b",x"b97e",x"400e",x"3775",x"3224",x"ad11",x"3bd3",x"3651",x"3077",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"b97b",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3653",x"303e",x"b97e",x"400e",x"3775",x"3224",x"ad11",x"3bd3",x"3651",x"3077",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040"),
(x"b97b",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3653",x"303e",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b"),
(x"b97d",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3658",x"3004",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003"),
(x"b97d",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3658",x"3004",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003",x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"b973",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5",x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd"),
(x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b973",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf"),
(x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee"),
(x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e"),
(x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079",x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079"),
(x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079",x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0",x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079"),
(x"b97e",x"400e",x"3775",x"3224",x"ad11",x"3bd3",x"3651",x"3077",x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079",x"b97b",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3653",x"303e"),
(x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b"),
(x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b97d",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3658",x"3004"),
(x"b973",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"b98d",x"4000",x"3770",x"3be7",x"a0ea",x"30f9",x"3661",x"2df3",x"b98f",x"400d",x"378a",x"3bdf",x"2581",x"319c",x"365f",x"2e8f",x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f"),
(x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03",x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50",x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03",x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f",x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50",x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74"),
(x"b98d",x"4024",x"37aa",x"3a75",x"b7d2",x"354a",x"3662",x"2f9c",x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89"),
(x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7",x"b98d",x"4024",x"37aa",x"3a75",x"b7d2",x"354a",x"3662",x"2f9c",x"b993",x"4023",x"37b7",x"39e1",x"b96b",x"23fc",x"365c",x"2f93"),
(x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7",x"b993",x"4023",x"37b7",x"39e1",x"b96b",x"23fc",x"365c",x"2f93",x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4",x"b993",x"4022",x"37c3",x"3af0",x"b4e6",x"b647",x"3658",x"2f91",x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c"),
(x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c",x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61",x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e",x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b98e",x"400d",x"37a5",x"3b77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b98f",x"3ffd",x"378d",x"3bfd",x"9d53",x"29ab",x"3655",x"2de8",x"b98e",x"400d",x"37a5",x"3b77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"b990",x"3ffd",x"3797",x"3be2",x"ab03",x"3119",x"3651",x"2de7",x"b98e",x"400d",x"37b0",x"3bfb",x"a724",x"2bb7",x"3651",x"2e9c",x"b98f",x"3ffd",x"378d",x"3bfd",x"9d53",x"29ab",x"3655",x"2de8"),
(x"b98e",x"400d",x"37a5",x"3b77",x"2f4d",x"b571",x"3655",x"2e9c",x"b98e",x"400d",x"37b0",x"3bfb",x"a724",x"2bb7",x"3651",x"2e9c",x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e",x"b98e",x"4017",x"37d0",x"3c00",x"9e59",x"868d",x"364a",x"2f1c",x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61",x"b98e",x"401d",x"37dc",x"3bfd",x"135f",x"a9d9",x"364a",x"2f66",x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c"),
(x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c",x"b98e",x"4022",x"37db",x"3bff",x"1b2b",x"2560",x"364e",x"2f95",x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4",x"b98e",x"4024",x"37cd",x"3bf5",x"2bb1",x"2d1b",x"3655",x"2fb0",x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7"),
(x"b98d",x"4024",x"37aa",x"3a75",x"b7d2",x"354a",x"3662",x"2f9c",x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7",x"b98d",x"4025",x"37a7",x"3bff",x"1fc8",x"25fd",x"3664",x"2fa8"),
(x"b98d",x"4024",x"37aa",x"3a75",x"b7d2",x"354a",x"3662",x"2f9c",x"b98d",x"4025",x"37a7",x"3bff",x"1fc8",x"25fd",x"3664",x"2fa8",x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f"),
(x"b98d",x"4022",x"378e",x"3bf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"b98c",x"4022",x"378b",x"3afb",x"aeb0",x"37a0",x"366e",x"2f82",x"b98c",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"366e",x"2f4e"),
(x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f",x"b98d",x"4022",x"378e",x"3bf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50"),
(x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50",x"b98c",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"366e",x"2f4e",x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03"),
(x"b98c",x"400d",x"3777",x"3bc5",x"a8b2",x"3387",x"3667",x"2e8b",x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"b98b",x"4017",x"377f",x"3bc6",x"a57a",x"3387",x"366c",x"2f00"),
(x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"b98c",x"400d",x"3777",x"3bc5",x"a8b2",x"3387",x"3667",x"2e8b",x"b98d",x"4000",x"3770",x"3be7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"b98f",x"3ffd",x"378d",x"3bfd",x"9d53",x"29ab",x"3655",x"2de8",x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b98d",x"4000",x"3770",x"3be7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"b98f",x"400d",x"378a",x"3bdf",x"2581",x"319c",x"365f",x"2e8f",x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05",x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e",x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74"),
(x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74",x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89"),
(x"b993",x"4022",x"37c3",x"3af0",x"b4e6",x"b647",x"3658",x"2f91",x"b993",x"4023",x"37b7",x"39e1",x"b96b",x"23fc",x"365c",x"2f93",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89"),
(x"b990",x"3ffd",x"3797",x"3851",x"b1da",x"3a92",x"35a6",x"3422",x"b9ae",x"3ffe",x"37c0",x"2418",x"b372",x"3bc7",x"35c2",x"341c",x"b98e",x"400d",x"37b0",x"3883",x"b339",x"3a5a",x"35a4",x"33e7"),
(x"b98e",x"400d",x"37b0",x"3883",x"b339",x"3a5a",x"35a4",x"33e7",x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b98e",x"4017",x"37d0",x"3883",x"b46b",x"3a39",x"35a5",x"33a3"),
(x"b98e",x"4017",x"37d0",x"3883",x"b46b",x"3a39",x"35a5",x"33a3",x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b98e",x"401d",x"37dc",x"388e",x"afce",x"3a80",x"35a7",x"337c"),
(x"b98e",x"401d",x"37dc",x"388e",x"afce",x"3a80",x"35a7",x"337c",x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b98e",x"4022",x"37db",x"3859",x"3581",x"3a1f",x"35a9",x"3362"),
(x"b98e",x"4024",x"37cd",x"3609",x"3a62",x"3783",x"35aa",x"334e",x"b98e",x"4022",x"37db",x"3859",x"3581",x"3a1f",x"35a9",x"3362",x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351"),
(x"b98d",x"4025",x"37b8",x"34be",x"3ba1",x"2a04",x"35a8",x"333e",x"b98e",x"4024",x"37cd",x"3609",x"3a62",x"3783",x"35aa",x"334e",x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341"),
(x"b98d",x"4025",x"37a7",x"34f8",x"3b04",x"b5db",x"35a6",x"3332",x"b98d",x"4025",x"37b8",x"34be",x"3ba1",x"2a04",x"35a8",x"333e",x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331"),
(x"b98d",x"4022",x"378e",x"38e6",x"391d",x"b76f",x"35a1",x"331c",x"b98d",x"4025",x"37a7",x"34f8",x"3b04",x"b5db",x"35a6",x"3332",x"b995",x"4024",x"3789",x"3533",x"3ac8",x"b6b3",x"35a9",x"3318"),
(x"b995",x"4024",x"3789",x"3533",x"3ac8",x"b6b3",x"35a9",x"3318",x"b990",x"4023",x"378b",x"37bd",x"3afd",x"2a63",x"35a4",x"331a",x"b98d",x"4022",x"378e",x"38e6",x"391d",x"b76f",x"35a1",x"331c"),
(x"b98c",x"4022",x"378b",x"b889",x"38bf",x"3891",x"3665",x"3446",x"b98e",x"4022",x"3782",x"b856",x"3952",x"381b",x"3662",x"3443",x"b987",x"4023",x"378c",x"b932",x"391d",x"3695",x"3664",x"344a"),
(x"b98d",x"4022",x"378e",x"38e6",x"391d",x"b76f",x"35a1",x"331c",x"b990",x"4023",x"378b",x"37bd",x"3afd",x"2a63",x"35a4",x"331a",x"b98c",x"4022",x"378b",x"371a",x"3b19",x"2ff2",x"35a0",x"3319"),
(x"b972",x"4001",x"376d",x"3a5f",x"af27",x"38c0",x"3663",x"34cf",x"b967",x"4002",x"3752",x"3ab1",x"af0f",x"3849",x"3656",x"34ce",x"b972",x"3ffb",x"376e",x"3ab9",x"ac8e",x"384b",x"3665",x"34da"),
(x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0",x"b972",x"4001",x"376d",x"303c",x"aa80",x"3beb",x"3641",x"30bf",x"b97b",x"3fff",x"3770",x"2d3d",x"28c9",x"3bf7",x"3647",x"30ce"),
(x"b97b",x"3fff",x"3770",x"2d3d",x"28c9",x"3bf7",x"3647",x"30ce",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2",x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0"),
(x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2",x"b97b",x"3fff",x"3770",x"2d3d",x"28c9",x"3bf7",x"3647",x"30ce",x"b98d",x"4000",x"3770",x"2c3e",x"a8a5",x"3bfa",x"3655",x"30cc"),
(x"b9e8",x"4002",x"376d",x"baf0",x"b0d8",x"3796",x"362f",x"33e9",x"b9e6",x"3ff8",x"376e",x"bafe",x"ac6a",x"37b1",x"3633",x"33c7",x"b9f0",x"4002",x"3752",x"bb07",x"b070",x"374f",x"3623",x"33e8"),
(x"b9e6",x"3ff8",x"376e",x"ad21",x"068d",x"3bf9",x"357c",x"34c0",x"b9e8",x"4002",x"376d",x"afac",x"ad49",x"3bea",x"357c",x"34d1",x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"b9e6",x"3ff8",x"376e",x"ad21",x"068d",x"3bf9",x"357c",x"34c0",x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"b9d5",x"3ffc",x"3770",x"a935",x"1d6d",x"3bfe",x"3589",x"34c5"),
(x"b9d5",x"3ffc",x"3770",x"a935",x"1d6d",x"3bfe",x"3589",x"34c5",x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9cd",x"3fff",x"3770",x"ae76",x"a942",x"3bf3",x"3590",x"34c9"),
(x"b9f8",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"3613",x"34eb",x"b9ff",x"404b",x"3786",x"baf5",x"afa4",x"37a8",x"3610",x"34de",x"ba05",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35fb",x"34ec"),
(x"b9f2",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"3615",x"34f1",x"b9f8",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"3613",x"34eb",x"b9fc",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35fd",x"34f4"),
(x"b9e7",x"4051",x"378f",x"25dc",x"3bcd",x"330b",x"3619",x"34f8",x"b9f2",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"3615",x"34f1",x"b9f4",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35ff",x"34f9"),
(x"b9f0",x"403d",x"3777",x"baf8",x"b403",x"36bf",x"3619",x"34b3",x"b9f8",x"403d",x"3752",x"bad1",x"b46a",x"371a",x"360a",x"34b0",x"b9ff",x"404b",x"3786",x"baf5",x"afa4",x"37a8",x"3610",x"34de"),
(x"b9e8",x"4034",x"376d",x"bae5",x"b1fa",x"378a",x"361e",x"3499",x"b9f0",x"4034",x"3752",x"bafe",x"b17b",x"3746",x"3612",x"3497",x"b9f0",x"403d",x"3777",x"baf8",x"b403",x"36bf",x"3619",x"34b3"),
(x"b9e7",x"4051",x"378f",x"25dc",x"3bcd",x"330b",x"3619",x"34f8",x"b9f4",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35ff",x"34f9",x"b9dc",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"361c",x"34ff"),
(x"b9d3",x"404e",x"378c",x"38cb",x"39b0",x"35e1",x"3620",x"3508",x"b9dc",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"361c",x"34ff",x"b9d5",x"404f",x"3782",x"385b",x"3ab4",x"a80e",x"361b",x"3507"),
(x"b9f0",x"403d",x"3777",x"253f",x"b05f",x"3bec",x"3611",x"3305",x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9e8",x"4034",x"376d",x"a5e3",x"adbf",x"3bf7",x"360e",x"333a"),
(x"b9ff",x"404b",x"3786",x"b0f8",x"b10b",x"3bcd",x"3619",x"32ae",x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9f0",x"403d",x"3777",x"253f",x"b05f",x"3bec",x"3611",x"3305"),
(x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9f8",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3613",x"3297"),
(x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9f2",x"4051",x"378e",x"ad5b",x"a187",x"3bf8",x"360e",x"328f"),
(x"b9e6",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3605",x"3292",x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9e7",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"b9dc",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"35fe",x"3292",x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9e7",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"b9d3",x"404e",x"378c",x"2877",x"ae68",x"3bf4",x"35f7",x"32a1",x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9dc",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"35fe",x"3292"),
(x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9cf",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"35f4",x"32a5",x"b9d7",x"404a",x"3788",x"ac6f",x"b1f6",x"3bd7",x"35fb",x"32b8"),
(x"b9cf",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"35f6",x"32d9",x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9ce",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"b9cf",x"403d",x"3777",x"abbb",x"ae16",x"3bf2",x"35f8",x"3309",x"b9d7",x"403d",x"3777",x"ac2a",x"afe7",x"3beb",x"35fe",x"3305",x"b9cf",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"35f6",x"32d9"),
(x"b9cd",x"4032",x"3770",x"ae75",x"aa87",x"3bf2",x"35fa",x"334a",x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b",x"b9cf",x"403d",x"3777",x"abbb",x"ae16",x"3bf2",x"35f8",x"3309"),
(x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302",x"b9d7",x"403d",x"3777",x"ac2a",x"afe7",x"3beb",x"35fe",x"3305",x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b"),
(x"b9df",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3602",x"32d4",x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"b9d7",x"404a",x"3788",x"ac6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4",x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"b9e3",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3603",x"329c",x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4"),
(x"b9e7",x"4050",x"3787",x"2710",x"b98f",x"39bf",x"3606",x"329a",x"b9e6",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3605",x"3292",x"b9e3",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3603",x"329c"),
(x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b",x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9e7",x"4050",x"3787",x"2710",x"b98f",x"39bf",x"3606",x"329a"),
(x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1",x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b"),
(x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0",x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1"),
(x"b9e5",x"403d",x"3773",x"2db8",x"ad34",x"3bf1",x"3609",x"3304",x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9e5",x"403d",x"3773",x"2db8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b",x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0",x"b9df",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3602",x"32d4",x"b9e5",x"403d",x"3773",x"2db8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7",x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b",x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4",x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1"),
(x"b9e7",x"4050",x"3787",x"2710",x"b98f",x"39bf",x"3606",x"329a",x"b9e3",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3603",x"329c",x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b"),
(x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9cd",x"4032",x"3770",x"bbc5",x"a836",x"338d",x"35a6",x"34c4",x"b9cd",x"403d",x"3783",x"bb8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"b9c8",x"4045",x"3794",x"bbbc",x"287e",x"3408",x"35a6",x"348a",x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9cd",x"404a",x"3790",x"bb17",x"ade0",x"3741",x"35ac",x"347b",x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9c6",x"404d",x"37a3",x"bbd3",x"a9fd",x"3272",x"35a4",x"3474",x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9cd",x"404f",x"37aa",x"b9e5",x"b8ae",x"3566",x"35a5",x"346b",x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468",x"b9c6",x"404e",x"37b6",x"b93b",x"b9e8",x"313a",x"359f",x"346f",x"b9cd",x"404f",x"37aa",x"b9e5",x"b8ae",x"3566",x"35a5",x"346b"),
(x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469",x"b9c6",x"404e",x"37c1",x"ba55",x"b865",x"b441",x"359c",x"346e",x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468"),
(x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e",x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477"),
(x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485"),
(x"b9ca",x"403d",x"379f",x"bbf7",x"2d6b",x"a836",x"359d",x"34a0",x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f"),
(x"b9cb",x"4031",x"378d",x"bbfd",x"1418",x"2a73",x"359b",x"34c3",x"b9ca",x"403d",x"379f",x"bbf7",x"2d6b",x"a836",x"359d",x"34a0",x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f"),
(x"b9cb",x"4031",x"378d",x"bbfd",x"1418",x"2a73",x"359b",x"34c3",x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f",x"b9ca",x"4031",x"3795",x"bbe2",x"acf4",x"30cc",x"3598",x"34c3"),
(x"b9cc",x"4045",x"37d1",x"bbf6",x"a9b5",x"2d99",x"358e",x"3485",x"b9cb",x"403d",x"37b2",x"bbec",x"ac1f",x"2fcd",x"3595",x"349f",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485"),
(x"b9cc",x"404a",x"37de",x"bbe7",x"a00b",x"30f2",x"358d",x"3476",x"b9cc",x"4045",x"37d1",x"bbf6",x"a9b5",x"2d99",x"358e",x"3485",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477"),
(x"b9cc",x"404d",x"37dc",x"bbd6",x"2b52",x"322d",x"3590",x"346c",x"b9cc",x"404a",x"37de",x"bbe7",x"a00b",x"30f2",x"358d",x"3476",x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469",x"b9cc",x"4050",x"37cc",x"bbe3",x"2d8f",x"3091",x"3598",x"3466",x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468",x"b9cd",x"4050",x"37b8",x"bbf8",x"2c13",x"2b34",x"35a1",x"3466",x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"b9cd",x"404f",x"37aa",x"b9e5",x"b8ae",x"3566",x"35a5",x"346b",x"b9cd",x"4050",x"37a7",x"bbff",x"232b",x"2518",x"35a7",x"3469",x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468"),
(x"b9ce",x"404e",x"378e",x"bbf3",x"a432",x"2ede",x"35af",x"3471",x"b9cd",x"4050",x"37a7",x"bbff",x"232b",x"2518",x"35a7",x"3469",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9cf",x"404e",x"378b",x"baf6",x"b023",x"379a",x"35b1",x"3471",x"b9ce",x"404e",x"378e",x"bbf3",x"a432",x"2ede",x"35af",x"3471",x"b9ce",x"404a",x"3784",x"bbd5",x"a532",x"3276",x"35b1",x"347c"),
(x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472",x"b9cd",x"404a",x"3790",x"bb17",x"ade0",x"3741",x"35ac",x"347b",x"b9ce",x"404e",x"378e",x"bbf3",x"a432",x"2ede",x"35af",x"3471"),
(x"b9cf",x"4045",x"377f",x"bbc6",x"a6c8",x"337e",x"35b0",x"348c",x"b9ce",x"404a",x"3784",x"bbd5",x"a532",x"3276",x"35b1",x"347c",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9cf",x"403d",x"3777",x"bbc6",x"a9a5",x"3365",x"35ac",x"34a4",x"b9cf",x"4045",x"377f",x"bbc6",x"a6c8",x"337e",x"35b0",x"348c",x"b9cd",x"403d",x"3783",x"bb8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"b9cf",x"403d",x"3777",x"bbc6",x"a9a5",x"3365",x"35ac",x"34a4",x"b9cd",x"403d",x"3783",x"bb8f",x"ab5c",x"3527",x"35a7",x"34a3",x"b9cd",x"4032",x"3770",x"bbc5",x"a836",x"338d",x"35a6",x"34c4"),
(x"b9cd",x"4032",x"3770",x"bbc5",x"a836",x"338d",x"35a6",x"34c4",x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9cb",x"4031",x"378d",x"bbfd",x"1418",x"2a73",x"359b",x"34c3"),
(x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9ca",x"403d",x"379f",x"bbf7",x"2d6b",x"a836",x"359d",x"34a0",x"b9c8",x"4045",x"3794",x"bbbc",x"287e",x"3408",x"35a6",x"348a"),
(x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c"),
(x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9c6",x"404d",x"37a3",x"bbd3",x"a9fd",x"3272",x"35a4",x"3474"),
(x"b9c6",x"404e",x"37c1",x"ba55",x"b865",x"b441",x"359c",x"346e",x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470"),
(x"b9c6",x"404e",x"37b6",x"b93b",x"b9e8",x"313a",x"359f",x"346f",x"b9c6",x"404e",x"37c1",x"ba55",x"b865",x"b441",x"359c",x"346e",x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470"),
(x"b9ca",x"4031",x"3795",x"b89a",x"b412",x"3a37",x"3679",x"2ae7",x"b9cb",x"403d",x"37b2",x"b86e",x"b47a",x"3a45",x"367a",x"29b1",x"b9ae",x"4031",x"37c0",x"1bc8",x"b48d",x"3bab",x"365d",x"2ab9"),
(x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b9cc",x"4045",x"37d1",x"b856",x"b5aa",x"3a18",x"3678",x"28cc"),
(x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b9cc",x"404a",x"37de",x"b892",x"b07e",x"3a77",x"3675",x"284f"),
(x"b9ac",x"4050",x"37fd",x"232b",x"38f3",x"3a48",x"365b",x"2806",x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b9cc",x"404d",x"37dc",x"b809",x"374a",x"39de",x"3673",x"27ef"),
(x"b9cc",x"4050",x"37cc",x"b4ee",x"3aeb",x"3653",x"3673",x"275d",x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e",x"b9cc",x"404d",x"37dc",x"b809",x"374a",x"39de",x"3673",x"27ef"),
(x"b9cd",x"4050",x"37b8",x"b361",x"3bc7",x"282c",x"3674",x"26df",x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709",x"b9cc",x"4050",x"37cc",x"b4ee",x"3aeb",x"3653",x"3673",x"275d"),
(x"b9cd",x"4050",x"37a7",x"b362",x"3b62",x"b4ea",x"3676",x"2679",x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c",x"b9cd",x"4050",x"37b8",x"b361",x"3bc7",x"282c",x"3674",x"26df"),
(x"b9ce",x"404e",x"378e",x"b62d",x"3aa4",x"b670",x"3679",x"25cc",x"b9c4",x"4050",x"379c",x"b458",x"3b15",x"b609",x"366f",x"2623",x"b9cd",x"4050",x"37a7",x"b362",x"3b62",x"b4ea",x"3676",x"2679"),
(x"b9ca",x"404e",x"378b",x"b819",x"3ad2",x"aea1",x"3676",x"25ba",x"b9c4",x"4050",x"379c",x"b458",x"3b15",x"b609",x"366f",x"2623",x"b9ce",x"404e",x"378e",x"b62d",x"3aa4",x"b670",x"3679",x"25cc"),
(x"b9cf",x"404e",x"378b",x"37f4",x"38dc",x"38f4",x"3622",x"350b",x"b9d3",x"404e",x"378c",x"38cb",x"39b0",x"35e1",x"3620",x"3508",x"b9cd",x"404e",x"3786",x"375f",x"39e5",x"37e9",x"3620",x"350c"),
(x"b9cf",x"404e",x"378b",x"b6fc",x"3ace",x"34aa",x"367a",x"25b5",x"b9cd",x"404e",x"3786",x"b5dc",x"3b09",x"34dc",x"3679",x"2599",x"b9ce",x"404e",x"378e",x"b62c",x"3aa4",x"b66f",x"3679",x"25cc"),
(x"b94b",x"404c",x"3752",x"3ac8",x"b025",x"381c",x"35de",x"2dda",x"b95b",x"404b",x"3786",x"3ae1",x"b000",x"37eb",x"35f5",x"2dd3",x"b956",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35e0",x"2d9e"),
(x"b956",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35e0",x"2d9e",x"b962",x"404f",x"378d",x"3a12",x"37fa",x"36b2",x"35f8",x"2da1",x"b95e",x"4053",x"3752",x"3848",x"3a10",x"35f5",x"35e2",x"2d7f"),
(x"b95e",x"4053",x"3752",x"3848",x"3a10",x"35f5",x"35e2",x"2d7f",x"b968",x"4051",x"378e",x"3610",x"3adf",x"357f",x"35fa",x"2d8a",x"b966",x"4053",x"3752",x"af69",x"3bdc",x"30a3",x"35e4",x"2d68"),
(x"b96c",x"403c",x"3775",x"3ab0",x"b345",x"37fd",x"35ff",x"2e87",x"b95b",x"404b",x"3786",x"3ae1",x"b000",x"37eb",x"35f5",x"2dd3",x"b962",x"403d",x"3752",x"3ab4",x"b44c",x"3799",x"35f0",x"2e8e"),
(x"b972",x"4033",x"376d",x"3a5a",x"b06c",x"38bc",x"3604",x"2ef0",x"b96c",x"403c",x"3775",x"3ab0",x"b345",x"37fd",x"35ff",x"2e87",x"b967",x"4034",x"3752",x"3aac",x"b05e",x"3846",x"35f7",x"2ef0"),
(x"b966",x"4053",x"3752",x"af69",x"3bdc",x"30a3",x"35e4",x"2d68",x"b973",x"4051",x"378f",x"a5dc",x"3bcb",x"332e",x"35fe",x"2d6c",x"b97e",x"4051",x"378e",x"b6f1",x"3b35",x"205a",x"3601",x"2d50"),
(x"b987",x"404e",x"378c",x"b8b4",x"39be",x"35f4",x"3605",x"2d2d",x"b985",x"404f",x"3782",x"b861",x"3ab1",x"a386",x"3600",x"2d31",x"b97e",x"4051",x"378e",x"b6f1",x"3b35",x"205a",x"3601",x"2d50"),
(x"b972",x"4033",x"376d",x"303b",x"ac06",x"3be9",x"3668",x"2c64",x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b96c",x"403c",x"3775",x"2dad",x"b0c1",x"3be1",x"3667",x"2cd0"),
(x"b95b",x"404b",x"3786",x"30f0",x"b192",x"3bc7",x"366a",x"2d86",x"b96c",x"403c",x"3775",x"2dad",x"b0c1",x"3be1",x"3667",x"2cd0",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"b95b",x"404b",x"3786",x"30f0",x"b192",x"3bc7",x"366a",x"2d86",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83",x"b962",x"404f",x"378d",x"2f46",x"b03f",x"3be0",x"3663",x"2db2"),
(x"b962",x"404f",x"378d",x"2f46",x"b03f",x"3be0",x"3663",x"2db2",x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8",x"b968",x"4051",x"378e",x"2d5c",x"a17a",x"3bf8",x"365d",x"2dbf"),
(x"b968",x"4051",x"378e",x"2d5c",x"a17a",x"3bf8",x"365d",x"2dbf",x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4",x"b973",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3655",x"2dc0"),
(x"b97e",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"364d",x"2db2",x"b973",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3655",x"2dc0",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"b987",x"404e",x"378c",x"a877",x"ae68",x"3bf4",x"3647",x"2d91",x"b97e",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"364d",x"2db2",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"b983",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"364c",x"2d65",x"b98c",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"3645",x"2d87",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"b98b",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"364a",x"2d20",x"b98c",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"b98c",x"403d",x"3777",x"2a04",x"ae02",x"3bf4",x"364f",x"2cc3",x"b98b",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"364a",x"2d20",x"b983",x"403d",x"3777",x"2c2f",x"afb9",x"3bec",x"3655",x"2cce"),
(x"b98d",x"4032",x"3770",x"2ca2",x"a97a",x"3bf8",x"3655",x"2c46",x"b98c",x"403d",x"3777",x"2a04",x"ae02",x"3bf4",x"364f",x"2cc3",x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"b983",x"403d",x"3777",x"2c2f",x"afb9",x"3bec",x"3655",x"2cce",x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"b97b",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3656",x"2d31",x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"b97b",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3656",x"2d31",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68"),
(x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"b977",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3654",x"2d9f",x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"b973",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3656",x"2da5",x"b977",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3654",x"2d9f",x"b975",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3654",x"2db4"),
(x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b973",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3656",x"2da5",x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4"),
(x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8"),
(x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"b975",x"403d",x"3773",x"adae",x"ad20",x"3bf1",x"3660",x"2cd4",x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b972",x"403d",x"3776",x"b31e",x"aca2",x"3bc7",x"3662",x"2cd4"),
(x"b972",x"403d",x"3776",x"b31e",x"aca2",x"3bc7",x"3662",x"2cd4",x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b975",x"403d",x"3773",x"adae",x"ad20",x"3bf1",x"3660",x"2cd4"),
(x"b975",x"403d",x"3773",x"adae",x"ad20",x"3bf1",x"3660",x"2cd4",x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5"),
(x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b975",x"403d",x"3773",x"adae",x"ad20",x"3bf1",x"3660",x"2cd4",x"b97b",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3656",x"2d31"),
(x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68"),
(x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d"),
(x"b973",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3656",x"2da5",x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b977",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3654",x"2d9f"),
(x"b98d",x"4032",x"3770",x"3be2",x"a025",x"3161",x"35f6",x"340d",x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8",x"b98d",x"403d",x"3782",x"3b88",x"abb1",x"354b",x"35f4",x"33d9"),
(x"b98d",x"403d",x"3782",x"3b88",x"abb1",x"354b",x"35f4",x"33d9",x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"b98d",x"404a",x"3790",x"3b10",x"ad8c",x"3760",x"35ed",x"338b",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa",x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b"),
(x"b98d",x"404a",x"3790",x"3b10",x"ad8c",x"3760",x"35ed",x"338b",x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b",x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"b98d",x"404f",x"37aa",x"3a13",x"b891",x"34fa",x"35f4",x"336a",x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b98d",x"404f",x"37aa",x"3a13",x"b891",x"34fa",x"35f4",x"336a",x"b993",x"404f",x"37b7",x"3977",x"b9c7",x"2ec0",x"35fa",x"336e"),
(x"b98d",x"404f",x"37c9",x"3b31",x"b5e3",x"b397",x"3600",x"3366",x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e"),
(x"b98d",x"404f",x"37c9",x"3b31",x"b5e3",x"b397",x"3600",x"3366",x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e",x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f",x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380",x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b"),
(x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b",x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1"),
(x"b990",x"403d",x"37a1",x"3bf5",x"2dc9",x"aa2b",x"3600",x"33d2",x"b98d",x"4030",x"378d",x"3bfe",x"28c2",x"2138",x"3602",x"340f",x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1"),
(x"b98e",x"403d",x"37b0",x"3bff",x"a3ef",x"2511",x"3606",x"33d1",x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1",x"b98e",x"4030",x"3797",x"3bf6",x"a3bb",x"2e0a",x"3606",x"340f"),
(x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1",x"b98e",x"403d",x"37b0",x"3bff",x"a3ef",x"2511",x"3606",x"33d1",x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b"),
(x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b",x"b98e",x"4045",x"37d0",x"3c00",x"9fe2",x"868d",x"360b",x"339c",x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380",x"b98e",x"404a",x"37dc",x"3bfd",x"1481",x"a9d9",x"360c",x"337d",x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"b98d",x"404f",x"37c9",x"3b31",x"b5e3",x"b397",x"3600",x"3366",x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f",x"b98e",x"4050",x"37cd",x"3bfa",x"2874",x"2c13",x"3601",x"3360"),
(x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b98d",x"404f",x"37c9",x"3b31",x"b5e3",x"b397",x"3600",x"3366",x"b98d",x"4050",x"37b8",x"3bfa",x"2a69",x"2a66",x"35f8",x"3360"),
(x"b98d",x"404f",x"37aa",x"3a13",x"b891",x"34fa",x"35f4",x"336a",x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b98d",x"4050",x"37a7",x"3bff",x"20dd",x"25fd",x"35f2",x"3366"),
(x"b98d",x"404f",x"37aa",x"3a13",x"b891",x"34fa",x"35f4",x"336a",x"b98d",x"4050",x"37a7",x"3bff",x"20dd",x"25fd",x"35f2",x"3366",x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"b98d",x"404e",x"378e",x"3bf3",x"a432",x"2f1d",x"35ea",x"3376",x"b98c",x"404e",x"378b",x"3af6",x"b023",x"379b",x"35e8",x"3377",x"b98c",x"404a",x"3784",x"3bd5",x"a532",x"3276",x"35e9",x"338d"),
(x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377",x"b98d",x"404e",x"378e",x"3bf3",x"a432",x"2f1d",x"35ea",x"3376",x"b98d",x"404a",x"3790",x"3b10",x"ad8c",x"3760",x"35ed",x"338b"),
(x"b98d",x"404a",x"3790",x"3b10",x"ad8c",x"3760",x"35ed",x"338b",x"b98c",x"404a",x"3784",x"3bd5",x"a532",x"3276",x"35e9",x"338d",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"b98c",x"403d",x"3777",x"3bc4",x"a9cc",x"3386",x"35ef",x"33db",x"b98d",x"403d",x"3782",x"3b88",x"abb1",x"354b",x"35f4",x"33d9",x"b98b",x"4045",x"377f",x"3bc5",x"a6cf",x"3387",x"35eb",x"33ac"),
(x"b98d",x"403d",x"3782",x"3b88",x"abb1",x"354b",x"35f4",x"33d9",x"b98c",x"403d",x"3777",x"3bc4",x"a9cc",x"3386",x"35ef",x"33db",x"b98d",x"4032",x"3770",x"3be2",x"a025",x"3161",x"35f6",x"340d"),
(x"b98d",x"4032",x"3770",x"3be2",x"a025",x"3161",x"35f6",x"340d",x"b98d",x"4030",x"378d",x"3bfe",x"28c2",x"2138",x"3602",x"340f",x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8"),
(x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8",x"b990",x"403d",x"37a1",x"3bf5",x"2dc9",x"aa2b",x"3600",x"33d2",x"b992",x"4045",x"3794",x"3bd9",x"292f",x"3209",x"35f5",x"33a8"),
(x"b992",x"4045",x"3794",x"3bd9",x"292f",x"3209",x"35f5",x"33a8",x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b"),
(x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b",x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b994",x"404d",x"37a3",x"3bda",x"aea9",x"311c",x"35f5",x"337c"),
(x"b994",x"404d",x"37a3",x"3bda",x"aea9",x"311c",x"35f5",x"337c",x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e",x"b993",x"404f",x"37b7",x"3977",x"b9c7",x"2ec0",x"35fa",x"336e",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"b98e",x"4030",x"3797",x"3813",x"b281",x"3ab0",x"3640",x"2b01",x"b9ae",x"4031",x"37c0",x"1bc8",x"b48d",x"3bab",x"365d",x"2ab9",x"b98e",x"403d",x"37b0",x"3860",x"b445",x"3a59",x"363e",x"29b6"),
(x"b98e",x"403d",x"37b0",x"3860",x"b445",x"3a59",x"363e",x"29b6",x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b98e",x"4045",x"37d0",x"386c",x"b560",x"3a19",x"3640",x"28d0"),
(x"b98e",x"4045",x"37d0",x"386c",x"b560",x"3a19",x"3640",x"28d0",x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b98e",x"404a",x"37dc",x"3889",x"b0d3",x"3a7a",x"3643",x"2852"),
(x"b98e",x"404a",x"37dc",x"3889",x"b0d3",x"3a7a",x"3643",x"2852",x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b98e",x"404d",x"37db",x"3837",x"36a0",x"39ef",x"3644",x"2800"),
(x"b98e",x"4050",x"37cd",x"3534",x"3ad6",x"367a",x"3644",x"2773",x"b98e",x"404d",x"37db",x"3837",x"36a0",x"39ef",x"3644",x"2800",x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e"),
(x"b98d",x"4050",x"37b8",x"33c4",x"3bc1",x"28ed",x"3642",x"26f2",x"b98e",x"4050",x"37cd",x"3534",x"3ad6",x"367a",x"3644",x"2773",x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709"),
(x"b98d",x"4050",x"37a7",x"342d",x"3b51",x"b4ec",x"3641",x"268d",x"b98d",x"4050",x"37b8",x"33c4",x"3bc1",x"28ed",x"3642",x"26f2",x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c"),
(x"b98d",x"404e",x"378e",x"386f",x"39bf",x"b6b9",x"363c",x"25e5",x"b98d",x"4050",x"37a7",x"342d",x"3b51",x"b4ec",x"3641",x"268d",x"b995",x"404f",x"3789",x"3469",x"3b25",x"b5af",x"3644",x"25c3"),
(x"b995",x"404f",x"3789",x"3469",x"3b25",x"b5af",x"3644",x"25c3",x"b990",x"404e",x"378b",x"3682",x"3b4c",x"2987",x"363f",x"25d0",x"b98d",x"404e",x"378e",x"386f",x"39bf",x"b6b9",x"363c",x"25e5"),
(x"b98c",x"404e",x"378b",x"b828",x"3967",x"382f",x"3606",x"2d1e",x"b98e",x"404e",x"3782",x"b7ca",x"39ef",x"375f",x"3603",x"2d14",x"b987",x"404e",x"378c",x"b8b4",x"39be",x"35f4",x"3605",x"2d2d"),
(x"b98d",x"404e",x"378e",x"386f",x"39bf",x"b6b9",x"363c",x"25e5",x"b990",x"404e",x"378b",x"3682",x"3b4c",x"2987",x"363f",x"25d0",x"b98c",x"404e",x"378b",x"35f3",x"3b61",x"2ea6",x"363c",x"25cf"),
(x"b972",x"4033",x"376d",x"3a5a",x"b06c",x"38bc",x"3604",x"2ef0",x"b967",x"4034",x"3752",x"3aac",x"b05e",x"3846",x"35f7",x"2ef0",x"b972",x"4030",x"376e",x"3ab7",x"ada6",x"384a",x"3606",x"2f15"),
(x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b972",x"4033",x"376d",x"303b",x"ac06",x"3be9",x"3668",x"2c64",x"b97b",x"4032",x"3770",x"2cfa",x"29bc",x"3bf7",x"3663",x"2c4b"),
(x"b97b",x"4032",x"3770",x"2cfa",x"29bc",x"3bf7",x"3663",x"2c4b",x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c",x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62"),
(x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c",x"b97b",x"4032",x"3770",x"2cfa",x"29bc",x"3bf7",x"3663",x"2c4b",x"b98d",x"4032",x"3770",x"2ca2",x"a97a",x"3bf8",x"3655",x"2c46"),
(x"b9e8",x"4034",x"376d",x"bae5",x"b1fa",x"378a",x"361e",x"3499",x"b9e6",x"402f",x"376e",x"bafb",x"ad7a",x"37ae",x"3622",x"348b",x"b9f0",x"4034",x"3752",x"bafe",x"b17b",x"3746",x"3612",x"3497"),
(x"b9e6",x"402f",x"376e",x"ad21",x"068d",x"3bf9",x"360e",x"3357",x"b9e8",x"4034",x"376d",x"a5e3",x"adbf",x"3bf7",x"360e",x"333a",x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a"),
(x"b9e6",x"402f",x"376e",x"ad21",x"068d",x"3bf9",x"360e",x"3357",x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9d5",x"4031",x"3770",x"a935",x"1ec2",x"3bfe",x"3601",x"3350"),
(x"b9d5",x"4031",x"3770",x"a935",x"1ec2",x"3bfe",x"3601",x"3350",x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b",x"b9cd",x"4032",x"3770",x"ae75",x"aa87",x"3bf2",x"35fa",x"334a"),
(x"b9e2",x"3f95",x"37cf",x"bafd",x"36b2",x"b3e9",x"3562",x"3530",x"ba0b",x"3f58",x"3752",x"bb05",x"36a0",x"b3ae",x"3504",x"34fb",x"b9f7",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518"),
(x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"b9e2",x"3f95",x"37cf",x"b33d",x"35ad",x"3b41",x"3604",x"30cf"),
(x"b970",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce",x"b9a9",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"b9aa",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"b96e",x"3f46",x"3752",x"330f",x"b68f",x"3b14",x"35af",x"2b2d",x"b985",x"3f77",x"37bd",x"367e",x"b50c",x"3adc",x"3585",x"2cb9",x"b95a",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88"),
(x"b94a",x"3f58",x"3752",x"374a",x"b488",x"3ac0",x"35c3",x"2c17",x"b95a",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88",x"b985",x"3f77",x"37bd",x"367e",x"b50c",x"3adc",x"3585",x"2cb9"),
(x"b970",x"3f95",x"37ce",x"3af6",x"36ac",x"b42c",x"359e",x"2d3c",x"b981",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a",x"b95d",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91"),
(x"b9ce",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"b9f1",x"3f48",x"3752",x"b5a1",x"b590",x"3af3",x"3506",x"349f",x"ba0b",x"3f58",x"3752",x"b6ba",x"b4d8",x"3ad7",x"34fb",x"34bd"),
(x"b9a9",x"3f49",x"380d",x"3ac4",x"b843",x"a386",x"35e1",x"2e92",x"b9a9",x"3f49",x"382e",x"3a6c",x"b8c3",x"9624",x"35c9",x"2e91",x"b9a6",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1"),
(x"b9a9",x"3f49",x"380d",x"ba6f",x"b8bf",x"a6fd",x"356a",x"3496",x"b9aa",x"3f4b",x"380c",x"bb52",x"b656",x"ac81",x"3569",x"3499",x"b9ad",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c"),
(x"b9a6",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1",x"b970",x"3f95",x"37ce",x"3b84",x"b57a",x"175f",x"35fa",x"3035",x"b985",x"3f77",x"37bd",x"3b7c",x"b5a3",x"a1ae",x"3602",x"2fb5"),
(x"b9ad",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c",x"b9aa",x"3f4b",x"380c",x"bb52",x"b656",x"ac81",x"3569",x"3499",x"b9ce",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd"),
(x"b98b",x"3f82",x"3752",x"381e",x"3818",x"b980",x"35d8",x"2d45",x"b95d",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91",x"b981",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a"),
(x"b9d3",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"b9f7",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518",x"b9d2",x"3f71",x"3752",x"b43c",x"3773",x"bac1",x"3517",x"3533"),
(x"b982",x"4072",x"3752",x"39fd",x"0000",x"394d",x"35ef",x"2c07",x"b982",x"405c",x"3752",x"39fd",x"0000",x"394d",x"35ef",x"2cfe",x"b9b1",x"405c",x"37be",x"39fd",x"0000",x"394d",x"3625",x"2d00"),
(x"b9e2",x"405e",x"3752",x"b9ee",x"0a8d",x"395e",x"360a",x"2d16",x"b9e2",x"4071",x"3752",x"b9ee",x"0cea",x"395e",x"360a",x"2df8",x"b9b1",x"4072",x"37be",x"b9ee",x"0a8d",x"395e",x"3641",x"2dfd"),
(x"b9b2",x"407a",x"3802",x"b837",x"b93f",x"3851",x"35b4",x"2aa4",x"b9b1",x"4072",x"37be",x"b8a6",x"b8cf",x"3862",x"35c5",x"2b97",x"b9e2",x"4071",x"3752",x"b837",x"b940",x"3851",x"35fc",x"2bb2"),
(x"b982",x"4072",x"3752",x"3854",x"b926",x"3853",x"3516",x"34a2",x"b9b1",x"4072",x"37be",x"38df",x"b892",x"3866",x"354c",x"349f",x"b9b2",x"407a",x"3802",x"3854",x"b926",x"3853",x"355f",x"3481"),
(x"b9e8",x"3f49",x"3754",x"bab7",x"9f2b",x"3858",x"34ae",x"259c",x"b9a9",x"3f4b",x"380f",x"bac7",x"a224",x"383e",x"3455",x"2566",x"b9aa",x"3dc3",x"3804",x"bab6",x"9af6",x"385a",x"345b",x"311f"),
(x"b96c",x"3f46",x"3755",x"3abd",x"9ffc",x"384e",x"34af",x"25db",x"b96c",x"3dc2",x"3752",x"3a9d",x"90ea",x"3880",x"34b4",x"3123",x"b9aa",x"3dc3",x"3804",x"3abc",x"9c9b",x"3850",x"3507",x"311e"),
(x"ba0f",x"3db3",x"3752",x"b8d1",x"395c",x"36f1",x"348c",x"3524",x"b9e7",x"3dc2",x"3752",x"b873",x"3a03",x"35ad",x"349d",x"3544",x"b9aa",x"3dc3",x"3804",x"b8d1",x"395c",x"36f1",x"34f0",x"3544"),
(x"b9aa",x"3dc3",x"3804",x"38d0",x"395f",x"36e9",x"3493",x"3520",x"b96c",x"3dc2",x"3752",x"388b",x"39de",x"35f7",x"34e6",x"3520",x"b945",x"3db3",x"3752",x"38d0",x"395f",x"36e9",x"34f7",x"3500"),
(x"ba10",x"3d4c",x"3752",x"ba6d",x"1c32",x"38c3",x"3512",x"263e",x"ba0f",x"3db3",x"3752",x"ba6b",x"19bc",x"38c5",x"3513",x"2bf1",x"b9a9",x"3db1",x"3832",x"ba6c",x"1b5f",x"38c4",x"358f",x"2bd9"),
(x"b9a9",x"3db1",x"3832",x"3a6f",x"1d6d",x"38c0",x"3587",x"3369",x"b945",x"3db3",x"3752",x"3a75",x"20ea",x"38b8",x"3507",x"3363",x"b942",x"3d4d",x"3752",x"3a6f",x"1d6d",x"38c0",x"3505",x"3446"),
(x"b946",x"3cfa",x"3872",x"9b5f",x"b9fc",x"394f",x"34fa",x"34f8",x"b943",x"3ca2",x"3752",x"928d",x"b9fe",x"394b",x"34fa",x"3435",x"ba11",x"3ca2",x"3752",x"9ac2",x"b9fc",x"394e",x"345f",x"3435"),
(x"b943",x"351b",x"3752",x"0e8d",x"3a2a",x"3918",x"34fa",x"32b2",x"b945",x"3397",x"3877",x"9ffc",x"3a32",x"390e",x"34fa",x"3130",x"ba10",x"3396",x"3874",x"0e8d",x"3a2a",x"3918",x"3461",x"3131"),
(x"ba10",x"3396",x"3874",x"96f6",x"ba26",x"391d",x"3465",x"3428",x"b945",x"3397",x"3877",x"9dd6",x"ba2a",x"3918",x"34f9",x"3428",x"b943",x"30ef",x"3752",x"9624",x"ba26",x"391d",x"34f9",x"32bf"),
(x"b9ff",x"401f",x"3786",x"baf9",x"ae2b",x"37ae",x"3620",x"344a",x"ba0f",x"4020",x"3752",x"bacd",x"aeb3",x"381f",x"3609",x"344a",x"ba05",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"360a",x"345b"),
(x"b9f8",x"4024",x"378d",x"ba5b",x"36b9",x"3703",x"3622",x"3459",x"ba05",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"360a",x"345b",x"b9fc",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"360c",x"3464"),
(x"b9f2",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3624",x"3460",x"b9fc",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"360c",x"3464",x"b9f4",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"360e",x"346a"),
(x"b9f8",x"400d",x"3752",x"bae9",x"b336",x"3733",x"361b",x"3412",x"ba0f",x"4020",x"3752",x"bacd",x"aeb3",x"381f",x"3609",x"344a",x"b9ff",x"401f",x"3786",x"baf9",x"ae2b",x"37ae",x"3620",x"344a"),
(x"b9f0",x"4002",x"3752",x"bb07",x"b070",x"374f",x"3623",x"33e8",x"b9f8",x"400d",x"3752",x"bae9",x"b336",x"3733",x"361b",x"3412",x"b9f0",x"400d",x"3777",x"bb0c",x"b28a",x"36d3",x"362a",x"3414"),
(x"b9dc",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"362c",x"346e",x"b9f4",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"360e",x"346a",x"b9d5",x"4024",x"3782",x"3904",x"3a39",x"a8ac",x"362c",x"3476"),
(x"b9f0",x"400d",x"3777",x"9d6d",x"aedf",x"3bf4",x"3578",x"34f2",x"b9e8",x"400d",x"3776",x"349f",x"a9d6",x"3ba6",x"357d",x"34f3",x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9e8",x"400d",x"3776",x"349f",x"a9d6",x"3ba6",x"357d",x"34f3",x"b9f0",x"400d",x"3777",x"9d6d",x"aedf",x"3bf4",x"3578",x"34f2"),
(x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9ff",x"401f",x"3786",x"b0fd",x"b014",x"3bd6",x"356f",x"3528",x"b9f8",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3575",x"3536"),
(x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9f8",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3575",x"3536",x"b9f2",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"357a",x"353b"),
(x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9f2",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"357a",x"353b",x"b9e7",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3582",x"353d"),
(x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9e7",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3582",x"353d",x"b9dc",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9e0",x"4025",x"378f",x"b17c",x"b4ab",x"3b87",x"3587",x"3537",x"b9dc",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"b9d7",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"358e",x"3523",x"b9cf",x"4022",x"378b",x"2ef6",x"b0cc",x"3bdc",x"3594",x"352f",x"b9ce",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9d3",x"4023",x"378c",x"287a",x"ad2b",x"3bf8",x"3591",x"3531",x"b9cf",x"4022",x"378b",x"2ef6",x"b0cc",x"3bdc",x"3594",x"352f"),
(x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9d7",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"358e",x"3523",x"b9ce",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"b9d7",x"400e",x"3777",x"ac2d",x"ae61",x"3bf1",x"358b",x"34f3",x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9cf",x"4017",x"377f",x"27d5",x"aef0",x"3bf2",x"3593",x"350f"),
(x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9d7",x"400e",x"3777",x"ac2d",x"ae61",x"3bf1",x"358b",x"34f3",x"b9cf",x"400d",x"3777",x"abbe",x"ace8",x"3bf6",x"3591",x"34f1"),
(x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9d7",x"400e",x"3777",x"ac2d",x"ae61",x"3bf1",x"358b",x"34f3",x"b9dc",x"400e",x"3775",x"b232",x"ad32",x"3bd2",x"3587",x"34f5"),
(x"b9d9",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"358b",x"3511",x"b9df",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3586",x"3512",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523"),
(x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9d7",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"358e",x"3523",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523"),
(x"b9d9",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"358c",x"3530",x"b9dd",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3589",x"352f",x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534"),
(x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9e0",x"4025",x"378f",x"b17c",x"b4ab",x"3b87",x"3587",x"3537",x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534"),
(x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9e6",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3583",x"3539",x"b9e7",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3581",x"3535"),
(x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9ee",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"357c",x"3538",x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534"),
(x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9f3",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3578",x"3534",x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"b9e8",x"400d",x"3776",x"349f",x"a9d6",x"3ba6",x"357d",x"34f3",x"b9f7",x"401f",x"3788",x"30d4",x"aed9",x"3bdc",x"3574",x"3528",x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527"),
(x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"b9df",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3586",x"3512",x"b9dc",x"400e",x"3775",x"b232",x"ad32",x"3bd2",x"3587",x"34f5",x"b9e5",x"400e",x"3773",x"2c3e",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523",x"b9df",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3586",x"3512",x"b9f3",x"401f",x"3782",x"3116",x"adf8",x"3bdc",x"3578",x"3527"),
(x"b9dd",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3589",x"352f",x"b9db",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"358a",x"3523",x"b9f0",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"b9e3",x"4024",x"3787",x"b4c3",x"b627",x"3afd",x"3585",x"3534",x"b9dd",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3589",x"352f",x"b9ec",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"357e",x"3534"),
(x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f",x"b9cb",x"400d",x"378a",x"bbec",x"2694",x"3049",x"3648",x"317b",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b"),
(x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b",x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f",x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140"),
(x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108",x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b",x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a"),
(x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff",x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108",x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"b9c6",x"4023",x"37b6",x"b9d1",x"b94b",x"31cf",x"3644",x"30fb",x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff",x"b9cd",x"4024",x"37aa",x"ba49",x"b805",x"35c1",x"364a",x"30f4"),
(x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9c6",x"4023",x"37b6",x"b9d1",x"b94b",x"31cf",x"3644",x"30fb",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9c6",x"4022",x"37c1",x"ba68",x"b74a",x"b638",x"3640",x"30fb",x"b9cd",x"4023",x"37c8",x"bb6a",x"b4dc",x"b301",x"363e",x"30f1",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112"),
(x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133"),
(x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133",x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174",x"b9cb",x"400d",x"37b2",x"bbee",x"a8fd",x"2fea",x"3638",x"3174",x"b9cc",x"3fff",x"3798",x"bbe2",x"a7a0",x"314e",x"363a",x"31c7"),
(x"b9cb",x"400d",x"37b2",x"bbee",x"a8fd",x"2fea",x"3638",x"3174",x"b9cc",x"400d",x"37a7",x"bbb8",x"2e24",x"b3c9",x"363c",x"3174",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133"),
(x"b9cc",x"4017",x"37d1",x"bbf6",x"a89b",x"2d9b",x"3632",x"3134",x"b9cc",x"4018",x"37c6",x"bb58",x"3009",x"b603",x"3636",x"3133",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112"),
(x"b9cc",x"401d",x"37de",x"bbe7",x"9e8d",x"30f2",x"3631",x"3110",x"b9cd",x"401d",x"37d4",x"bb44",x"2839",x"b6a9",x"3635",x"3112",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"b9cc",x"4022",x"37dc",x"bbdb",x"2a31",x"31d8",x"3635",x"30f7",x"b9cd",x"4021",x"37d2",x"bb5b",x"afb9",x"b5f8",x"3638",x"30fb",x"b9cd",x"4023",x"37c8",x"bb6a",x"b4dc",x"b301",x"363e",x"30f1"),
(x"b9cc",x"4024",x"37cc",x"bbf1",x"2b1a",x"2ec3",x"363d",x"30ea",x"b9cd",x"4023",x"37c8",x"bb6a",x"b4dc",x"b301",x"363e",x"30f1",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9cd",x"4025",x"37a7",x"bbff",x"21bc",x"2518",x"364c",x"30ed",x"b9cd",x"4025",x"37b8",x"bbfc",x"2752",x"2a48",x"3645",x"30e8",x"b9cd",x"4024",x"37b7",x"bb1c",x"b755",x"a280",x"3645",x"30ee"),
(x"b9cd",x"4025",x"37a7",x"bbff",x"21bc",x"2518",x"364c",x"30ed",x"b9cd",x"4024",x"37aa",x"ba49",x"b805",x"35c1",x"364a",x"30f4",x"b9cd",x"4021",x"3799",x"bafb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a",x"b9ce",x"401e",x"3784",x"bbd5",x"a432",x"3276",x"3656",x"311b",x"b9ce",x"4022",x"378e",x"bbf3",x"a2c2",x"2ede",x"3654",x"3100"),
(x"b9ce",x"401e",x"3784",x"bbd5",x"a432",x"3276",x"3656",x"311b",x"b9cd",x"401e",x"3790",x"bad6",x"aec5",x"3810",x"3651",x"311a",x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140"),
(x"b9cf",x"4017",x"377f",x"bbc6",x"a57a",x"337e",x"3654",x"3142",x"b9cd",x"4017",x"378b",x"baba",x"aa69",x"384e",x"364f",x"3140",x"b9cd",x"400d",x"3783",x"bb43",x"aa24",x"36a7",x"364a",x"317b"),
(x"b9cb",x"400d",x"378a",x"bbec",x"2694",x"3049",x"3648",x"317b",x"b9ca",x"400d",x"379f",x"bbf8",x"2d3a",x"a850",x"3640",x"3175",x"b9cd",x"3fff",x"3790",x"bbfe",x"2874",x"9fc8",x"363d",x"31c9"),
(x"b9ca",x"400d",x"379f",x"bbf8",x"2d3a",x"a850",x"3640",x"3175",x"b9cb",x"400d",x"378a",x"bbec",x"2694",x"3049",x"3648",x"317b",x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f"),
(x"b9c6",x"4018",x"37ba",x"bbdd",x"2e26",x"b0f1",x"363d",x"3133",x"b9c8",x"4017",x"3794",x"bbb1",x"25b5",x"345f",x"364a",x"313f",x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b"),
(x"b9c6",x"401d",x"37c9",x"bbcd",x"2c2d",x"b2c5",x"363b",x"3114",x"b9c8",x"401d",x"3798",x"bbae",x"a82f",x"3470",x"364c",x"311b",x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108"),
(x"b9c6",x"4021",x"37c7",x"bb8c",x"a849",x"b548",x"363e",x"3102",x"b9c6",x"4021",x"37a3",x"bbab",x"abf9",x"346d",x"3649",x"3108",x"b9c6",x"4022",x"37ac",x"bb0b",x"b542",x"3578",x"3647",x"30ff"),
(x"b9cb",x"400d",x"37b2",x"b866",x"b31b",x"3a70",x"35df",x"33e6",x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b9ae",x"3ffe",x"37c0",x"2418",x"b372",x"3bc7",x"35c2",x"341c"),
(x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b9cb",x"400d",x"37b2",x"b866",x"b31b",x"3a70",x"35df",x"33e6",x"b9cc",x"4017",x"37d1",x"b86f",x"b4aa",x"3a3c",x"35de",x"33a2"),
(x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b9cc",x"4017",x"37d1",x"b86f",x"b4aa",x"3a3c",x"35de",x"33a2",x"b9cc",x"401d",x"37de",x"b896",x"af43",x"3a7d",x"35db",x"337c"),
(x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b9cc",x"401d",x"37de",x"b896",x"af43",x"3a7d",x"35db",x"337c",x"b9cc",x"4022",x"37dc",x"b830",x"3619",x"3a17",x"35d9",x"3360"),
(x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351",x"b9ac",x"4024",x"37fd",x"23bb",x"3849",x"3ac0",x"35c1",x"3362",x"b9cc",x"4022",x"37dc",x"b830",x"3619",x"3a17",x"35d9",x"3360"),
(x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341",x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351",x"b9cc",x"4024",x"37cc",x"b5be",x"3a7e",x"375e",x"35d9",x"334c"),
(x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331",x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341",x"b9cd",x"4025",x"37b8",x"b483",x"3bab",x"291b",x"35da",x"333c"),
(x"b9c4",x"4025",x"379c",x"b51a",x"3ab3",x"b716",x"35d5",x"3325",x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331",x"b9cd",x"4025",x"37a7",x"b469",x"3b1b",x"b5df",x"35db",x"332f"),
(x"b9d3",x"4023",x"378c",x"3949",x"390d",x"367c",x"3632",x"3477",x"b9d5",x"4024",x"3782",x"3904",x"3a39",x"a8ac",x"362c",x"3476",x"b9cd",x"4022",x"3786",x"3818",x"3947",x"3865",x"3631",x"347c"),
(x"b9cd",x"4022",x"3786",x"b6de",x"3aa3",x"35b2",x"35df",x"3313",x"b9ca",x"4023",x"378b",x"b8bf",x"3a5d",x"afac",x"35dc",x"3317",x"b9ce",x"4022",x"378e",x"b717",x"3a25",x"b764",x"35e0",x"3319"),
(x"b95b",x"401f",x"3786",x"3ae5",x"ae76",x"37f1",x"3652",x"3477",x"b962",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3655",x"3468",x"b956",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"363c",x"3466"),
(x"b962",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3655",x"3468",x"b968",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3656",x"3461",x"b95e",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"363e",x"345e"),
(x"b968",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3656",x"3461",x"b973",x"4027",x"378f",x"a731",x"3bb3",x"3450",x"365a",x"345a",x"b966",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"3640",x"3458"),
(x"b95b",x"401f",x"3786",x"3ae5",x"ae76",x"37f1",x"3652",x"3477",x"b94b",x"4020",x"3752",x"3acd",x"aeb3",x"381f",x"363b",x"3478",x"b962",x"400d",x"3752",x"3aca",x"b303",x"37b2",x"364e",x"34af"),
(x"b96c",x"400d",x"3775",x"3abf",x"b1e9",x"3808",x"365d",x"34ae",x"b962",x"400d",x"3752",x"3aca",x"b303",x"37b2",x"364e",x"34af",x"b967",x"4002",x"3752",x"3ab1",x"af0f",x"3849",x"3656",x"34ce"),
(x"b985",x"4024",x"3782",x"b907",x"3a38",x"a54c",x"365e",x"344b",x"b966",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"3640",x"3458",x"b97e",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"365e",x"3453"),
(x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0",x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079",x"b96c",x"400d",x"3775",x"2b97",x"ae90",x"3bf1",x"3642",x"307d"),
(x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079",x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e",x"b95b",x"401f",x"3786",x"2e5c",x"b067",x"3be2",x"363e",x"300d"),
(x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e",x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee",x"b962",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3645",x"2fe4"),
(x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee",x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf",x"b968",x"4026",x"378e",x"2d5c",x"a067",x"3bf8",x"364b",x"2fd2"),
(x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf",x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd",x"b973",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3653",x"2fce"),
(x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd",x"b97a",x"4025",x"378f",x"317c",x"b4aa",x"3b87",x"3658",x"2fe7",x"b97e",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"365b",x"2fdd"),
(x"b97e",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"365b",x"2fdd",x"b97a",x"4025",x"378f",x"317c",x"b4aa",x"3b87",x"3658",x"2fe7",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003"),
(x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003",x"b98c",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3664",x"3007",x"b987",x"4023",x"378c",x"a87a",x"ad2b",x"3bf8",x"3661",x"3001"),
(x"b983",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"365c",x"301d",x"b98c",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3662",x"3020",x"b98c",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3664",x"3007"),
(x"b98c",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3662",x"3020",x"b983",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"365c",x"301d",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040"),
(x"b98b",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"365f",x"3047",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040",x"b983",x"400e",x"3777",x"2c32",x"ae3d",x"3bf1",x"3654",x"307b"),
(x"b98c",x"400d",x"3777",x"296a",x"ace7",x"3bf8",x"365a",x"3081",x"b983",x"400e",x"3777",x"2c32",x"ae3d",x"3bf1",x"3654",x"307b",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"b97e",x"400e",x"3775",x"3224",x"ad11",x"3bd3",x"3651",x"3077",x"b983",x"400e",x"3777",x"2c32",x"ae3d",x"3bf1",x"3654",x"307b",x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040"),
(x"b981",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"3658",x"3040",x"b983",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"365c",x"301d",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b"),
(x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b",x"b983",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"365c",x"301d",x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003"),
(x"b981",x"4022",x"378c",x"327a",x"b213",x"3baf",x"365c",x"3003",x"b97a",x"4025",x"378f",x"317c",x"b4aa",x"3b87",x"3658",x"2fe7",x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5",x"b97a",x"4025",x"378f",x"317c",x"b4aa",x"3b87",x"3658",x"2fe7",x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd"),
(x"b973",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"b975",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3654",x"2fdd",x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf"),
(x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b96c",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"364d",x"2fdf",x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee"),
(x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b967",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3648",x"2fee",x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e"),
(x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b963",x"401f",x"3788",x"b153",x"afe4",x"3bd3",x"3643",x"300e",x"b972",x"400d",x"3776",x"aff7",x"ad4e",x"3be9",x"3647",x"3079"),
(x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079",x"b979",x"4001",x"376f",x"2217",x"aa2e",x"3bfd",x"3646",x"30c0",x"b985",x"4002",x"3770",x"2bef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"b975",x"400e",x"3773",x"ac28",x"abec",x"3bf7",x"3649",x"3079",x"b97e",x"400e",x"3775",x"3224",x"ad11",x"3bd3",x"3651",x"3077",x"b97b",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3653",x"303e"),
(x"b967",x"401f",x"3782",x"b115",x"adfa",x"3bdc",x"3647",x"3011",x"b97b",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3653",x"303e",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b"),
(x"b96a",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"364b",x"2ffc",x"b97f",x"401e",x"3782",x"315c",x"b078",x"3bce",x"3658",x"301b",x"b97d",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3658",x"3004"),
(x"b96e",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"364e",x"2ff0",x"b97d",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3658",x"3004",x"b977",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"b98f",x"400d",x"378a",x"3bdf",x"2581",x"319c",x"365f",x"2e8f",x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03",x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05",x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50",x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e",x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74"),
(x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f",x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89"),
(x"b98d",x"4024",x"37aa",x"3a75",x"b7d2",x"354a",x"3662",x"2f9c",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89",x"b993",x"4023",x"37b7",x"39e1",x"b96b",x"23fc",x"365c",x"2f93"),
(x"b993",x"4023",x"37b7",x"39e1",x"b96b",x"23fc",x"365c",x"2f93",x"b993",x"4022",x"37c3",x"3af0",x"b4e6",x"b647",x"3658",x"2f91",x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"b993",x"4022",x"37c3",x"3af0",x"b4e6",x"b647",x"3658",x"2f91",x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c"),
(x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b98e",x"400d",x"37a5",x"3b77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"b98e",x"400d",x"37b0",x"3bfb",x"a724",x"2bb7",x"3651",x"2e9c",x"b98e",x"400d",x"37a5",x"3b77",x"2f4d",x"b571",x"3655",x"2e9c",x"b98f",x"3ffd",x"378d",x"3bfd",x"9d53",x"29ab",x"3655",x"2de8"),
(x"b98e",x"400d",x"37b0",x"3bfb",x"a724",x"2bb7",x"3651",x"2e9c",x"b98e",x"4017",x"37d0",x"3c00",x"9e59",x"868d",x"364a",x"2f1c",x"b98e",x"4018",x"37c6",x"3b32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"b98e",x"4017",x"37d0",x"3c00",x"9e59",x"868d",x"364a",x"2f1c",x"b98e",x"401d",x"37dc",x"3bfd",x"135f",x"a9d9",x"364a",x"2f66",x"b98e",x"401d",x"37d2",x"3afe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"b98e",x"401d",x"37dc",x"3bfd",x"135f",x"a9d9",x"364a",x"2f66",x"b98e",x"4022",x"37db",x"3bff",x"1b2b",x"2560",x"364e",x"2f95",x"b98e",x"4021",x"37d0",x"3b35",x"af71",x"b6b0",x"3651",x"2f8c"),
(x"b98e",x"4022",x"37db",x"3bff",x"1b2b",x"2560",x"364e",x"2f95",x"b98e",x"4024",x"37cd",x"3bf5",x"2bb1",x"2d1b",x"3655",x"2fb0",x"b98d",x"4023",x"37c9",x"3b3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"b98e",x"4024",x"37cd",x"3bf5",x"2bb1",x"2d1b",x"3655",x"2fb0",x"b98d",x"4025",x"37b8",x"3bfd",x"20a8",x"29ed",x"365e",x"2fb3",x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7"),
(x"b98d",x"4024",x"37b7",x"3b7d",x"b59c",x"2594",x"365e",x"2fa7",x"b98d",x"4025",x"37b8",x"3bfd",x"20a8",x"29ed",x"365e",x"2fb3",x"b98d",x"4025",x"37a7",x"3bff",x"1fc8",x"25fd",x"3664",x"2fa8"),
(x"b98d",x"4025",x"37a7",x"3bff",x"1fc8",x"25fd",x"3664",x"2fa8",x"b98d",x"4022",x"378e",x"3bf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"b98d",x"4021",x"3798",x"3aff",x"b392",x"36c4",x"3668",x"2f7f"),
(x"b98d",x"4022",x"378e",x"3bf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"b98c",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"366e",x"2f4e",x"b98d",x"401e",x"3790",x"3ad4",x"ae75",x"3815",x"3669",x"2f50"),
(x"b98c",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"366e",x"2f4e",x"b98b",x"4017",x"377f",x"3bc6",x"a57a",x"3387",x"366c",x"2f00",x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03"),
(x"b98d",x"400d",x"3782",x"3b3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"b98d",x"4017",x"378b",x"3aba",x"aab1",x"384d",x"3667",x"2f03",x"b98b",x"4017",x"377f",x"3bc6",x"a57a",x"3387",x"366c",x"2f00"),
(x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b98f",x"400d",x"378a",x"3bdf",x"2581",x"319c",x"365f",x"2e8f",x"b98d",x"4000",x"3770",x"3be7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"b990",x"400d",x"37a1",x"3bfd",x"2a97",x"9553",x"3657",x"2e9c",x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b992",x"4017",x"3794",x"3bcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"b993",x"4018",x"37be",x"3be0",x"2e19",x"b0b1",x"3654",x"2f20",x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b992",x"401d",x"3798",x"3bbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"b994",x"401d",x"37c9",x"3bcf",x"2b2e",x"b2a8",x"3653",x"2f5a",x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b994",x"4021",x"37a3",x"3bbc",x"ae61",x"3382",x"3662",x"2f74"),
(x"b993",x"4021",x"37c9",x"3b92",x"ad65",x"b4fc",x"3655",x"2f83",x"b993",x"4022",x"37c3",x"3af0",x"b4e6",x"b647",x"3658",x"2f91",x"b993",x"4022",x"37ac",x"3b40",x"b55d",x"341d",x"3660",x"2f89"),
(x"b9ae",x"3ffe",x"37c0",x"2418",x"b372",x"3bc7",x"35c2",x"341c",x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b98e",x"400d",x"37b0",x"3883",x"b339",x"3a5a",x"35a4",x"33e7"),
(x"b9ac",x"400d",x"37dc",x"21fd",x"b51b",x"3b94",x"35c1",x"33de",x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b98e",x"4017",x"37d0",x"3883",x"b46b",x"3a39",x"35a5",x"33a3"),
(x"b9ae",x"4019",x"3800",x"22f6",x"b49e",x"3ba8",x"35c2",x"3397",x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b98e",x"401d",x"37dc",x"388e",x"afce",x"3a80",x"35a7",x"337c"),
(x"b9ad",x"401f",x"3804",x"2194",x"2a70",x"3bfd",x"35c2",x"3379",x"b9ac",x"4024",x"37fd",x"23bb",x"3849",x"3ac0",x"35c1",x"3362",x"b98e",x"4022",x"37db",x"3859",x"3581",x"3a1f",x"35a9",x"3362"),
(x"b98e",x"4022",x"37db",x"3859",x"3581",x"3a1f",x"35a9",x"3362",x"b9ac",x"4024",x"37fd",x"23bb",x"3849",x"3ac0",x"35c1",x"3362",x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351"),
(x"b98e",x"4024",x"37cd",x"3609",x"3a62",x"3783",x"35aa",x"334e",x"b9ac",x"4026",x"37e2",x"1c81",x"3a99",x"3885",x"35c1",x"3351",x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341"),
(x"b98d",x"4025",x"37b8",x"34be",x"3ba1",x"2a04",x"35a8",x"333e",x"b9ac",x"4027",x"37c9",x"1987",x"3bd9",x"322d",x"35c1",x"3341",x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331"),
(x"b98d",x"4025",x"37a7",x"34f8",x"3b04",x"b5db",x"35a6",x"3332",x"b9ac",x"4027",x"37b3",x"2887",x"3bce",x"b2e4",x"35c0",x"3331",x"b995",x"4024",x"3789",x"3533",x"3ac8",x"b6b3",x"35a9",x"3318"),
(x"b98e",x"4022",x"3782",x"b856",x"3952",x"381b",x"3662",x"3443",x"b985",x"4024",x"3782",x"b907",x"3a38",x"a54c",x"365e",x"344b",x"b987",x"4023",x"378c",x"b932",x"391d",x"3694",x"3664",x"344a"),
(x"b990",x"4023",x"378b",x"37bd",x"3afd",x"2a63",x"35a4",x"331a",x"b98e",x"4022",x"3782",x"3717",x"3b28",x"2aab",x"35a3",x"3313",x"b98c",x"4022",x"378b",x"371a",x"3b19",x"2ff2",x"35a0",x"3319"),
(x"b967",x"4002",x"3752",x"3ab1",x"af0f",x"3849",x"3656",x"34ce",x"b96d",x"3ff0",x"3752",x"3ae0",x"aed4",x"37ff",x"365d",x"34ec",x"b972",x"3ffb",x"376e",x"3ab9",x"ac8e",x"384b",x"3665",x"34da"),
(x"b972",x"4001",x"376d",x"303c",x"aa80",x"3beb",x"3641",x"30bf",x"b972",x"3ffb",x"376e",x"312d",x"21ae",x"3be4",x"363f",x"30d7",x"b97b",x"3fff",x"3770",x"2d3d",x"28c9",x"3bf7",x"3647",x"30ce"),
(x"b9e6",x"3ff8",x"376e",x"bafe",x"ac6a",x"37b1",x"3633",x"33c7",x"b9ec",x"3fef",x"3752",x"bb01",x"ac96",x"37a2",x"362b",x"33a9",x"b9f0",x"4002",x"3752",x"bb07",x"b070",x"374f",x"3623",x"33e8"),
(x"b9e1",x"4002",x"376f",x"8e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"b9d5",x"4002",x"3770",x"ac6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"b9d5",x"3ffc",x"3770",x"a935",x"1d6d",x"3bfe",x"3589",x"34c5"),
(x"b9ff",x"404b",x"3786",x"baf5",x"afa4",x"37a8",x"3610",x"34de",x"ba0f",x"404c",x"3752",x"bac8",x"b025",x"381c",x"35f9",x"34dd",x"ba05",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35fb",x"34ec"),
(x"b9f8",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"3613",x"34eb",x"ba05",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35fb",x"34ec",x"b9fc",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35fd",x"34f4"),
(x"b9f2",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"3615",x"34f1",x"b9fc",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35fd",x"34f4",x"b9f4",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35ff",x"34f9"),
(x"b9f8",x"403d",x"3752",x"bad1",x"b46a",x"371a",x"360a",x"34b0",x"ba0f",x"404c",x"3752",x"bac8",x"b025",x"381c",x"35f9",x"34dd",x"b9ff",x"404b",x"3786",x"baf5",x"afa4",x"37a8",x"3610",x"34de"),
(x"b9f0",x"4034",x"3752",x"bafe",x"b17b",x"3746",x"3612",x"3497",x"b9f8",x"403d",x"3752",x"bad1",x"b46a",x"371a",x"360a",x"34b0",x"b9f0",x"403d",x"3777",x"baf8",x"b403",x"36bf",x"3619",x"34b3"),
(x"b9dc",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"361c",x"34ff",x"b9f4",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35ff",x"34f9",x"b9d5",x"404f",x"3782",x"385b",x"3ab4",x"a80e",x"361b",x"3507"),
(x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9e8",x"4034",x"376d",x"a5e3",x"adbf",x"3bf7",x"360e",x"333a"),
(x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9f0",x"403d",x"3777",x"253f",x"b05f",x"3bec",x"3611",x"3305"),
(x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9ff",x"404b",x"3786",x"b0f8",x"b10b",x"3bcd",x"3619",x"32ae",x"b9f8",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3613",x"3297"),
(x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9f8",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3613",x"3297",x"b9f2",x"4051",x"378e",x"ad5b",x"a187",x"3bf8",x"360e",x"328f"),
(x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9f2",x"4051",x"378e",x"ad5b",x"a187",x"3bf8",x"360e",x"328f",x"b9e7",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9e6",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3605",x"3292",x"b9e7",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9dc",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"35fe",x"3292"),
(x"b9d7",x"404a",x"3788",x"ac6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"b9cf",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"35f4",x"32a5",x"b9ce",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9d3",x"404e",x"378c",x"2877",x"ae68",x"3bf4",x"35f7",x"32a1",x"b9cf",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"35f4",x"32a5"),
(x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9d7",x"404a",x"3788",x"ac6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"b9ce",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"b9d7",x"403d",x"3777",x"ac2a",x"afe7",x"3beb",x"35fe",x"3305",x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9cf",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"35f6",x"32d9"),
(x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b",x"b9d7",x"403d",x"3777",x"ac2a",x"afe7",x"3beb",x"35fe",x"3305",x"b9cf",x"403d",x"3777",x"abbb",x"ae16",x"3bf2",x"35f8",x"3309"),
(x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9d7",x"403d",x"3777",x"ac2a",x"afe7",x"3beb",x"35fe",x"3305",x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"b9d9",x"4045",x"3780",x"b169",x"b087",x"3bcd",x"35fd",x"32d5",x"b9df",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3602",x"32d4",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9d7",x"404a",x"3788",x"ac6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9d9",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"35fc",x"32a3",x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4"),
(x"b9e6",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3605",x"3292",x"b9e0",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3601",x"3296",x"b9e3",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3603",x"329c"),
(x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9e6",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3605",x"3292",x"b9e7",x"4050",x"3787",x"2710",x"b98f",x"39bf",x"3606",x"329a"),
(x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9ee",x"4050",x"378f",x"2d72",x"b63f",x"3b55",x"360c",x"3294",x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b"),
(x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9f3",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3610",x"329a",x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1"),
(x"b9e8",x"403d",x"3776",x"3339",x"accc",x"3bc5",x"360c",x"3304",x"b9f7",x"404c",x"3788",x"30d1",x"b03c",x"3bd6",x"3614",x"32ae",x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9e5",x"403d",x"3773",x"2db8",x"ad34",x"3bf1",x"3609",x"3304",x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"b9df",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3602",x"32d4",x"b9dc",x"403e",x"3775",x"b0b9",x"adbc",x"3be1",x"3602",x"3302",x"b9e5",x"403d",x"3773",x"2db8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7",x"b9df",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3602",x"32d4",x"b9f3",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4",x"b9db",x"404b",x"3782",x"b155",x"b185",x"3bc4",x"35fe",x"32b7",x"b9f0",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"360d",x"32a1"),
(x"b9e3",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3603",x"329c",x"b9dd",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"35ff",x"32a4",x"b9ec",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"360a",x"329b"),
(x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9cd",x"403d",x"3783",x"bb8f",x"ab5c",x"3527",x"35a7",x"34a3",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c",x"b9c8",x"4045",x"3794",x"bbbc",x"287e",x"3408",x"35a6",x"348a",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c",x"b9cd",x"404a",x"3790",x"bb17",x"ade0",x"3741",x"35ac",x"347b",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470",x"b9c6",x"404d",x"37a3",x"bbd3",x"a9fd",x"3272",x"35a4",x"3474",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9c6",x"404e",x"37b6",x"b93b",x"b9e8",x"313a",x"359f",x"346f",x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470",x"b9cd",x"404f",x"37aa",x"b9e5",x"b8ae",x"3566",x"35a5",x"346b"),
(x"b9c6",x"404e",x"37c1",x"ba55",x"b865",x"b441",x"359c",x"346e",x"b9c6",x"404e",x"37b6",x"b93b",x"b9e8",x"313a",x"359f",x"346f",x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468"),
(x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9c6",x"404e",x"37c1",x"ba55",x"b865",x"b441",x"359c",x"346e",x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477"),
(x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485"),
(x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485",x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f"),
(x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f",x"b9cb",x"403d",x"37b2",x"bbec",x"ac1f",x"2fcd",x"3595",x"349f",x"b9ca",x"4031",x"3795",x"bbe2",x"acf4",x"30cb",x"3598",x"34c3"),
(x"b9cb",x"403d",x"37b2",x"bbec",x"ac1f",x"2fcd",x"3595",x"349f",x"b9cc",x"403d",x"37a7",x"bbbc",x"2e02",x"b38e",x"3599",x"349f",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485"),
(x"b9cc",x"4045",x"37d1",x"bbf6",x"a9b5",x"2d99",x"358e",x"3485",x"b9cc",x"4046",x"37c6",x"bb50",x"30fd",x"b5fd",x"3592",x"3485",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477"),
(x"b9cc",x"404a",x"37de",x"bbe7",x"a00b",x"30f2",x"358d",x"3476",x"b9cd",x"404a",x"37d4",x"bb44",x"293f",x"b6a9",x"3590",x"3477",x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"b9cc",x"4050",x"37cc",x"bbe3",x"2d8f",x"3091",x"3598",x"3466",x"b9cc",x"404d",x"37dc",x"bbd6",x"2b52",x"322d",x"3590",x"346c",x"b9cd",x"404d",x"37d2",x"bbb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"b9cd",x"4050",x"37b8",x"bbf8",x"2c13",x"2b34",x"35a1",x"3466",x"b9cc",x"4050",x"37cc",x"bbe3",x"2d8f",x"3091",x"3598",x"3466",x"b9cd",x"404f",x"37c8",x"baa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"b9cd",x"4050",x"37a7",x"bbff",x"232b",x"2518",x"35a7",x"3469",x"b9cd",x"4050",x"37b8",x"bbf8",x"2c13",x"2b34",x"35a1",x"3466",x"b9cd",x"4050",x"37b7",x"ba3a",x"b904",x"a765",x"35a0",x"3468"),
(x"b9cd",x"4050",x"37a7",x"bbff",x"232b",x"2518",x"35a7",x"3469",x"b9cd",x"404f",x"37aa",x"b9e5",x"b8ae",x"3566",x"35a5",x"346b",x"b9cd",x"404d",x"3799",x"ba98",x"b4cf",x"37ab",x"35ab",x"3472"),
(x"b9cd",x"404a",x"3790",x"bb17",x"ade0",x"3741",x"35ac",x"347b",x"b9ce",x"404a",x"3784",x"bbd5",x"a532",x"3276",x"35b1",x"347c",x"b9ce",x"404e",x"378e",x"bbf3",x"a432",x"2ede",x"35af",x"3471"),
(x"b9ce",x"404a",x"3784",x"bbd5",x"a532",x"3276",x"35b1",x"347c",x"b9cd",x"404a",x"3790",x"bb17",x"ade0",x"3741",x"35ac",x"347b",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b"),
(x"b9cf",x"4045",x"377f",x"bbc6",x"a6c8",x"337e",x"35b0",x"348c",x"b9cd",x"4045",x"378b",x"baba",x"ab10",x"384d",x"35ab",x"348b",x"b9cd",x"403d",x"3783",x"bb8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9ca",x"403d",x"379f",x"bbf7",x"2d6b",x"a836",x"359d",x"34a0",x"b9cb",x"4031",x"378d",x"bbfd",x"1418",x"2a73",x"359b",x"34c3"),
(x"b9ca",x"403d",x"379f",x"bbf7",x"2d6b",x"a836",x"359d",x"34a0",x"b9cb",x"403d",x"378a",x"bbb7",x"a074",x"3436",x"35a4",x"34a2",x"b9c8",x"4045",x"3794",x"bbbc",x"287e",x"3408",x"35a6",x"348a"),
(x"b9c6",x"4046",x"37ba",x"bbd9",x"2f7e",x"b0f2",x"3599",x"3485",x"b9c8",x"4045",x"3794",x"bbbc",x"287e",x"3408",x"35a6",x"348a",x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c"),
(x"b9c6",x"404a",x"37c9",x"bbcb",x"2cfc",x"b2c5",x"3597",x"3478",x"b9c8",x"404a",x"3798",x"bb91",x"ab6f",x"3519",x"35a7",x"347c",x"b9c6",x"404d",x"37a3",x"bbd3",x"a9fd",x"3272",x"35a4",x"3474"),
(x"b9c6",x"404d",x"37c7",x"bb5f",x"ae12",x"b605",x"3599",x"3471",x"b9c6",x"404d",x"37a3",x"bbd3",x"a9fd",x"3272",x"35a4",x"3474",x"b9c6",x"404e",x"37ac",x"bad8",x"b658",x"3550",x"35a2",x"3470"),
(x"b9cb",x"403d",x"37b2",x"b86e",x"b47a",x"3a45",x"367a",x"29b1",x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b9ae",x"4031",x"37c0",x"1bc8",x"b48d",x"3bab",x"365d",x"2ab9"),
(x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b9cb",x"403d",x"37b2",x"b86e",x"b47a",x"3a45",x"367a",x"29b1",x"b9cc",x"4045",x"37d1",x"b856",x"b5aa",x"3a18",x"3678",x"28cc"),
(x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b9cc",x"4045",x"37d1",x"b856",x"b5aa",x"3a18",x"3678",x"28cc",x"b9cc",x"404a",x"37de",x"b892",x"b07e",x"3a77",x"3675",x"284f"),
(x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b9cc",x"404a",x"37de",x"b892",x"b07e",x"3a77",x"3675",x"284f",x"b9cc",x"404d",x"37dc",x"b809",x"374a",x"39de",x"3673",x"27ef"),
(x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e",x"b9ac",x"4050",x"37fd",x"232b",x"38f3",x"3a48",x"365b",x"2806",x"b9cc",x"404d",x"37dc",x"b809",x"374a",x"39de",x"3673",x"27ef"),
(x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709",x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e",x"b9cc",x"4050",x"37cc",x"b4ee",x"3aeb",x"3653",x"3673",x"275d"),
(x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c",x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709",x"b9cd",x"4050",x"37b8",x"b361",x"3bc7",x"282c",x"3674",x"26df"),
(x"b9c4",x"4050",x"379c",x"b458",x"3b15",x"b609",x"366f",x"2623",x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c",x"b9cd",x"4050",x"37a7",x"b362",x"3b62",x"b4ea",x"3676",x"2679"),
(x"b9d3",x"404e",x"378c",x"38cb",x"39b0",x"35e1",x"3620",x"3508",x"b9d5",x"404f",x"3782",x"385b",x"3ab4",x"a80e",x"361b",x"3507",x"b9cd",x"404e",x"3786",x"375f",x"39e5",x"37e9",x"3620",x"350c"),
(x"b9cd",x"404e",x"3786",x"b5de",x"3b08",x"34dc",x"3679",x"2599",x"b9ca",x"404e",x"378b",x"b819",x"3ad2",x"aea1",x"3676",x"25ba",x"b9ce",x"404e",x"378e",x"b62d",x"3aa4",x"b670",x"3679",x"25cc"),
(x"b95b",x"404b",x"3786",x"3ae1",x"b000",x"37eb",x"35f5",x"2dd3",x"b962",x"404f",x"378d",x"3a12",x"37fa",x"36b2",x"35f8",x"2da1",x"b956",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35e0",x"2d9e"),
(x"b962",x"404f",x"378d",x"3a12",x"37fa",x"36b2",x"35f8",x"2da1",x"b968",x"4051",x"378e",x"3610",x"3adf",x"357f",x"35fa",x"2d8a",x"b95e",x"4053",x"3752",x"3848",x"3a10",x"35f5",x"35e2",x"2d7f"),
(x"b968",x"4051",x"378e",x"3610",x"3adf",x"357f",x"35fa",x"2d8a",x"b973",x"4051",x"378f",x"a5dc",x"3bcb",x"332e",x"35fe",x"2d6c",x"b966",x"4053",x"3752",x"af69",x"3bdc",x"30a3",x"35e4",x"2d68"),
(x"b95b",x"404b",x"3786",x"3ae1",x"b000",x"37eb",x"35f5",x"2dd3",x"b94b",x"404c",x"3752",x"3ac8",x"b025",x"381c",x"35de",x"2dda",x"b962",x"403d",x"3752",x"3ab4",x"b44c",x"3799",x"35f0",x"2e8e"),
(x"b96c",x"403c",x"3775",x"3ab0",x"b345",x"37fd",x"35ff",x"2e87",x"b962",x"403d",x"3752",x"3ab4",x"b44c",x"3799",x"35f0",x"2e8e",x"b967",x"4034",x"3752",x"3aac",x"b05e",x"3846",x"35f7",x"2ef0"),
(x"b985",x"404f",x"3782",x"b861",x"3ab1",x"a386",x"3600",x"2d31",x"b966",x"4053",x"3752",x"af69",x"3bdc",x"30a3",x"35e4",x"2d68",x"b97e",x"4051",x"378e",x"b6f1",x"3b35",x"205a",x"3601",x"2d50"),
(x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b972",x"403d",x"3776",x"b31e",x"aca2",x"3bc7",x"3662",x"2cd4",x"b96c",x"403c",x"3775",x"2dad",x"b0c1",x"3be1",x"3667",x"2cd0"),
(x"b96c",x"403c",x"3775",x"2dad",x"b0c1",x"3be1",x"3667",x"2cd0",x"b972",x"403d",x"3776",x"b31e",x"aca2",x"3bc7",x"3662",x"2cd4",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83",x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8",x"b962",x"404f",x"378d",x"2f46",x"b03f",x"3be0",x"3663",x"2db2"),
(x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8",x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4",x"b968",x"4051",x"378e",x"2d5c",x"a17a",x"3bf8",x"365d",x"2dbf"),
(x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4",x"b975",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3654",x"2db4",x"b973",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3655",x"2dc0"),
(x"b973",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3655",x"2dc0",x"b975",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3654",x"2db4",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"b97e",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"364d",x"2db2",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f",x"b98c",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"3645",x"2d87",x"b987",x"404e",x"378c",x"a877",x"ae68",x"3bf4",x"3647",x"2d91"),
(x"b983",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"364c",x"2d65",x"b98c",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"b98c",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"3645",x"2d87"),
(x"b98c",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"b983",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"364c",x"2d65",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"b98b",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"364a",x"2d20",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c",x"b983",x"403d",x"3777",x"2c2f",x"afb9",x"3bec",x"3655",x"2cce"),
(x"b98c",x"403d",x"3777",x"2a04",x"ae02",x"3bf4",x"364f",x"2cc3",x"b983",x"403d",x"3777",x"2c2f",x"afb9",x"3bec",x"3655",x"2cce",x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"b983",x"403d",x"3777",x"2c2f",x"afb9",x"3bec",x"3655",x"2cce",x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"b981",x"4045",x"3780",x"3169",x"b087",x"3bcd",x"3651",x"2d2c",x"b983",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"364c",x"2d65",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68"),
(x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68",x"b983",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"364c",x"2d65",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d",x"b981",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"364c",x"2d8f",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"b977",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3654",x"2d9f",x"b97a",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3650",x"2daa",x"b975",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3654",x"2db4"),
(x"b973",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3656",x"2da5",x"b975",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3654",x"2db4",x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4"),
(x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b96c",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"365b",x"2db4",x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8"),
(x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b967",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3660",x"2da8",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b963",x"404c",x"3788",x"aed5",x"b0dc",x"3bdc",x"3665",x"2d83",x"b972",x"403d",x"3776",x"b31e",x"aca2",x"3bc7",x"3662",x"2cd4"),
(x"b979",x"4034",x"376f",x"25ae",x"abef",x"3bfb",x"3663",x"2c62",x"b985",x"4034",x"3770",x"2c25",x"ab90",x"3bf8",x"365a",x"2c5c",x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5"),
(x"b975",x"403d",x"3773",x"adae",x"ad20",x"3bf1",x"3660",x"2cd4",x"b97e",x"403e",x"3775",x"30a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"b97b",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3656",x"2d31"),
(x"b967",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3661",x"2d7d",x"b97b",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3656",x"2d31",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68"),
(x"b96a",x"404e",x"3785",x"ae64",x"b275",x"3bcb",x"365d",x"2d9b",x"b97f",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"3650",x"2d68",x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d"),
(x"b96e",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"365a",x"2da4",x"b97d",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"3650",x"2d8d",x"b977",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3654",x"2d9f"),
(x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8",x"b992",x"4045",x"3794",x"3bd9",x"292f",x"3209",x"35f5",x"33a8",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa",x"b992",x"4045",x"3794",x"3bd9",x"292f",x"3209",x"35f5",x"33a8",x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b"),
(x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b",x"b994",x"404d",x"37a3",x"3bda",x"aea9",x"311c",x"35f5",x"337c",x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377",x"b994",x"404d",x"37a3",x"3bda",x"aea9",x"311c",x"35f5",x"337c",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"b98d",x"404f",x"37aa",x"3a13",x"b891",x"34fa",x"35f4",x"336a",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373",x"b993",x"404f",x"37b7",x"3977",x"b9c7",x"2ec0",x"35fa",x"336e"),
(x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b993",x"404f",x"37b7",x"3977",x"b9c7",x"2ec0",x"35fa",x"336e",x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e"),
(x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e",x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b"),
(x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b990",x"403d",x"37a1",x"3bf5",x"2dc9",x"aa2b",x"3600",x"33d2",x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1"),
(x"b98e",x"403d",x"37a5",x"3bc3",x"2ec2",x"b2f5",x"3601",x"33d1",x"b98d",x"4030",x"378d",x"3bfe",x"28c2",x"2138",x"3602",x"340f",x"b98e",x"4030",x"3797",x"3bf6",x"a3bb",x"2e0a",x"3606",x"340f"),
(x"b98e",x"403d",x"37b0",x"3bff",x"a3ef",x"2511",x"3606",x"33d1",x"b98e",x"4045",x"37d0",x"3c00",x"9fe2",x"868d",x"360b",x"339c",x"b98e",x"4046",x"37c6",x"3b29",x"3144",x"b6a0",x"3608",x"339b"),
(x"b98e",x"4045",x"37d0",x"3c00",x"9fe2",x"868d",x"360b",x"339c",x"b98e",x"404a",x"37dc",x"3bfd",x"1481",x"a9d9",x"360c",x"337d",x"b98e",x"404a",x"37d2",x"3afe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"b98e",x"404a",x"37dc",x"3bfd",x"1481",x"a9d9",x"360c",x"337d",x"b98e",x"404d",x"37db",x"3bff",x"9018",x"a31d",x"3608",x"336a",x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"b98e",x"404d",x"37d0",x"3b62",x"afb4",x"b5d8",x"3604",x"336f",x"b98e",x"404d",x"37db",x"3bff",x"9018",x"a31d",x"3608",x"336a",x"b98e",x"4050",x"37cd",x"3bfa",x"2874",x"2c13",x"3601",x"3360"),
(x"b98d",x"404f",x"37c9",x"3b31",x"b5e3",x"b397",x"3600",x"3366",x"b98e",x"4050",x"37cd",x"3bfa",x"2874",x"2c13",x"3601",x"3360",x"b98d",x"4050",x"37b8",x"3bfa",x"2a69",x"2a66",x"35f8",x"3360"),
(x"b98d",x"404f",x"37b7",x"3a7d",x"b8a9",x"a953",x"35f9",x"3365",x"b98d",x"4050",x"37b8",x"3bfa",x"2a69",x"2a66",x"35f8",x"3360",x"b98d",x"4050",x"37a7",x"3bff",x"20dd",x"25fd",x"35f2",x"3366"),
(x"b98d",x"4050",x"37a7",x"3bff",x"20dd",x"25fd",x"35f2",x"3366",x"b98d",x"404e",x"378e",x"3bf3",x"a432",x"2f1d",x"35ea",x"3376",x"b98d",x"404d",x"3798",x"3a9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"b98d",x"404e",x"378e",x"3bf3",x"a432",x"2f1d",x"35ea",x"3376",x"b98c",x"404a",x"3784",x"3bd5",x"a532",x"3276",x"35e9",x"338d",x"b98d",x"404a",x"3790",x"3b10",x"ad8c",x"3760",x"35ed",x"338b"),
(x"b98c",x"404a",x"3784",x"3bd5",x"a532",x"3276",x"35e9",x"338d",x"b98b",x"4045",x"377f",x"3bc5",x"a6cf",x"3387",x"35eb",x"33ac",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"b98d",x"403d",x"3782",x"3b88",x"abb1",x"354b",x"35f4",x"33d9",x"b98d",x"4045",x"378b",x"3abf",x"ab14",x"3846",x"35ef",x"33aa",x"b98b",x"4045",x"377f",x"3bc5",x"a6cf",x"3387",x"35eb",x"33ac"),
(x"b98d",x"4030",x"378d",x"3bfe",x"28c2",x"2138",x"3602",x"340f",x"b990",x"403d",x"37a1",x"3bf5",x"2dc9",x"aa2b",x"3600",x"33d2",x"b98f",x"403d",x"378a",x"3bd9",x"243f",x"3220",x"35f7",x"33d8"),
(x"b990",x"403d",x"37a1",x"3bf5",x"2dc9",x"aa2b",x"3600",x"33d2",x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b992",x"4045",x"3794",x"3bd9",x"292f",x"3209",x"35f5",x"33a8"),
(x"b993",x"4046",x"37be",x"3bdb",x"2f8d",x"b0af",x"3602",x"339b",x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b992",x"404a",x"3798",x"3ba3",x"a849",x"34bc",x"35f2",x"338b"),
(x"b994",x"404a",x"37c9",x"3bce",x"2c74",x"b2a7",x"3603",x"3383",x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b994",x"404d",x"37a3",x"3bda",x"aea9",x"311c",x"35f5",x"337c"),
(x"b993",x"404d",x"37c9",x"3b8e",x"aeae",x"b4f9",x"3601",x"3374",x"b993",x"404e",x"37c3",x"3a5f",x"b7e4",x"b595",x"35fe",x"336e",x"b993",x"404e",x"37ac",x"3b0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"b9ae",x"4031",x"37c0",x"1bc8",x"b48d",x"3bab",x"365d",x"2ab9",x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b98e",x"403d",x"37b0",x"3860",x"b445",x"3a59",x"363e",x"29b6"),
(x"b9ac",x"403d",x"37dc",x"21d6",x"b62a",x"3b61",x"365c",x"298f",x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b98e",x"4045",x"37d0",x"386c",x"b560",x"3a19",x"3640",x"28d0"),
(x"b9ae",x"4046",x"3800",x"22cf",x"b59c",x"3b7d",x"365c",x"28a9",x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b98e",x"404a",x"37dc",x"3889",x"b0d3",x"3a7a",x"3643",x"2852"),
(x"b9ad",x"404b",x"3804",x"2194",x"2bfc",x"3bfb",x"365c",x"284f",x"b9ac",x"4050",x"37fd",x"232b",x"38f3",x"3a48",x"365b",x"2806",x"b98e",x"404d",x"37db",x"3837",x"36a0",x"39ef",x"3644",x"2800"),
(x"b98e",x"404d",x"37db",x"3837",x"36a0",x"39ef",x"3644",x"2800",x"b9ac",x"4050",x"37fd",x"232b",x"38f3",x"3a48",x"365b",x"2806",x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e"),
(x"b98e",x"4050",x"37cd",x"3534",x"3ad6",x"367a",x"3644",x"2773",x"b9ac",x"4051",x"37e2",x"1bc8",x"3b01",x"37bb",x"365b",x"278e",x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709"),
(x"b98d",x"4050",x"37b8",x"33c4",x"3bc1",x"28ed",x"3642",x"26f2",x"b9ac",x"4052",x"37c9",x"1881",x"3be6",x"3101",x"365b",x"2709",x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c"),
(x"b98d",x"4050",x"37a7",x"342d",x"3b51",x"b4ec",x"3641",x"268d",x"b9ac",x"4052",x"37b3",x"275f",x"3bdf",x"b19a",x"365b",x"268c",x"b995",x"404f",x"3789",x"3469",x"3b25",x"b5af",x"3644",x"25c3"),
(x"b98e",x"404e",x"3782",x"b7c9",x"39ef",x"375f",x"3603",x"2d14",x"b985",x"404f",x"3782",x"b861",x"3ab1",x"a386",x"3600",x"2d31",x"b987",x"404e",x"378c",x"b8b4",x"39be",x"35f4",x"3605",x"2d2d"),
(x"b990",x"404e",x"378b",x"3682",x"3b4c",x"2987",x"363f",x"25d0",x"b98e",x"404e",x"3782",x"35ed",x"3b6c",x"2991",x"363e",x"2598",x"b98c",x"404e",x"378b",x"35f3",x"3b61",x"2ea6",x"363c",x"25cf"),
(x"b967",x"4034",x"3752",x"3aac",x"b05e",x"3846",x"35f7",x"2ef0",x"b96d",x"402c",x"3752",x"3ada",x"b039",x"37f9",x"35fe",x"2f4f",x"b972",x"4030",x"376e",x"3ab7",x"ada6",x"384a",x"3606",x"2f15"),
(x"b972",x"4033",x"376d",x"303b",x"ac06",x"3be9",x"3668",x"2c64",x"b972",x"4030",x"376e",x"312d",x"2310",x"3be4",x"366a",x"2c3f",x"b97b",x"4032",x"3770",x"2cfa",x"29bc",x"3bf7",x"3663",x"2c4b"),
(x"b9e6",x"402f",x"376e",x"bafb",x"ad7a",x"37ae",x"3622",x"348b",x"b9ec",x"402b",x"3752",x"baff",x"adb0",x"379f",x"3619",x"347e",x"b9f0",x"4034",x"3752",x"bafe",x"b17b",x"3746",x"3612",x"3497"),
(x"b9e1",x"4034",x"376f",x"a7bb",x"a9c9",x"3bfc",x"3609",x"333a",x"b9d5",x"4034",x"3770",x"ac95",x"ac08",x"3bf6",x"3600",x"333b",x"b9d5",x"4031",x"3770",x"a935",x"1ec2",x"3bfe",x"3601",x"3350"),
(x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5",x"3ac5",x"4000",x"377d",x"35fa",x"3ae9",x"3563",x"3641",x"34e8",x"3ac6",x"3ffd",x"3794",x"3663",x"3a38",x"37c6",x"363b",x"34f0"),
(x"3acf",x"3ffd",x"377a",x"3866",x"3a42",x"34ab",x"3647",x"34ee",x"3ac5",x"4000",x"377d",x"35fa",x"3ae9",x"3563",x"3641",x"34e8",x"3acb",x"4001",x"3752",x"324e",x"3bb3",x"31e9",x"364f",x"34df"),
(x"3acf",x"3ffd",x"377a",x"3068",x"a815",x"3beb",x"35ed",x"20c2",x"3ac4",x"3ff5",x"377c",x"3068",x"a815",x"3beb",x"35f4",x"1e8d",x"3ac5",x"4000",x"377d",x"3068",x"a815",x"3beb",x"35f4",x"2148"),
(x"3ac6",x"3ffd",x"3794",x"3be8",x"aaec",x"b08c",x"35fb",x"305f",x"3ac5",x"4000",x"377d",x"3be8",x"aaec",x"b08c",x"35fb",x"3073",x"3ac4",x"3ff5",x"377c",x"3be8",x"aaec",x"b08c",x"35ed",x"3063"),
(x"3acf",x"3ffd",x"377a",x"3a72",x"b86b",x"32c9",x"3669",x"31b3",x"3ad6",x"3ffe",x"3752",x"3a94",x"b7fc",x"345d",x"365a",x"31b1",x"3ac4",x"3ff5",x"377c",x"39d9",x"b836",x"36f0",x"366f",x"3198"),
(x"3a98",x"3fdf",x"3787",x"38c1",x"b811",x"38fb",x"3686",x"3146",x"3ab4",x"3ffc",x"37b2",x"38ae",x"b826",x"38fc",x"3686",x"31ae",x"3abb",x"3fec",x"376e",x"38f8",x"b816",x"38c1",x"366f",x"3179"),
(x"3ab4",x"3ffc",x"37b2",x"b422",x"b30f",x"3b86",x"3632",x"2b49",x"3a98",x"3fdf",x"3787",x"b776",x"b053",x"3afe",x"3632",x"2c6d",x"3aaa",x"3ffd",x"37ae",x"b776",x"b054",x"3afe",x"362b",x"2b5e"),
(x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5",x"3ab4",x"3ffc",x"37b2",x"348b",x"3a04",x"38c2",x"362a",x"34ed",x"3aaa",x"3ffd",x"37ae",x"b35d",x"39d9",x"3923",x"3626",x"34e7"),
(x"3aaa",x"3ffd",x"37ae",x"b776",x"b054",x"3afe",x"362b",x"2b5e",x"3a98",x"3fdf",x"3787",x"b776",x"b053",x"3afe",x"3632",x"2c6d",x"3aa1",x"3ffe",x"379f",x"b8fe",x"ab38",x"3a3b",x"3623",x"2b7a"),
(x"3aa1",x"3ffe",x"379f",x"b54f",x"39c9",x"38d8",x"3624",x"34df",x"3a94",x"4000",x"3780",x"acbe",x"3bc6",x"3329",x"3626",x"34ce",x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"3aad",x"4001",x"3752",x"1da1",x"3bf5",x"2e87",x"3640",x"34ce",x"3acb",x"4001",x"3752",x"324e",x"3bb3",x"31e9",x"364f",x"34df",x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5",x"3acb",x"4001",x"3752",x"324e",x"3bb3",x"31e9",x"364f",x"34df",x"3ac5",x"4000",x"377d",x"35fa",x"3ae9",x"3563",x"3641",x"34e8"),
(x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e",x"3a81",x"3fff",x"37ca",x"2393",x"3b79",x"35b2",x"362a",x"2f26",x"3a78",x"3ffc",x"37d9",x"b146",x"3a67",x"389c",x"3623",x"2f40"),
(x"3a81",x"3fff",x"37ca",x"2393",x"3b79",x"35b2",x"362a",x"2f26",x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3a9b",x"3ffd",x"37d0",x"31ec",x"3b16",x"36cd",x"363e",x"2f34"),
(x"3a89",x"3ffd",x"37d9",x"b950",x"a0ea",x"39fa",x"35f6",x"208e",x"3a81",x"3ff6",x"37ca",x"b950",x"a0ea",x"39fa",x"35fe",x"1e8d",x"3a81",x"3fff",x"37ca",x"b950",x"a0ea",x"39fa",x"35fe",x"210b"),
(x"3a78",x"3ffc",x"37d9",x"393c",x"95bc",x"3a0c",x"35df",x"2d1a",x"3a81",x"3fff",x"37ca",x"393c",x"95bc",x"3a0c",x"35e8",x"2d07",x"3a81",x"3ff6",x"37ca",x"393c",x"95bc",x"3a0c",x"35e8",x"2d3f"),
(x"3a89",x"3ffd",x"37d9",x"3325",x"b878",x"3a63",x"3671",x"322e",x"3a9b",x"3ffd",x"37d0",x"333b",x"b811",x"3aa5",x"367e",x"322f",x"3a81",x"3ff6",x"37ca",x"9e0a",x"b823",x"3ad8",x"366b",x"3246"),
(x"3a65",x"3fe3",x"3791",x"b252",x"b816",x"3ab1",x"3657",x"328b",x"3a63",x"3ffc",x"37cd",x"b1e7",x"b81a",x"3ab5",x"3654",x"3237",x"3a81",x"3fe8",x"37ad",x"23bb",x"b81b",x"3add",x"366c",x"3272"),
(x"3a63",x"3ffc",x"37cd",x"baf6",x"b475",x"367c",x"35a3",x"3029",x"3a65",x"3fe3",x"3791",x"bae1",x"b415",x"370f",x"35b4",x"2fb8",x"3a5e",x"3ffc",x"37ba",x"bb3a",x"b41e",x"357a",x"35ab",x"3028"),
(x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e",x"3a63",x"3ffc",x"37cd",x"b58a",x"3a1b",x"385c",x"3613",x"2f2b",x"3a5e",x"3ffc",x"37ba",x"b926",x"39b7",x"3464",x"360f",x"2f0f"),
(x"3a5e",x"3ffc",x"37ba",x"bb3a",x"b41e",x"357a",x"35ab",x"3028",x"3a65",x"3fe3",x"3791",x"bae1",x"b415",x"370f",x"35b4",x"2fb8",x"3a59",x"3ffc",x"379b",x"bad4",x"b3bd",x"3761",x"35b7",x"3027"),
(x"3a59",x"3ffc",x"379b",x"b825",x"3acf",x"2d30",x"360b",x"2ee1",x"3a66",x"3fff",x"3781",x"b1af",x"3bdf",x"1c18",x"3615",x"2eb7",x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"3a94",x"4000",x"3780",x"16f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e",x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3a81",x"3fff",x"37ca",x"2393",x"3b79",x"35b2",x"362a",x"2f26"),
(x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3a94",x"4000",x"3780",x"16f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"3aa1",x"3ffe",x"379f",x"394b",x"39eb",x"af9c",x"3644",x"2eeb"),
(x"3a9b",x"3ffd",x"37d0",x"31ec",x"3b16",x"36cd",x"363e",x"2f34",x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3aa3",x"3ffd",x"37ba",x"392f",x"39d8",x"32de",x"3644",x"2f14"),
(x"3a9b",x"3ffd",x"37d0",x"39f1",x"b5fe",x"3870",x"3609",x"314d",x"3aa3",x"3ffd",x"37ba",x"3b76",x"b463",x"3373",x"35ff",x"3145",x"3a98",x"3fdf",x"3787",x"3b76",x"b463",x"3373",x"3609",x"30e6"),
(x"3aa1",x"3ffe",x"379f",x"3bda",x"afe2",x"b0aa",x"35f6",x"313b",x"3a98",x"3fdf",x"3787",x"3b76",x"b463",x"3373",x"3609",x"30e6",x"3aa3",x"3ffd",x"37ba",x"3b76",x"b463",x"3373",x"35ff",x"3145"),
(x"3a61",x"3fe3",x"378f",x"b45c",x"b0de",x"3b99",x"35b7",x"2fb9",x"3a59",x"3ffc",x"379b",x"bad4",x"b3bd",x"3760",x"35b7",x"3027",x"3a65",x"3fe3",x"3791",x"bae1",x"b415",x"370f",x"35b4",x"2fb8"),
(x"3a59",x"3ffc",x"379b",x"366b",x"ac20",x"3b4f",x"369d",x"307f",x"3a61",x"3fe3",x"378f",x"28e0",x"aefd",x"3bf2",x"369d",x"30c9",x"3a5f",x"3fdf",x"378e",x"b496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"3a3c",x"3fec",x"376e",x"b931",x"b7c9",x"38ad",x"367c",x"30b4",x"3a44",x"3ffc",x"37af",x"b5ad",x"b6ed",x"3aa0",x"368c",x"3079",x"3a5f",x"3fdf",x"378e",x"b496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"3a44",x"3ffc",x"37af",x"b5ad",x"b6ed",x"3aa0",x"368c",x"3079",x"3a33",x"3ff5",x"377b",x"b9d9",x"b840",x"36d9",x"3678",x"3096",x"3a31",x"3ffb",x"378b",x"b815",x"b8b5",x"3904",x"3679",x"3081"),
(x"3a28",x"3ffd",x"3775",x"ba73",x"b85c",x"3350",x"366e",x"3082",x"3a33",x"3ff5",x"377b",x"b9d9",x"b840",x"36d9",x"3678",x"3096",x"3a22",x"3ffe",x"3752",x"ba86",x"b81f",x"3433",x"3660",x"3089"),
(x"3a33",x"4000",x"3780",x"bbd2",x"3047",x"b133",x"35cc",x"200a",x"3a33",x"3ffd",x"3797",x"bb81",x"34c0",x"31b8",x"35cc",x"214e",x"3a31",x"3ffb",x"378b",x"bbd2",x"3047",x"b133",x"35c7",x"210d"),
(x"3a33",x"4000",x"3780",x"b66b",x"ad14",x"3b4c",x"35d6",x"1e80",x"3a33",x"3ff5",x"377b",x"b612",x"af46",x"3b58",x"35d6",x"214e",x"3a28",x"3ffd",x"3775",x"b66c",x"ad14",x"3b4c",x"35cd",x"1ffb"),
(x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec",x"3a44",x"3ffc",x"37af",x"9fc8",x"3964",x"39e8",x"35ca",x"32fc",x"3a33",x"3ffd",x"3797",x"b553",x"3a2a",x"3859",x"35bc",x"3307"),
(x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec",x"3a60",x"4001",x"3777",x"3179",x"3b46",x"3611",x"35c7",x"32bf",x"3a59",x"3ffc",x"379b",x"35ee",x"392f",x"3951",x"35d0",x"32dc"),
(x"3a59",x"3ffc",x"379b",x"35ee",x"392f",x"3951",x"35d0",x"32dc",x"3a60",x"4001",x"3777",x"3179",x"3b46",x"3611",x"35c7",x"32bf",x"3a66",x"3fff",x"3781",x"3106",x"3a66",x"38a1",x"35cd",x"32bf"),
(x"3a56",x"4001",x"375e",x"a8c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"3a60",x"4001",x"3777",x"3179",x"3b46",x"3611",x"35c7",x"32bf",x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec"),
(x"3a2b",x"4001",x"3752",x"b411",x"3b93",x"3249",x"35a3",x"32ec",x"3a2b",x"3fff",x"3777",x"b91c",x"39e9",x"32d4",x"35ae",x"32ff",x"3a28",x"3ffd",x"3775",x"b9ba",x"391c",x"347b",x"35ab",x"3307"),
(x"3a51",x"4001",x"3752",x"a4f0",x"3bea",x"309d",x"35b4",x"32bf",x"3a56",x"4001",x"375e",x"a8c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"3a33",x"4000",x"3780",x"ade0",x"3bd5",x"31bf",x"35b4",x"32f9"),
(x"3a33",x"4000",x"3780",x"ade0",x"3bd5",x"31bf",x"35b4",x"32f9",x"3a2b",x"3fff",x"3777",x"b91c",x"39e9",x"32d4",x"35ae",x"32ff",x"3a2b",x"4001",x"3752",x"b411",x"3b93",x"3249",x"35a3",x"32ec"),
(x"3ab4",x"3ffc",x"37b2",x"348b",x"3a04",x"38c2",x"362a",x"34ed",x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5",x"3ac6",x"3ffd",x"3794",x"3663",x"3a38",x"37c6",x"363b",x"34f0"),
(x"3ad6",x"3ffe",x"3752",x"3892",x"3a2a",x"3480",x"3655",x"34e7",x"3acf",x"3ffd",x"377a",x"3866",x"3a42",x"34ab",x"3647",x"34ee",x"3acb",x"4001",x"3752",x"324e",x"3bb3",x"31e9",x"364f",x"34df"),
(x"3ac3",x"3fee",x"3752",x"3a96",x"b7a7",x"34e2",x"3663",x"317c",x"3ac4",x"3ff5",x"377c",x"39d9",x"b836",x"36f0",x"366f",x"3198",x"3ad6",x"3ffe",x"3752",x"3a94",x"b7fc",x"345d",x"365a",x"31b1"),
(x"3abb",x"3fec",x"376e",x"38f8",x"b816",x"38c1",x"366f",x"3179",x"3ac4",x"3ff5",x"377c",x"39d9",x"b836",x"36f0",x"366f",x"3198",x"3ac3",x"3fee",x"3752",x"3a96",x"b7a7",x"34e2",x"3663",x"317c"),
(x"3ac4",x"3ff5",x"377c",x"39d9",x"b836",x"36f0",x"366f",x"3198",x"3ab4",x"3ffc",x"37b2",x"38ae",x"b826",x"38fc",x"3686",x"31ae",x"3ac6",x"3ffd",x"3794",x"3839",x"b89f",x"38fa",x"3675",x"31b3"),
(x"3abb",x"3fec",x"376e",x"38f8",x"b816",x"38c1",x"366f",x"3179",x"3ab4",x"3ffc",x"37b2",x"38ae",x"b826",x"38fc",x"3686",x"31ae",x"3ac4",x"3ff5",x"377c",x"39d9",x"b836",x"36f0",x"366f",x"3198"),
(x"3aaa",x"3ffd",x"37ae",x"b35d",x"39d9",x"3923",x"3626",x"34e7",x"3aa1",x"3ffe",x"379f",x"b54f",x"39c9",x"38d8",x"3624",x"34df",x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"3a94",x"4000",x"3780",x"acbf",x"3bc6",x"3329",x"3626",x"34ce",x"3aad",x"4001",x"3752",x"1da1",x"3bf5",x"2e87",x"3640",x"34ce",x"3aaf",x"4000",x"37a1",x"2b52",x"3bb2",x"3444",x"362d",x"34e5"),
(x"3a63",x"3ffc",x"37cd",x"b58a",x"3a1b",x"385c",x"3613",x"2f2b",x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e",x"3a78",x"3ffc",x"37d9",x"b146",x"3a67",x"389c",x"3623",x"2f40"),
(x"3a89",x"3ffd",x"37d9",x"2e09",x"3b05",x"3784",x"3631",x"2f41",x"3a81",x"3fff",x"37ca",x"2393",x"3b79",x"35b2",x"362a",x"2f26",x"3a9b",x"3ffd",x"37d0",x"31ec",x"3b16",x"36cd",x"363e",x"2f34"),
(x"3a98",x"3fdf",x"3787",x"3409",x"b819",x"3a90",x"367e",x"3296",x"3a81",x"3fe8",x"37ad",x"23bb",x"b81b",x"3add",x"366c",x"3272",x"3a9b",x"3ffd",x"37d0",x"333b",x"b811",x"3aa5",x"367e",x"322f"),
(x"3a81",x"3ff6",x"37ca",x"9e0a",x"b823",x"3ad8",x"366b",x"3246",x"3a9b",x"3ffd",x"37d0",x"333b",x"b811",x"3aa5",x"367e",x"322f",x"3a81",x"3fe8",x"37ad",x"23bb",x"b81b",x"3add",x"366c",x"3272"),
(x"3a81",x"3ff6",x"37ca",x"9e0a",x"b823",x"3ad8",x"366b",x"3246",x"3a63",x"3ffc",x"37cd",x"b1e7",x"b81a",x"3ab5",x"3654",x"3237",x"3a78",x"3ffc",x"37d9",x"b24d",x"b8ad",x"3a4b",x"3664",x"3230"),
(x"3a81",x"3fe8",x"37ad",x"23bb",x"b81b",x"3add",x"366c",x"3272",x"3a63",x"3ffc",x"37cd",x"b1e7",x"b81a",x"3ab5",x"3654",x"3237",x"3a81",x"3ff6",x"37ca",x"9e0a",x"b823",x"3ad8",x"366b",x"3246"),
(x"3a5e",x"3ffc",x"37ba",x"b926",x"39b7",x"3464",x"360f",x"2f0f",x"3a59",x"3ffc",x"379b",x"b825",x"3acf",x"2d30",x"360b",x"2ee1",x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"3a66",x"3fff",x"3781",x"b1af",x"3bdf",x"1c18",x"3615",x"2eb7",x"3a94",x"4000",x"3780",x"16f6",x"3bfe",x"27c1",x"3638",x"2eb7",x"3a67",x"4000",x"37bc",x"b0a0",x"3bd5",x"3081",x"3618",x"2f0e"),
(x"3aa3",x"3ffd",x"37ba",x"392f",x"39d8",x"32de",x"3644",x"2f14",x"3a9d",x"4000",x"37b1",x"2f93",x"3bda",x"30c0",x"363e",x"2f02",x"3aa1",x"3ffe",x"379f",x"394b",x"39eb",x"af9c",x"3644",x"2eeb"),
(x"3a44",x"3ffc",x"37af",x"b5ad",x"b6ed",x"3aa0",x"368c",x"3079",x"3a59",x"3ffc",x"379b",x"366b",x"ac20",x"3b4f",x"369d",x"307f",x"3a5f",x"3fdf",x"378e",x"b496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"3a59",x"3fdf",x"377f",x"b92b",x"b842",x"385f",x"3694",x"30d7",x"3a3c",x"3fec",x"376e",x"b931",x"b7c9",x"38ad",x"367c",x"30b4",x"3a5f",x"3fdf",x"378e",x"b496",x"b62e",x"3b03",x"369b",x"30d4"),
(x"3a44",x"3ffc",x"37af",x"b5ad",x"b6ed",x"3aa0",x"368c",x"3079",x"3a31",x"3ffb",x"378b",x"b815",x"b8b5",x"3904",x"3679",x"3081",x"3a33",x"3ffd",x"3797",x"b810",x"b8bd",x"3900",x"367c",x"3079"),
(x"3a3c",x"3fec",x"376e",x"b931",x"b7c9",x"38ad",x"367c",x"30b4",x"3a33",x"3ff5",x"377b",x"b9d9",x"b840",x"36d9",x"3678",x"3096",x"3a44",x"3ffc",x"37af",x"b5ad",x"b6ed",x"3aa0",x"368c",x"3079"),
(x"3a36",x"3fee",x"3752",x"ba94",x"b7fd",x"345a",x"3671",x"30b8",x"3a33",x"3ff5",x"377b",x"b9d9",x"b840",x"36d9",x"3678",x"3096",x"3a3c",x"3fec",x"376e",x"b931",x"b7c9",x"38ad",x"367c",x"30b4"),
(x"3a22",x"3ffe",x"3752",x"ba86",x"b81f",x"3433",x"3660",x"3089",x"3a33",x"3ff5",x"377b",x"b9d9",x"b840",x"36d9",x"3678",x"3096",x"3a36",x"3fee",x"3752",x"ba94",x"b7fd",x"345a",x"3671",x"30b8"),
(x"3a33",x"3ff5",x"377b",x"bb82",x"286a",x"b57a",x"35bc",x"20d5",x"3a33",x"4000",x"3780",x"bbd2",x"3047",x"b133",x"35cc",x"200a",x"3a31",x"3ffb",x"378b",x"bbd2",x"3047",x"b133",x"35c7",x"210d"),
(x"3a2b",x"3fff",x"3777",x"b827",x"3037",x"3ac1",x"35cf",x"1efe",x"3a33",x"4000",x"3780",x"b66b",x"ad14",x"3b4c",x"35d6",x"1e80",x"3a28",x"3ffd",x"3775",x"b66c",x"ad14",x"3b4c",x"35cd",x"1ffb"),
(x"3a33",x"4000",x"3780",x"ade0",x"3bd5",x"31bf",x"35b4",x"32f9",x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec",x"3a33",x"3ffd",x"3797",x"b553",x"3a2a",x"3859",x"35bc",x"3307"),
(x"3a44",x"3ffc",x"37af",x"9fc8",x"3964",x"39e8",x"35ca",x"32fc",x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec",x"3a59",x"3ffc",x"379b",x"35ee",x"392f",x"3951",x"35d0",x"32dc"),
(x"3a33",x"4000",x"3780",x"ade0",x"3bd5",x"31bf",x"35b4",x"32f9",x"3a56",x"4001",x"375e",x"a8c6",x"3bf3",x"2e87",x"35ba",x"32bf",x"3a49",x"4000",x"37a0",x"90ea",x"3b79",x"35b5",x"35c6",x"32ec"),
(x"3a22",x"3ffe",x"3752",x"b8cb",x"39c5",x"358d",x"359e",x"32fc",x"3a2b",x"4001",x"3752",x"b411",x"3b93",x"3249",x"35a3",x"32ec",x"3a28",x"3ffd",x"3775",x"b9ba",x"391c",x"347b",x"35ab",x"3307"),
(x"3a2b",x"4001",x"3752",x"b411",x"3b93",x"3249",x"35a3",x"32ec",x"3a51",x"4001",x"3752",x"a4f0",x"3bea",x"309d",x"35b4",x"32bf",x"3a33",x"4000",x"3780",x"ade0",x"3bd5",x"31bf",x"35b4",x"32f9"),
(x"3aae",x"3ce9",x"376e",x"3bb7",x"8000",x"b434",x"3277",x"3554",x"3aae",x"1ef5",x"376e",x"3b33",x"0000",x"b6f8",x"3276",x"21dd",x"3ab0",x"22af",x"3794",x"3bff",x"0000",x"a460",x"32a3",x"2363"),
(x"3ab0",x"3ce9",x"3794",x"3bfe",x"8000",x"27ef",x"32a6",x"3554",x"3ab0",x"22af",x"3794",x"3bff",x"0000",x"a460",x"32a3",x"2363",x"3aad",x"2680",x"37e5",x"3be2",x"0000",x"315e",x"32d0",x"2479"),
(x"3aad",x"3ce9",x"37e5",x"3b99",x"8000",x"34ff",x"32d4",x"3554",x"3aad",x"2680",x"37e5",x"3be2",x"0000",x"315e",x"32d0",x"2479",x"3aa1",x"2805",x"3807",x"3a4b",x"8000",x"38f0",x"3301",x"253c"),
(x"3aa1",x"3ce9",x"3807",x"3970",x"0000",x"39dd",x"3302",x"3554",x"3aa1",x"2805",x"3807",x"3a4b",x"8000",x"38f0",x"3301",x"253c",x"3a90",x"2869",x"3813",x"368f",x"0000",x"3b4b",x"332f",x"25a6"),
(x"3a90",x"3ce9",x"3813",x"34a7",x"0000",x"3ba7",x"3330",x"3555",x"3a90",x"2869",x"3813",x"368f",x"0000",x"3b4b",x"332f",x"25a6",x"3a76",x"28ad",x"3818",x"a495",x"0000",x"3bff",x"335d",x"25cb"),
(x"3a5e",x"3ce9",x"3812",x"b61b",x"0000",x"3b64",x"338c",x"3555",x"3a76",x"3ce9",x"3818",x"a495",x"0000",x"3bff",x"335e",x"3555",x"3a76",x"28ad",x"3818",x"a495",x"0000",x"3bff",x"335d",x"25cb"),
(x"3a4b",x"3ce9",x"3802",x"b9c4",x"868d",x"398b",x"33ba",x"3554",x"3a5e",x"3ce9",x"3812",x"b61b",x"0000",x"3b64",x"338c",x"3555",x"3a5e",x"2870",x"3812",x"b81e",x"0000",x"3adb",x"338b",x"2594"),
(x"3a43",x"3ce9",x"37e4",x"bb9c",x"0000",x"34ef",x"33e9",x"3554",x"3a4b",x"3ce9",x"3802",x"b9c4",x"868d",x"398b",x"33ba",x"3554",x"3a4b",x"27a4",x"3802",x"ba87",x"8000",x"389f",x"33b9",x"2503"),
(x"3a41",x"3ce9",x"37ba",x"bbfc",x"0000",x"2bdf",x"340b",x"3554",x"3a43",x"3ce9",x"37e4",x"bb9c",x"0000",x"34ef",x"33e9",x"3554",x"3a43",x"2661",x"37e4",x"bbd4",x"8000",x"328e",x"33e7",x"2438"),
(x"3a41",x"3ce9",x"3775",x"bbfd",x"068d",x"aac8",x"3423",x"3554",x"3a41",x"3ce9",x"37ba",x"bbfc",x"0000",x"2bdf",x"340b",x"3554",x"3a41",x"24c7",x"37ba",x"bbff",x"0000",x"26a1",x"340b",x"22bc"),
(x"3a45",x"3ce9",x"3764",x"baa9",x"0000",x"b86d",x"343b",x"3554",x"3a41",x"3ce9",x"3775",x"bbfd",x"068d",x"aac8",x"3423",x"3554",x"3a41",x"2065",x"3775",x"bbe7",x"0000",x"b0fd",x"3423",x"2104"),
(x"3a4e",x"3ce9",x"3752",x"b98d",x"8000",x"b9c2",x"3453",x"3554",x"3a45",x"3ce9",x"3764",x"baa9",x"0000",x"b86d",x"343b",x"3554",x"3a45",x"1d1b",x"3764",x"ba17",x"0000",x"b92f",x"343b",x"1d79"),
(x"3aa3",x"3ce9",x"3752",x"3a65",x"8000",x"b8cd",x"3248",x"3554",x"3aa3",x"1a08",x"3752",x"3a65",x"8000",x"b8cd",x"3245",x"207d",x"3aae",x"1ef5",x"376e",x"3b33",x"0000",x"b6f8",x"3276",x"21dd"),
(x"3a4b",x"27a4",x"3802",x"a352",x"bab1",x"3860",x"35fb",x"3474",x"3a5e",x"2870",x"3812",x"19bc",x"bac2",x"3846",x"35ed",x"3482",x"3a76",x"28ad",x"3818",x"a495",x"ba9b",x"3881",x"35db",x"3487"),
(x"3a45",x"1d1b",x"3764",x"0a8d",x"baca",x"383a",x"35fd",x"342e",x"3aae",x"1ef5",x"376e",x"9c81",x"baa0",x"387b",x"35af",x"3433",x"3aa3",x"1a08",x"3752",x"1a24",x"bb18",x"3761",x"35b6",x"3427"),
(x"3aae",x"1ef5",x"376e",x"9c81",x"baa0",x"387b",x"35af",x"3433",x"3a45",x"1d1b",x"3764",x"0a8d",x"baca",x"383a",x"35fd",x"342e",x"3a41",x"2065",x"3775",x"9da1",x"bab0",x"3862",x"3600",x"3436"),
(x"3ab0",x"22af",x"3794",x"9953",x"bac8",x"383d",x"35ae",x"3444",x"3a41",x"2065",x"3775",x"9da1",x"bab0",x"3862",x"3600",x"3436",x"3a41",x"24c7",x"37ba",x"128d",x"bad3",x"382c",x"3601",x"3454"),
(x"3aad",x"2680",x"37e5",x"1af6",x"bad3",x"382b",x"35b1",x"3467",x"3a41",x"24c7",x"37ba",x"128d",x"bad3",x"382c",x"3601",x"3454",x"3a43",x"2661",x"37e4",x"1b5f",x"badf",x"3817",x"3600",x"3466"),
(x"3a43",x"2661",x"37e4",x"1b5f",x"badf",x"3817",x"3600",x"3466",x"3a4b",x"27a4",x"3802",x"a352",x"bab1",x"3860",x"35fb",x"3474",x"3a90",x"2869",x"3813",x"9e3f",x"bacb",x"3838",x"35c8",x"3482"),
(x"3ab0",x"3ce9",x"3794",x"3bfe",x"8000",x"27ef",x"32a6",x"3554",x"3aae",x"3ce9",x"376e",x"3bb7",x"8000",x"b434",x"3277",x"3554",x"3ab0",x"22af",x"3794",x"3bff",x"0000",x"a460",x"32a3",x"2363"),
(x"3aad",x"3ce9",x"37e5",x"3b99",x"8000",x"34ff",x"32d4",x"3554",x"3ab0",x"3ce9",x"3794",x"3bfe",x"8000",x"27ef",x"32a6",x"3554",x"3aad",x"2680",x"37e5",x"3be2",x"0000",x"315e",x"32d0",x"2479"),
(x"3aa1",x"3ce9",x"3807",x"3970",x"0000",x"39dd",x"3302",x"3554",x"3aad",x"3ce9",x"37e5",x"3b99",x"8000",x"34ff",x"32d4",x"3554",x"3aa1",x"2805",x"3807",x"3a4b",x"8000",x"38f0",x"3301",x"253c"),
(x"3a90",x"3ce9",x"3813",x"34a7",x"0000",x"3ba7",x"3330",x"3555",x"3aa1",x"3ce9",x"3807",x"3970",x"0000",x"39dd",x"3302",x"3554",x"3a90",x"2869",x"3813",x"368f",x"0000",x"3b4b",x"332f",x"25a6"),
(x"3a76",x"3ce9",x"3818",x"a495",x"0000",x"3bff",x"335e",x"3555",x"3a90",x"3ce9",x"3813",x"34a7",x"0000",x"3ba7",x"3330",x"3555",x"3a76",x"28ad",x"3818",x"a495",x"0000",x"3bff",x"335d",x"25cb"),
(x"3a5e",x"2870",x"3812",x"b81e",x"0000",x"3adb",x"338b",x"2594",x"3a5e",x"3ce9",x"3812",x"b61b",x"0000",x"3b64",x"338c",x"3555",x"3a76",x"28ad",x"3818",x"a495",x"0000",x"3bff",x"335d",x"25cb"),
(x"3a4b",x"27a4",x"3802",x"ba87",x"8000",x"389f",x"33b9",x"2503",x"3a4b",x"3ce9",x"3802",x"b9c4",x"868d",x"398b",x"33ba",x"3554",x"3a5e",x"2870",x"3812",x"b81e",x"0000",x"3adb",x"338b",x"2594"),
(x"3a43",x"2661",x"37e4",x"bbd4",x"8000",x"328e",x"33e7",x"2438",x"3a43",x"3ce9",x"37e4",x"bb9c",x"0000",x"34ef",x"33e9",x"3554",x"3a4b",x"27a4",x"3802",x"ba87",x"8000",x"389f",x"33b9",x"2503"),
(x"3a41",x"24c7",x"37ba",x"bbff",x"0000",x"26a1",x"340b",x"22bc",x"3a41",x"3ce9",x"37ba",x"bbfc",x"0000",x"2bdf",x"340b",x"3554",x"3a43",x"2661",x"37e4",x"bbd4",x"8000",x"328e",x"33e7",x"2438"),
(x"3a41",x"2065",x"3775",x"bbe7",x"0000",x"b0fd",x"3423",x"2104",x"3a41",x"3ce9",x"3775",x"bbfd",x"068d",x"aac8",x"3423",x"3554",x"3a41",x"24c7",x"37ba",x"bbff",x"0000",x"26a1",x"340b",x"22bc"),
(x"3a45",x"1d1b",x"3764",x"ba17",x"0000",x"b92f",x"343b",x"1d79",x"3a45",x"3ce9",x"3764",x"baa9",x"0000",x"b86d",x"343b",x"3554",x"3a41",x"2065",x"3775",x"bbe7",x"0000",x"b0fd",x"3423",x"2104"),
(x"3a4e",x"1a6a",x"3752",x"b98d",x"8000",x"b9c2",x"3453",x"1b5d",x"3a4e",x"3ce9",x"3752",x"b98d",x"8000",x"b9c2",x"3453",x"3554",x"3a45",x"1d1b",x"3764",x"ba17",x"0000",x"b92f",x"343b",x"1d79"),
(x"3aae",x"3ce9",x"376e",x"3bb7",x"8000",x"b434",x"3277",x"3554",x"3aa3",x"3ce9",x"3752",x"3a65",x"8000",x"b8cd",x"3248",x"3554",x"3aae",x"1ef5",x"376e",x"3b33",x"0000",x"b6f8",x"3276",x"21dd"),
(x"3a90",x"2869",x"3813",x"9e3f",x"bacb",x"3838",x"35c8",x"3482",x"3a4b",x"27a4",x"3802",x"a352",x"bab1",x"3860",x"35fb",x"3474",x"3a76",x"28ad",x"3818",x"a495",x"ba9b",x"3881",x"35db",x"3487"),
(x"3a4e",x"1a6a",x"3752",x"9c32",x"bb56",x"3661",x"35f6",x"3427",x"3a45",x"1d1b",x"3764",x"0a8d",x"baca",x"383a",x"35fd",x"342e",x"3aa3",x"1a08",x"3752",x"1a24",x"bb18",x"3761",x"35b6",x"3427"),
(x"3ab0",x"22af",x"3794",x"9953",x"bac8",x"383d",x"35ae",x"3444",x"3aae",x"1ef5",x"376e",x"9c81",x"baa0",x"387b",x"35af",x"3433",x"3a41",x"2065",x"3775",x"9da1",x"bab0",x"3862",x"3600",x"3436"),
(x"3aad",x"2680",x"37e5",x"1af6",x"bad3",x"382b",x"35b1",x"3467",x"3ab0",x"22af",x"3794",x"9953",x"bac8",x"383d",x"35ae",x"3444",x"3a41",x"24c7",x"37ba",x"128d",x"bad3",x"382c",x"3601",x"3454"),
(x"3aa1",x"2805",x"3807",x"1e73",x"baea",x"3806",x"35bb",x"3479",x"3aad",x"2680",x"37e5",x"1af6",x"bad3",x"382b",x"35b1",x"3467",x"3a43",x"2661",x"37e4",x"1b5f",x"badf",x"3817",x"3600",x"3466"),
(x"3aa1",x"2805",x"3807",x"1e73",x"baea",x"3806",x"35bb",x"3479",x"3a43",x"2661",x"37e4",x"1b5f",x"badf",x"3817",x"3600",x"3466",x"3a90",x"2869",x"3813",x"9e3f",x"bacb",x"3838",x"35c8",x"3482"),
(x"3ac4",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"3639",x"3346",x"3ad1",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"3620",x"334e",x"3adb",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"361f",x"3321"),
(x"3abe",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"363a",x"3356",x"3ac9",x"3ff0",x"3752",x"38fd",x"390a",x"3765",x"3622",x"3363",x"3ad1",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"3620",x"334e"),
(x"3abe",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"363a",x"3356",x"3ab3",x"3fec",x"378f",x"a8a8",x"3b7d",x"3597",x"363e",x"3365",x"3ac1",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"3624",x"336f"),
(x"3ac5",x"3fa8",x"3752",x"3afd",x"b17a",x"3748",x"3634",x"328d",x"3abc",x"3fa7",x"3777",x"3b1d",x"b0f4",x"36e3",x"3643",x"3291",x"3acb",x"3fd8",x"3786",x"3af1",x"b04f",x"37a7",x"3637",x"331f"),
(x"3abd",x"3f8b",x"3752",x"3b0e",x"aeb1",x"3757",x"363e",x"323c",x"3ab5",x"3f8a",x"376d",x"3af9",x"af50",x"37a0",x"3649",x"323c",x"3abc",x"3fa7",x"3777",x"3b1d",x"b0f4",x"36e3",x"3643",x"3291"),
(x"3ac1",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"3624",x"336f",x"3ab3",x"3fec",x"378f",x"a8a8",x"3b7d",x"3597",x"363e",x"3365",x"3aa9",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"3644",x"3373"),
(x"3aa9",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"3644",x"3373",x"3aa0",x"3fe2",x"378c",x"b9d1",x"382c",x"3723",x"364c",x"3387",x"3aa2",x"3fe5",x"3782",x"b9d9",x"3972",x"a970",x"3645",x"3385"),
(x"3abc",x"3fa7",x"3777",x"ab80",x"ac13",x"3bf8",x"35a9",x"31f0",x"3ab5",x"3f8a",x"376d",x"2faf",x"abf2",x"3bed",x"35ad",x"319a",x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3ac4",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"35a5",x"327f",x"3acb",x"3fd8",x"3786",x"282c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3ac4",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"35a6",x"32a5",x"3acb",x"3fd8",x"3786",x"282c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3abe",x"3fea",x"378e",x"2da8",x"257a",x"3bf7",x"35ab",x"32b3",x"3ac4",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"35a6",x"32a5"),
(x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ab2",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"3ab3",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"35b3",x"32b8"),
(x"3ab2",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3aa9",x"3fea",x"378e",x"ae38",x"2687",x"3bf5",x"35bc",x"32b1"),
(x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3aa0",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"35c2",x"329a"),
(x"3a9b",x"3fe0",x"378b",x"aefe",x"af3d",x"3be6",x"35c6",x"3293",x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274"),
(x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3a9b",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"35c4",x"323e",x"3a9b",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"3aa4",x"3faa",x"3777",x"2c2f",x"accc",x"3bf5",x"35bc",x"31f5",x"3a9b",x"3fa8",x"3777",x"2bc1",x"ab62",x"3bf8",x"35c2",x"31f0",x"3a9b",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"35c4",x"323e"),
(x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3a9a",x"3f83",x"3770",x"2e76",x"a7e2",x"3bf4",x"35c1",x"3184",x"3a9b",x"3fa8",x"3777",x"2bc1",x"ab62",x"3bf8",x"35c2",x"31f0"),
(x"3aa4",x"3faa",x"3777",x"2c2f",x"accc",x"3bf5",x"35bc",x"31f5",x"3aa8",x"3fab",x"3775",x"3235",x"abce",x"3bd5",x"35b8",x"31f9",x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c"),
(x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245",x"3aa8",x"3fab",x"3775",x"3235",x"abce",x"3bd5",x"35b8",x"31f9"),
(x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3aa7",x"3fd5",x"3782",x"2e90",x"aed5",x"3be9",x"35bb",x"3274",x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245"),
(x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293"),
(x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3aaf",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"35b6",x"32a0"),
(x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3ab2",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"3ab4",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1",x"3ab4",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"3ac4",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"35a5",x"327f",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298"),
(x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3aa8",x"3fab",x"3775",x"3235",x"abce",x"3bd5",x"35b8",x"31f9",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"3aa7",x"3fd5",x"3782",x"2e90",x"aed5",x"3be9",x"35bb",x"3274",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298"),
(x"3aaf",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"35b6",x"32a0",x"3ab4",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"35b3",x"32a3",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"3a9a",x"3f83",x"3770",x"3be8",x"9d04",x"30d3",x"35e4",x"32f1",x"3a98",x"3fa7",x"378a",x"3bec",x"2581",x"3053",x"35e3",x"3284",x"3a9a",x"3fa8",x"3783",x"3b1f",x"a907",x"3740",x"35e6",x"3285"),
(x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236",x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236",x"3a9a",x"3fa8",x"3783",x"3b1f",x"a907",x"3740",x"35e6",x"3285"),
(x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203",x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236"),
(x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203"),
(x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5"),
(x"3a93",x"3fe1",x"37b6",x"3a64",x"b8cb",x"29c5",x"35e0",x"31dc",x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"3a93",x"3fe1",x"37b6",x"3a64",x"b8cb",x"29c5",x"35e0",x"31dc",x"3a93",x"3fe1",x"37c1",x"3add",x"b464",x"b6f2",x"35dc",x"31dd",x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"3a93",x"3fe1",x"37c1",x"3add",x"b464",x"b6f2",x"35dc",x"31dd",x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a99",x"3fc5",x"37c6",x"3af7",x"2fc0",x"b79e",x"35d2",x"322a"),
(x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a97",x"3fa9",x"379f",x"3bfa",x"2c34",x"a7c1",x"35dc",x"327e",x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"3a97",x"3fa9",x"379f",x"3bfa",x"2c34",x"a7c1",x"35dc",x"327e",x"3a99",x"3f8a",x"3790",x"3bff",x"25e3",x"1e73",x"35da",x"32db",x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"3a99",x"3f8a",x"3790",x"3bff",x"25e3",x"1e73",x"35da",x"32db",x"3a99",x"3f88",x"3798",x"3be2",x"a70a",x"315a",x"35d6",x"32dd",x"3a98",x"3fa8",x"37b2",x"3be6",x"a82f",x"30eb",x"35d4",x"327f"),
(x"3a99",x"3fc3",x"37d1",x"3bf3",x"a804",x"2ec5",x"35cd",x"322c",x"3a99",x"3fc5",x"37c6",x"3af7",x"2fc0",x"b79e",x"35d2",x"322a",x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"3a99",x"3fc3",x"37d1",x"3bf3",x"a804",x"2ec5",x"35cd",x"322c",x"3a98",x"3fd3",x"37de",x"3be7",x"9cea",x"30f2",x"35cc",x"31fd",x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"3a98",x"3fd3",x"37de",x"3be7",x"9cea",x"30f2",x"35cc",x"31fd",x"3a98",x"3fdf",x"37dc",x"3bdc",x"28a8",x"31da",x"35d0",x"31db",x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"3a98",x"3fdf",x"37dc",x"3bdc",x"28a8",x"31da",x"35d0",x"31db",x"3a99",x"3fe6",x"37cc",x"3bf2",x"2959",x"2ec5",x"35d9",x"31c8",x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"3a99",x"3fe6",x"37cc",x"3bf2",x"2959",x"2ec5",x"35d9",x"31c8",x"3a9a",x"3fe8",x"37b8",x"3bfd",x"2587",x"2a48",x"35e1",x"31c5",x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"3a9a",x"3fe7",x"37a7",x"3bff",x"1ec2",x"2532",x"35e8",x"31ca",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3",x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"3a9a",x"3fe0",x"378e",x"3bf9",x"1818",x"2d46",x"35f0",x"31e1",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"3a9a",x"3fe0",x"378e",x"3bf9",x"1818",x"2d46",x"35f0",x"31e1",x"3a9b",x"3fe0",x"378b",x"3aff",x"ad07",x"37a5",x"35f2",x"31e1",x"3a9b",x"3fd4",x"3784",x"3beb",x"a025",x"3083",x"35f2",x"3204"),
(x"3a9b",x"3fd4",x"3784",x"3beb",x"a025",x"3083",x"35f2",x"3204",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5"),
(x"3a9b",x"3fc3",x"377f",x"3bd2",x"a2f6",x"32b9",x"35f0",x"3237",x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203"),
(x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236",x"3a9b",x"3fc3",x"377f",x"3bd2",x"a2f6",x"32b9",x"35f0",x"3237",x"3a9b",x"3fa8",x"3777",x"3bc7",x"a659",x"336e",x"35eb",x"3285"),
(x"3a9a",x"3fa8",x"3783",x"3b1f",x"a907",x"3740",x"35e6",x"3285",x"3a9b",x"3fa8",x"3777",x"3bc7",x"a659",x"336e",x"35eb",x"3285",x"3a9a",x"3f83",x"3770",x"3be8",x"9d04",x"30d3",x"35e4",x"32f1"),
(x"3a98",x"3fa7",x"378a",x"3bec",x"2581",x"3053",x"35e3",x"3284",x"3a9a",x"3f83",x"3770",x"3be8",x"9d04",x"30d3",x"35e4",x"32f1",x"3a99",x"3f8a",x"3790",x"3bff",x"25e3",x"1e73",x"35da",x"32db"),
(x"3a97",x"3fa9",x"379f",x"3bfa",x"2c34",x"a7c1",x"35dc",x"327e",x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236"),
(x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205"),
(x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec"),
(x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a93",x"3fe1",x"37c1",x"3add",x"b464",x"b6f2",x"35dc",x"31dd",x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"3a93",x"3fe1",x"37c1",x"3add",x"b464",x"b6f2",x"35dc",x"31dd",x"3a93",x"3fe1",x"37b6",x"3a64",x"b8cb",x"29c5",x"35e0",x"31dc",x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"3a98",x"3fa8",x"37b2",x"3870",x"b1f2",x"3a7c",x"35f5",x"3500",x"3a99",x"3f88",x"3798",x"386c",x"b134",x"3a89",x"35f5",x"3530",x"3a7a",x"3f87",x"37c0",x"a48e",x"b255",x"3bd7",x"35d8",x"352f"),
(x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a99",x"3fc3",x"37d1",x"3885",x"b324",x"3a5a",x"35f4",x"34d4"),
(x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a98",x"3fd3",x"37de",x"389a",x"ad78",x"3a82",x"35f2",x"34bc"),
(x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a98",x"3fdf",x"37dc",x"3869",x"323c",x"3a7d",x"35f0",x"34aa"),
(x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a79",x"3feb",x"37e2",x"9953",x"3ada",x"3821",x"35d7",x"349e",x"3a99",x"3fe6",x"37cc",x"3783",x"398b",x"385f",x"35ef",x"349c"),
(x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495",x"3a9a",x"3fe8",x"37b8",x"35d5",x"3b70",x"2a94",x"35f1",x"3494",x"3a99",x"3fe6",x"37cc",x"3783",x"398b",x"385f",x"35ef",x"349c"),
(x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e",x"3a9a",x"3fe7",x"37a7",x"3572",x"3a96",x"b740",x"35f3",x"348e",x"3a9a",x"3fe8",x"37b8",x"35d5",x"3b70",x"2a94",x"35f1",x"3494"),
(x"3a91",x"3fe7",x"379c",x"3620",x"3a0a",x"b841",x"35ed",x"3488",x"3a9a",x"3fe0",x"378e",x"381d",x"395a",x"b849",x"35f9",x"3481",x"3a9a",x"3fe7",x"37a7",x"3572",x"3a96",x"b740",x"35f3",x"348e"),
(x"3a91",x"3fe7",x"379c",x"3620",x"3a0a",x"b841",x"35ed",x"3488",x"3a97",x"3fe1",x"378b",x"3994",x"399e",x"b083",x"35f6",x"3480",x"3a9a",x"3fe0",x"378e",x"381d",x"395a",x"b849",x"35f9",x"3481"),
(x"3aa0",x"3fe2",x"378c",x"b9d1",x"382c",x"3723",x"364c",x"3387",x"3a9b",x"3fe0",x"378b",x"b88b",x"36b7",x"39a9",x"364e",x"338f",x"3a9a",x"3fe1",x"3786",x"b88d",x"3867",x"38e2",x"364c",x"3391"),
(x"3a9a",x"3fe1",x"3786",x"381b",x"39f5",x"36cf",x"35f8",x"347e",x"3a9b",x"3fe0",x"378b",x"38bf",x"3999",x"3659",x"35fa",x"3480",x"3a9a",x"3fe0",x"378e",x"381d",x"395a",x"b849",x"35f9",x"3481"),
(x"3a18",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"35ab",x"2e93",x"3a22",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"35ab",x"2e39",x"3a2f",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"35c4",x"2e47"),
(x"3a22",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"35ab",x"2e39",x"3a2a",x"3ff0",x"3752",x"b8fd",x"390a",x"3765",x"35ad",x"2e10",x"3a35",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"35c6",x"2e27"),
(x"3a35",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"35c6",x"2e27",x"3a2a",x"3ff0",x"3752",x"b8fd",x"390a",x"3765",x"35ad",x"2e10",x"3a33",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"35af",x"2df7"),
(x"3a28",x"3fd8",x"3786",x"bad9",x"b071",x"37f4",x"35c2",x"2e97",x"3a38",x"3fa6",x"3775",x"bacd",x"b078",x"380f",x"35cf",x"2fb9",x"3a2e",x"3fa8",x"3752",x"badc",x"b152",x"37c7",x"35c0",x"2fbb"),
(x"3a38",x"3fa6",x"3775",x"bacd",x"b078",x"380f",x"35cf",x"2fb9",x"3a3f",x"3f88",x"376d",x"ba64",x"ad63",x"38c3",x"35d7",x"3033",x"3a34",x"3f8b",x"3752",x"bab6",x"ad4f",x"384d",x"35c9",x"302f"),
(x"3a40",x"3fec",x"378f",x"28ac",x"3b7d",x"3597",x"35ca",x"2e09",x"3a33",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"35af",x"2df7",x"3a4b",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"3a52",x"3fe5",x"3782",x"39dc",x"3971",x"a62b",x"35d1",x"2dca",x"3a54",x"3fe2",x"378c",x"39bb",x"383c",x"3743",x"35d7",x"2dc5",x"3a4b",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e",x"3a3f",x"3f88",x"376d",x"b03d",x"a8e0",x"3bec",x"3614",x"3130",x"3a38",x"3fa6",x"3775",x"ab9a",x"acf0",x"3bf6",x"3611",x"30d8"),
(x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2",x"3a38",x"3fa6",x"3775",x"ab9a",x"acf0",x"3bf6",x"3611",x"30d8",x"3a28",x"3fd8",x"3786",x"ae54",x"ae94",x"3beb",x"3607",x"3046"),
(x"3a28",x"3fd8",x"3786",x"ae54",x"ae94",x"3beb",x"3607",x"3046",x"3a2f",x"3fe5",x"378d",x"ae28",x"ac9e",x"3bf1",x"360d",x"3020",x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026"),
(x"3a2f",x"3fe5",x"378d",x"ae28",x"ac9e",x"3bf1",x"360d",x"3020",x"3a35",x"3fea",x"378e",x"ada8",x"257a",x"3bf7",x"3612",x"3012",x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a",x"3a35",x"3fea",x"378e",x"ada8",x"257a",x"3bf7",x"3612",x"3012",x"3a40",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"361b",x"300d"),
(x"3a41",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"361b",x"3016",x"3a40",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"361b",x"300d",x"3a4b",x"3fea",x"378e",x"2e38",x"2687",x"3bf5",x"3623",x"3014"),
(x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a4b",x"3fea",x"378e",x"2e38",x"2687",x"3bf5",x"3623",x"3014",x"3a54",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"3a58",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"362d",x"3032",x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051",x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f"),
(x"3a59",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"362d",x"3054",x"3a58",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"362b",x"3087",x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082"),
(x"3a58",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"362b",x"3087",x"3a58",x"3fa8",x"3777",x"a6fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"3a50",x"3faa",x"3777",x"ac34",x"acb0",x"3bf5",x"3623",x"30d0"),
(x"3a58",x"3fa8",x"3777",x"a6fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"3a5a",x"3f89",x"3770",x"a987",x"a828",x"3bfc",x"3628",x"312f",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"3a4b",x"3fab",x"3775",x"b227",x"ab9d",x"3bd6",x"361f",x"30cb",x"3a50",x"3faa",x"3777",x"ac34",x"acb0",x"3bf5",x"3623",x"30d0",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"3a4b",x"3fab",x"3775",x"b227",x"ab9d",x"3bd6",x"361f",x"30cb",x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080",x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082"),
(x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080",x"3a4c",x"3fd5",x"3782",x"ae90",x"aed5",x"3be9",x"3623",x"3050",x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051"),
(x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051",x"3a4c",x"3fd5",x"3782",x"ae90",x"aed5",x"3be9",x"3623",x"3050",x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f",x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032",x"3a44",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"361d",x"3025"),
(x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a44",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"361d",x"3025",x"3a40",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"361a",x"3022"),
(x"3a40",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"361a",x"3022",x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026"),
(x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a2f",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"360d",x"3046"),
(x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2"),
(x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e",x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2",x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0"),
(x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"3a4b",x"3fab",x"3775",x"b227",x"ab9d",x"3bd6",x"361f",x"30cb",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080"),
(x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a4c",x"3fd5",x"3782",x"ae90",x"aed5",x"3be9",x"3623",x"3050"),
(x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a40",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"361a",x"3022",x"3a44",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"361d",x"3025"),
(x"3a5c",x"3fa8",x"378a",x"bbe0",x"2467",x"319c",x"360d",x"31c3",x"3a5a",x"3f89",x"3770",x"bbf0",x"1d6d",x"2fcb",x"360f",x"3168",x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4"),
(x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4",x"3a5a",x"3fc2",x"378b",x"ba70",x"a9d2",x"38bb",x"3615",x"3211",x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"3a5a",x"3fc2",x"378b",x"ba70",x"a9d2",x"38bb",x"3615",x"3211",x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263",x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b"),
(x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263",x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268"),
(x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b",x"3a5f",x"3fe2",x"37b7",x"ba93",x"b88d",x"2474",x"360a",x"326f"),
(x"3a5f",x"3fe2",x"37b7",x"ba93",x"b88d",x"2474",x"360a",x"326f",x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277"),
(x"3a5f",x"3fe1",x"37c3",x"bb15",x"b383",x"b669",x"3606",x"326c",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266",x"3a5b",x"3fd3",x"37d2",x"ba75",x"2987",x"b8b5",x"35fc",x"3249"),
(x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a5b",x"3fd3",x"37d2",x"ba75",x"2987",x"b8b5",x"35fc",x"3249",x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e"),
(x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e",x"3a5b",x"3fa9",x"37a5",x"bbef",x"2703",x"afed",x"3603",x"31c9",x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9"),
(x"3a5a",x"3f85",x"378d",x"bbff",x"2504",x"1d87",x"3604",x"3160",x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9",x"3a5b",x"3fa9",x"37a5",x"bbef",x"2703",x"afed",x"3603",x"31c9"),
(x"3a5b",x"3fa8",x"37b0",x"bbfa",x"a20a",x"2ca3",x"35ff",x"31c8",x"3a5b",x"3f84",x"3797",x"bbe3",x"a752",x"313e",x"3600",x"315e",x"3a5a",x"3f85",x"378d",x"bbff",x"2504",x"1d87",x"3604",x"3160"),
(x"3a5b",x"3fa9",x"37a5",x"bbef",x"2703",x"afed",x"3603",x"31c9",x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e",x"3a5b",x"3fc3",x"37d0",x"bbff",x"a2f6",x"24f0",x"35f8",x"321b"),
(x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e",x"3a5b",x"3fd3",x"37d2",x"ba75",x"2987",x"b8b5",x"35fc",x"3249",x"3a5a",x"3fd3",x"37dc",x"bbff",x"15bc",x"a66c",x"35f8",x"324b"),
(x"3a5a",x"3fd3",x"37dc",x"bbff",x"15bc",x"a66c",x"35f8",x"324b",x"3a5b",x"3fd3",x"37d2",x"ba75",x"2987",x"b8b5",x"35fc",x"3249",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"3a5a",x"3fde",x"37db",x"bbff",x"1953",x"2560",x"35fb",x"326b",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277"),
(x"3a5a",x"3fe6",x"37cd",x"bbf7",x"29c5",x"2d1b",x"3603",x"327f",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277",x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b"),
(x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b",x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a5a",x"3fe7",x"37a7",x"bbff",x"0a8d",x"2694",x"3612",x"327d"),
(x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263",x"3a59",x"3fe0",x"378e",x"bbf8",x"1553",x"2d82",x"361b",x"3266"),
(x"3a58",x"3fe0",x"378b",x"baff",x"ad09",x"37a5",x"361c",x"3266",x"3a59",x"3fe0",x"378e",x"bbf8",x"1553",x"2d82",x"361b",x"3266",x"3a59",x"3fd4",x"3784",x"bbea",x"a025",x"3095",x"361c",x"3243"),
(x"3a59",x"3fd4",x"3784",x"bbea",x"a025",x"3095",x"361c",x"3243",x"3a59",x"3fe0",x"378e",x"bbf8",x"1553",x"2d82",x"361b",x"3266",x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263"),
(x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a5a",x"3fc2",x"378b",x"ba70",x"a9d2",x"38bb",x"3615",x"3211",x"3a58",x"3fc3",x"377f",x"bbce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4",x"3a58",x"3fa8",x"3777",x"bbc5",x"a793",x"3388",x"3615",x"31c2",x"3a58",x"3fc3",x"377f",x"bbce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"3a58",x"3fa8",x"3777",x"bbc5",x"a793",x"3388",x"3615",x"31c2",x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4",x"3a5a",x"3f89",x"3770",x"bbf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9",x"3a5a",x"3f85",x"378d",x"bbff",x"2504",x"1d87",x"3604",x"3160",x"3a5a",x"3f89",x"3770",x"bbf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9",x"3a5c",x"3fa8",x"378a",x"bbe0",x"2467",x"319c",x"360d",x"31c3",x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"3a60",x"3fc5",x"37be",x"bbeb",x"2c4d",x"b006",x"3601",x"321f",x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211",x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242",x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b"),
(x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b",x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268"),
(x"3a5f",x"3fe2",x"37b7",x"ba93",x"b88d",x"2474",x"360a",x"326f",x"3a5f",x"3fe1",x"37c3",x"bb15",x"b383",x"b669",x"3606",x"326c",x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268"),
(x"3a7a",x"3f87",x"37c0",x"a48e",x"b255",x"3bd7",x"35d8",x"352f",x"3a5b",x"3f84",x"3797",x"b82d",x"b0b5",x"3ab8",x"35bc",x"3537",x"3a5b",x"3fa8",x"37b0",x"b87f",x"b1e6",x"3a73",x"35ba",x"3500"),
(x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a5b",x"3fa8",x"37b0",x"b87f",x"b1e6",x"3a73",x"35ba",x"3500",x"3a5b",x"3fc3",x"37d0",x"b896",x"b2c0",x"3a54",x"35bb",x"34d5"),
(x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a5b",x"3fc3",x"37d0",x"b896",x"b2c0",x"3a54",x"35bb",x"34d5",x"3a5a",x"3fd3",x"37dc",x"b892",x"ade1",x"3a86",x"35bc",x"34bc"),
(x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a5a",x"3fd3",x"37dc",x"b892",x"ade1",x"3a86",x"35bc",x"34bc",x"3a5a",x"3fde",x"37db",x"b885",x"3126",x"3a79",x"35be",x"34ab"),
(x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a5a",x"3fde",x"37db",x"b885",x"3126",x"3a79",x"35be",x"34ab",x"3a5a",x"3fe6",x"37cd",x"b7e6",x"396d",x"385a",x"35bf",x"349d"),
(x"3a5a",x"3fe6",x"37cd",x"b7e6",x"396d",x"385a",x"35bf",x"349d",x"3a5a",x"3fe8",x"37b8",x"b61b",x"3b60",x"2bbe",x"35be",x"3495",x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495"),
(x"3a5a",x"3fe8",x"37b8",x"b61b",x"3b60",x"2bbe",x"35be",x"3495",x"3a5a",x"3fe7",x"37a7",x"b619",x"3a76",x"b730",x"35bb",x"348f",x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e"),
(x"3a5a",x"3fe7",x"37a7",x"b619",x"3a76",x"b730",x"35bb",x"348f",x"3a59",x"3fe0",x"378e",x"b967",x"383c",x"b81a",x"35b4",x"3483",x"3a61",x"3fe4",x"3789",x"b646",x"3a25",x"b80b",x"35bd",x"3481"),
(x"3a5d",x"3fe1",x"378b",x"b8bd",x"3a6d",x"2c06",x"35b7",x"3482",x"3a61",x"3fe4",x"3789",x"b646",x"3a25",x"b80b",x"35bd",x"3481",x"3a59",x"3fe0",x"378e",x"b967",x"383c",x"b81a",x"35b4",x"3483"),
(x"3a5b",x"3fe1",x"3782",x"38d3",x"3873",x"3892",x"35d6",x"2daa",x"3a58",x"3fe0",x"378b",x"38ee",x"37c0",x"38f6",x"35d9",x"2db4",x"3a54",x"3fe2",x"378c",x"39bb",x"383c",x"3743",x"35d7",x"2dc5"),
(x"3a5d",x"3fe1",x"378b",x"b8bd",x"3a6d",x"2c06",x"35b7",x"3482",x"3a59",x"3fe0",x"378e",x"b967",x"383c",x"b81a",x"35b4",x"3483",x"3a58",x"3fe0",x"378b",x"b862",x"3a94",x"30e6",x"35b3",x"3481"),
(x"3a34",x"3f8b",x"3752",x"bab6",x"ad4f",x"384d",x"35c9",x"302f",x"3a3f",x"3f88",x"376d",x"ba64",x"ad63",x"38c3",x"35d7",x"3033",x"3a3e",x"3f7e",x"376e",x"babb",x"aad9",x"384d",x"35d9",x"3052"),
(x"3a3f",x"3f88",x"376d",x"b03d",x"a8e0",x"3bec",x"3614",x"3130",x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e",x"3a48",x"3f83",x"3770",x"ae2b",x"280b",x"3bf5",x"361a",x"3141"),
(x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e",x"3a48",x"3f83",x"3770",x"ae2b",x"280b",x"3bf5",x"361a",x"3141",x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e"),
(x"3a48",x"3f83",x"3770",x"ae2b",x"280b",x"3bf5",x"361a",x"3141",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e",x"3a5a",x"3f89",x"3770",x"a987",x"a828",x"3bfc",x"3628",x"312f"),
(x"3ab3",x"3f7a",x"376e",x"3b00",x"aaa4",x"37b3",x"364e",x"320e",x"3ab5",x"3f8a",x"376d",x"3af9",x"af50",x"37a0",x"3649",x"323c",x"3abd",x"3f8b",x"3752",x"3b0e",x"aeb1",x"3757",x"363e",x"323c"),
(x"3ab5",x"3f8a",x"376d",x"2faf",x"abf2",x"3bed",x"35ad",x"319a",x"3ab3",x"3f7a",x"376e",x"2d23",x"068d",x"3bf9",x"35ad",x"316b",x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"3ab3",x"3f7a",x"376e",x"2d23",x"068d",x"3bf9",x"35ad",x"316b",x"3aa2",x"3f7f",x"3770",x"2938",x"1b93",x"3bfe",x"35ba",x"3179"),
(x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3aa2",x"3f7f",x"3770",x"2938",x"1b93",x"3bfe",x"35ba",x"3179",x"3a9a",x"3f83",x"3770",x"2e76",x"a7e2",x"3bf4",x"35c1",x"3184"),
(x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9",x"3ac6",x"4032",x"377d",x"3601",x"3ae5",x"3571",x"3629",x"2fc2",x"3ac7",x"4030",x"3794",x"3663",x"3a38",x"37c6",x"3623",x"2fe3"),
(x"3ad0",x"4030",x"377a",x"3864",x"3a40",x"34bc",x"3630",x"2fdb",x"3ac6",x"4032",x"377d",x"3601",x"3ae5",x"3571",x"3629",x"2fc2",x"3acc",x"4033",x"3752",x"324d",x"3bb2",x"31fb",x"3638",x"2fa0"),
(x"3ad0",x"4030",x"377a",x"3068",x"a815",x"3beb",x"362f",x"3205",x"3ac4",x"402c",x"377c",x"3068",x"a815",x"3beb",x"362f",x"3221",x"3ac6",x"4032",x"377d",x"3068",x"a815",x"3beb",x"3626",x"3206"),
(x"3ac7",x"4030",x"3794",x"3be8",x"aaec",x"b08c",x"35d7",x"1fd1",x"3ac6",x"4032",x"377d",x"3be8",x"aaec",x"b08c",x"35e0",x"1e8d",x"3ac4",x"402c",x"377c",x"3be8",x"aaec",x"b08c",x"35e0",x"214e"),
(x"3ad0",x"4030",x"377a",x"3a71",x"b86a",x"32e4",x"3645",x"3436",x"3ad7",x"4031",x"3752",x"3a9b",x"b7a9",x"34c2",x"3635",x"3436",x"3ac4",x"402c",x"377c",x"39ed",x"b7fd",x"372e",x"364a",x"3429"),
(x"3a98",x"4021",x"3787",x"388f",x"b80c",x"392d",x"3662",x"3401",x"3ab4",x"4030",x"37b3",x"389d",x"b810",x"391d",x"3662",x"3434",x"3abc",x"4027",x"376e",x"38ec",x"b7ef",x"38e6",x"364a",x"3418"),
(x"3ab4",x"4030",x"37b3",x"b422",x"b30f",x"3b86",x"359c",x"33ee",x"3a98",x"4021",x"3787",x"b776",x"b053",x"3afe",x"359c",x"3429",x"3aab",x"4030",x"37ae",x"b777",x"b053",x"3afe",x"3595",x"33f3"),
(x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9",x"3ab4",x"4030",x"37b3",x"348b",x"3a03",x"38c2",x"3611",x"2fda",x"3aab",x"4030",x"37ae",x"b35d",x"39d9",x"3923",x"360d",x"2fc2"),
(x"3aab",x"4030",x"37ae",x"b777",x"b053",x"3afe",x"3595",x"33f3",x"3a98",x"4021",x"3787",x"b776",x"b053",x"3afe",x"359c",x"3429",x"3aa2",x"4031",x"379f",x"b8fe",x"ab38",x"3a3c",x"358d",x"33fa"),
(x"3aa2",x"4031",x"379f",x"b54f",x"39c9",x"38d8",x"360b",x"2fa1",x"3a94",x"4033",x"3780",x"acce",x"3bc5",x"3335",x"360d",x"2f61",x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"3aae",x"4033",x"3752",x"1d38",x"3bf5",x"2e94",x"3627",x"2f61",x"3acc",x"4033",x"3752",x"324d",x"3bb2",x"31fb",x"3638",x"2fa0",x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9",x"3acc",x"4033",x"3752",x"324d",x"3bb2",x"31fb",x"3638",x"2fa0",x"3ac6",x"4032",x"377d",x"3601",x"3ae5",x"3571",x"3629",x"2fc2"),
(x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349",x"3a81",x"4031",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"3355",x"3a78",x"4030",x"37da",x"b146",x"3a67",x"389c",x"3659",x"3362"),
(x"3a81",x"4031",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"3355",x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3a9b",x"4030",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"335c"),
(x"3a8a",x"4030",x"37da",x"b950",x"a0dd",x"39fa",x"35e9",x"2ccc",x"3a81",x"402d",x"37cb",x"b950",x"a0dd",x"39fa",x"35e9",x"2d02",x"3a81",x"4031",x"37cb",x"b950",x"a0dd",x"39fa",x"35df",x"2cd5"),
(x"3a78",x"4030",x"37da",x"393c",x"95bc",x"3a0c",x"35ec",x"2c9f",x"3a81",x"4031",x"37cb",x"393c",x"95bc",x"3a0c",x"35ec",x"2cc6",x"3a81",x"402d",x"37cb",x"393c",x"95bc",x"3a0c",x"35df",x"2cab"),
(x"3a8a",x"4030",x"37da",x"3325",x"b878",x"3a63",x"367b",x"30d7",x"3a9b",x"4030",x"37d1",x"333b",x"b811",x"3aa5",x"3689",x"30d9",x"3a81",x"402d",x"37cb",x"9e0a",x"b823",x"3ad8",x"3676",x"30ef"),
(x"3a64",x"4023",x"3791",x"b252",x"b816",x"3ab1",x"3661",x"3135",x"3a62",x"4030",x"37cd",x"b1e7",x"b81a",x"3ab5",x"365e",x"30e1",x"3a82",x"4026",x"37ad",x"23bb",x"b81b",x"3add",x"3677",x"311b"),
(x"3a62",x"4030",x"37cd",x"baf6",x"b475",x"367c",x"35a4",x"3094",x"3a64",x"4023",x"3791",x"bad4",x"b414",x"3743",x"35b5",x"3046",x"3a5e",x"4030",x"37ba",x"bb3a",x"b41e",x"357a",x"35ac",x"3093"),
(x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349",x"3a62",x"4030",x"37cd",x"b58a",x"3a1b",x"385c",x"3649",x"3358",x"3a5e",x"4030",x"37ba",x"b926",x"39b7",x"3463",x"3645",x"334a"),
(x"3a5e",x"4030",x"37ba",x"bb3a",x"b41e",x"357a",x"35ac",x"3093",x"3a64",x"4023",x"3791",x"bad4",x"b414",x"3743",x"35b5",x"3046",x"3a59",x"4030",x"379b",x"babf",x"b3b7",x"37af",x"35b9",x"3091"),
(x"3a59",x"4030",x"379b",x"b825",x"3acf",x"2d30",x"3640",x"3332",x"3a66",x"4032",x"3781",x"b1af",x"3bdf",x"1c18",x"364b",x"331d",x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"3a94",x"4033",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"331d",x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349",x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3a81",x"4031",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"3355"),
(x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3a94",x"4033",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"331d",x"3aa2",x"4031",x"379f",x"394b",x"39eb",x"af9d",x"367a",x"3337"),
(x"3a9b",x"4030",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"335c",x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3aa3",x"4030",x"37ba",x"392f",x"39d8",x"32de",x"367a",x"334c"),
(x"3a9b",x"4030",x"37d1",x"39f1",x"b5fe",x"3870",x"3649",x"2eb4",x"3aa3",x"4030",x"37ba",x"3b76",x"b463",x"3373",x"3640",x"2ea4",x"3a98",x"4021",x"3787",x"3b76",x"b463",x"3373",x"3649",x"2de4"),
(x"3aa2",x"4031",x"379f",x"3bda",x"afe2",x"b0aa",x"3637",x"2e90",x"3a98",x"4021",x"3787",x"3b76",x"b463",x"3373",x"3649",x"2de4",x"3aa3",x"4030",x"37ba",x"3b76",x"b463",x"3373",x"3640",x"2ea4"),
(x"3a60",x"4023",x"378f",x"b2ea",x"b07f",x"3bba",x"35b9",x"3044",x"3a59",x"4030",x"379b",x"babf",x"b3b7",x"37ae",x"35b9",x"3091",x"3a64",x"4023",x"3791",x"bad4",x"b414",x"3743",x"35b5",x"3046"),
(x"3a59",x"4030",x"379b",x"365b",x"ac2a",x"3b52",x"366b",x"3506",x"3a60",x"4023",x"378f",x"a822",x"af6e",x"3bf1",x"366b",x"352d",x"3a5e",x"4021",x"378e",x"b4a7",x"b630",x"3b00",x"3668",x"3531"),
(x"3a3b",x"4028",x"376e",x"b92f",x"b7c9",x"38af",x"3649",x"3520",x"3a44",x"4030",x"37b0",x"b5ad",x"b6ed",x"3aa0",x"3659",x"3502",x"3a5e",x"4021",x"378e",x"b4a7",x"b630",x"3b00",x"3668",x"3531"),
(x"3a44",x"4030",x"37b0",x"b5ad",x"b6ed",x"3aa0",x"3659",x"3502",x"3a32",x"402c",x"377a",x"b9d4",x"b83f",x"36e9",x"3645",x"3511",x"3a30",x"402f",x"378b",x"b815",x"b8b5",x"3904",x"3646",x"3507"),
(x"3a28",x"4030",x"3775",x"ba72",x"b85a",x"3373",x"363b",x"3507",x"3a32",x"402c",x"377a",x"b9d4",x"b83f",x"36e9",x"3645",x"3511",x"3a21",x"4031",x"3752",x"ba84",x"b81e",x"3444",x"362e",x"350b"),
(x"3a32",x"4032",x"3780",x"bbd2",x"3047",x"b134",x"35bb",x"2006",x"3a32",x"4030",x"3797",x"bb81",x"34c0",x"31b8",x"35bb",x"214e",x"3a30",x"402f",x"378b",x"bbd2",x"3047",x"b133",x"35b6",x"210c"),
(x"3a32",x"4032",x"3780",x"b66c",x"ad14",x"3b4c",x"362f",x"31e1",x"3a32",x"402c",x"377a",x"b612",x"af46",x"3b58",x"362f",x"3202",x"3a28",x"4030",x"3775",x"b66c",x"ad14",x"3b4c",x"3626",x"31ed"),
(x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f",x"3a44",x"4030",x"37b0",x"9fc8",x"3964",x"39e8",x"360f",x"2e1f",x"3a32",x"4030",x"3797",x"b553",x"3a2a",x"3858",x"361e",x"2e0a"),
(x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f",x"3a60",x"4033",x"3777",x"3179",x"3b46",x"3611",x"3613",x"2e9a",x"3a59",x"4030",x"379b",x"35ee",x"392f",x"3951",x"3609",x"2e60"),
(x"3a59",x"4030",x"379b",x"35ee",x"392f",x"3951",x"3609",x"2e60",x"3a60",x"4033",x"3777",x"3179",x"3b46",x"3611",x"3613",x"2e9a",x"3a66",x"4032",x"3781",x"3106",x"3a66",x"38a1",x"360c",x"2e9b"),
(x"3a55",x"4033",x"375d",x"a8bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"3a60",x"4033",x"3777",x"3179",x"3b46",x"3611",x"3613",x"2e9a",x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f"),
(x"3a2a",x"4033",x"3752",x"b410",x"3b92",x"3261",x"3637",x"2e3f",x"3a2a",x"4032",x"3777",x"b91e",x"39e6",x"32f0",x"362c",x"2e19",x"3a28",x"4030",x"3775",x"b9b9",x"391a",x"348e",x"362e",x"2e0a"),
(x"3a50",x"4033",x"3752",x"a4bc",x"3be9",x"30b5",x"3625",x"2e99",x"3a55",x"4033",x"375d",x"a8bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"3a32",x"4032",x"3780",x"ade3",x"3bd5",x"31ce",x"3625",x"2e26"),
(x"3a32",x"4032",x"3780",x"ade3",x"3bd5",x"31ce",x"3625",x"2e26",x"3a2a",x"4032",x"3777",x"b91e",x"39e6",x"32f0",x"362c",x"2e19",x"3a2a",x"4033",x"3752",x"b410",x"3b92",x"3261",x"3637",x"2e3f"),
(x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db",x"3ac6",x"405d",x"377d",x"3600",x"3ae5",x"3571",x"365f",x"33e0",x"3ac7",x"405b",x"3794",x"3663",x"3a38",x"37c6",x"3659",x"33f1"),
(x"3ad0",x"405b",x"377a",x"3865",x"3a40",x"34bc",x"3665",x"33ed",x"3ac6",x"405d",x"377d",x"3600",x"3ae5",x"3571",x"365f",x"33e0",x"3acc",x"405e",x"3752",x"324d",x"3bb2",x"31fb",x"366d",x"33ce"),
(x"3ad0",x"405b",x"377a",x"3068",x"a815",x"3beb",x"362f",x"3224",x"3ac4",x"4057",x"377c",x"3068",x"a815",x"3beb",x"362f",x"3241",x"3ac6",x"405d",x"377d",x"3068",x"a815",x"3beb",x"3626",x"3226"),
(x"3ac7",x"405b",x"3794",x"3be8",x"aaec",x"b08c",x"35eb",x"210c",x"3ac6",x"405d",x"377d",x"3be8",x"aaec",x"b08c",x"35e1",x"20e0",x"3ac4",x"4057",x"377c",x"3be8",x"aaec",x"b08c",x"35eb",x"1e8d"),
(x"3ad0",x"405b",x"377a",x"3a71",x"b86a",x"32e5",x"3655",x"3309",x"3ad7",x"405c",x"3752",x"3a92",x"b7f9",x"346d",x"3646",x"3307",x"3ac4",x"4057",x"377c",x"39d5",x"b835",x"3700",x"365a",x"32ee"),
(x"3a98",x"404c",x"3787",x"38c1",x"b811",x"38fb",x"3671",x"329b",x"3ab4",x"405b",x"37b3",x"38ae",x"b826",x"38fc",x"3671",x"3303",x"3abc",x"4053",x"376e",x"38f6",x"b815",x"38c2",x"365a",x"32ce"),
(x"3ab4",x"405b",x"37b3",x"b422",x"b30f",x"3b86",x"359b",x"337d",x"3a98",x"404c",x"3787",x"b776",x"b053",x"3afe",x"359b",x"33e2",x"3aab",x"405b",x"37ae",x"b776",x"b053",x"3afe",x"3594",x"3382"),
(x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db",x"3ab4",x"405b",x"37b3",x"348b",x"3a04",x"38c2",x"3648",x"33ec",x"3aab",x"405b",x"37ae",x"b35e",x"39d9",x"3923",x"3644",x"33e0"),
(x"3aab",x"405b",x"37ae",x"b776",x"b053",x"3afe",x"3594",x"3382",x"3a98",x"404c",x"3787",x"b776",x"b053",x"3afe",x"359b",x"33e2",x"3aa2",x"405b",x"379f",x"b8fe",x"ab38",x"3a3b",x"358c",x"3389"),
(x"3aa2",x"405b",x"379f",x"b54f",x"39c9",x"38d8",x"3642",x"33cf",x"3a94",x"405d",x"3780",x"acce",x"3bc5",x"3334",x"3644",x"33ae",x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db"),
(x"3aae",x"405e",x"3752",x"1d38",x"3bf5",x"2e94",x"365d",x"33ae",x"3acc",x"405e",x"3752",x"324d",x"3bb2",x"31fb",x"366d",x"33ce",x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db"),
(x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db",x"3acc",x"405e",x"3752",x"324d",x"3bb2",x"31fb",x"366d",x"33ce",x"3ac6",x"405d",x"377d",x"3600",x"3ae5",x"3571",x"365f",x"33e0"),
(x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9",x"3a81",x"405c",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"252a",x"3a78",x"405b",x"37da",x"b146",x"3a67",x"389c",x"3659",x"2595"),
(x"3a81",x"405c",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"252a",x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3a9b",x"405b",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"2563"),
(x"3a8a",x"405b",x"37da",x"b950",x"a0dd",x"39fa",x"35c9",x"1fba",x"3a81",x"4057",x"37cb",x"b950",x"a0dd",x"39fa",x"35bc",x"1ee4",x"3a81",x"405c",x"37cb",x"b950",x"a0dd",x"39fa",x"35c9",x"1d62"),
(x"3a78",x"405b",x"37da",x"393c",x"95bc",x"3a0c",x"35e3",x"3069",x"3a81",x"405c",x"37cb",x"393c",x"95bc",x"3a0c",x"35eb",x"305f",x"3a81",x"4057",x"37cb",x"393c",x"95bc",x"3a0c",x"35eb",x"307c"),
(x"3a8a",x"405b",x"37da",x"3325",x"b878",x"3a63",x"35f3",x"28c6",x"3a9b",x"405b",x"37d1",x"333b",x"b811",x"3aa5",x"3600",x"28cc",x"3a81",x"4057",x"37cb",x"9e0a",x"b823",x"3ad8",x"35ed",x"2927"),
(x"3a64",x"404e",x"3791",x"b252",x"b816",x"3ab1",x"35d8",x"2a3e",x"3a62",x"405a",x"37cd",x"b1e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"3a82",x"4051",x"37ad",x"23bb",x"b81b",x"3add",x"35ee",x"29d8"),
(x"3a62",x"405a",x"37cd",x"baf6",x"b475",x"367c",x"362a",x"3154",x"3a64",x"404e",x"3791",x"baf1",x"b416",x"36d1",x"362a",x"31a9",x"3a5e",x"405a",x"37ba",x"bb3a",x"b41e",x"357a",x"3622",x"315a"),
(x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9",x"3a62",x"405a",x"37cd",x"b58a",x"3a1b",x"385c",x"3649",x"253f",x"3a5e",x"405a",x"37ba",x"b926",x"39b7",x"3463",x"3645",x"24cf"),
(x"3a5e",x"405a",x"37ba",x"bb3a",x"b41e",x"357a",x"3622",x"315a",x"3a64",x"404e",x"3791",x"baf1",x"b416",x"36d1",x"362a",x"31a9",x"3a59",x"405b",x"379b",x"baed",x"b3c2",x"36ff",x"3617",x"3165"),
(x"3a59",x"405b",x"379b",x"b825",x"3acf",x"2d30",x"3640",x"2413",x"3a66",x"405c",x"3781",x"b1af",x"3bdf",x"1c18",x"364b",x"22d3",x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"3a94",x"405d",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"22d4",x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9",x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3a81",x"405c",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"252a"),
(x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3a94",x"405d",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"22d4",x"3aa2",x"405b",x"379f",x"394b",x"39eb",x"af9d",x"367a",x"243b"),
(x"3a9b",x"405b",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"2563",x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3aa3",x"405b",x"37ba",x"392f",x"39d8",x"32de",x"367a",x"24e0"),
(x"3a9b",x"405b",x"37d1",x"39f1",x"b5fe",x"3870",x"35a0",x"3460",x"3aa3",x"405b",x"37ba",x"3b76",x"b463",x"3372",x"3596",x"345c",x"3a98",x"404c",x"3787",x"3b76",x"b463",x"3372",x"35a0",x"342c"),
(x"3aa2",x"405b",x"379f",x"3bda",x"afe2",x"b0aa",x"358d",x"3457",x"3a98",x"404c",x"3787",x"3b76",x"b463",x"3372",x"35a0",x"342c",x"3aa3",x"405b",x"37ba",x"3b76",x"b463",x"3372",x"3596",x"345c"),
(x"3a60",x"404e",x"378f",x"b5a5",x"b161",x"3b5d",x"3626",x"31a8",x"3a59",x"405b",x"379b",x"baed",x"b3c3",x"3700",x"3617",x"3165",x"3a64",x"404e",x"3791",x"baf1",x"b416",x"36d1",x"362a",x"31a9"),
(x"3a60",x"404e",x"378f",x"367e",x"ac15",x"3b4b",x"3689",x"3214",x"3a5e",x"404c",x"378e",x"b850",x"b763",x"39a2",x"3686",x"3221",x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"3a3b",x"4052",x"376e",x"b92e",x"b7c8",x"38b1",x"3668",x"3200",x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5",x"3a5e",x"404c",x"378e",x"b850",x"b763",x"39a2",x"3686",x"3221"),
(x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5",x"3a32",x"4057",x"377a",x"b9d3",x"b83b",x"36f5",x"3663",x"31e2",x"3a30",x"405a",x"378b",x"b815",x"b8b5",x"3904",x"3664",x"31ce"),
(x"3a28",x"405b",x"3775",x"ba72",x"b85a",x"3373",x"365a",x"31ce",x"3a32",x"4057",x"377a",x"b9d3",x"b83b",x"36f5",x"3663",x"31e2",x"3a21",x"405c",x"3752",x"ba86",x"b816",x"3455",x"364c",x"31d5"),
(x"3a32",x"405d",x"3780",x"bbd2",x"3047",x"b134",x"35a0",x"1f3a",x"3a32",x"405b",x"3797",x"bb81",x"34c0",x"31b9",x"35aa",x"1ea6",x"3a30",x"405a",x"378b",x"bbd2",x"3048",x"b133",x"35aa",x"2000"),
(x"3a32",x"405d",x"3780",x"b66b",x"ad14",x"3b4c",x"362f",x"31bd",x"3a32",x"4057",x"377a",x"b612",x"af46",x"3b58",x"362f",x"31de",x"3a28",x"405b",x"3775",x"b66b",x"ad14",x"3b4c",x"3626",x"31c9"),
(x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b",x"3a44",x"405a",x"37b0",x"9fc8",x"3964",x"39e8",x"3641",x"2b5a",x"3a32",x"405b",x"3797",x"b553",x"3a2a",x"3858",x"3650",x"2b30"),
(x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b",x"3a60",x"405d",x"3777",x"3179",x"3b46",x"3611",x"3645",x"2c28",x"3a59",x"405b",x"379b",x"35ee",x"392f",x"3951",x"363c",x"2bdc"),
(x"3a59",x"405b",x"379b",x"35ee",x"392f",x"3951",x"363c",x"2bdc",x"3a60",x"405d",x"3777",x"3179",x"3b46",x"3611",x"3645",x"2c28",x"3a66",x"405c",x"3781",x"3106",x"3a66",x"38a1",x"363f",x"2c29"),
(x"3a55",x"405d",x"375d",x"a8bc",x"3bf3",x"2e92",x"3652",x"2c29",x"3a60",x"405d",x"3777",x"3179",x"3b46",x"3611",x"3645",x"2c28",x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b"),
(x"3a2a",x"405d",x"3752",x"b410",x"3b92",x"3261",x"3669",x"2b9b",x"3a2a",x"405c",x"3777",x"b91e",x"39e6",x"32f0",x"365f",x"2b4f",x"3a28",x"405b",x"3775",x"b9b9",x"391a",x"348e",x"3661",x"2b30"),
(x"3a50",x"405e",x"3752",x"a4c2",x"3be9",x"30b5",x"3658",x"2c27",x"3a55",x"405d",x"375d",x"a8bc",x"3bf3",x"2e92",x"3652",x"2c29",x"3a32",x"405d",x"3780",x"ade3",x"3bd5",x"31ce",x"3658",x"2b68"),
(x"3a32",x"405d",x"3780",x"ade3",x"3bd5",x"31ce",x"3658",x"2b68",x"3a2a",x"405c",x"3777",x"b91e",x"39e6",x"32f0",x"365f",x"2b4f",x"3a2a",x"405d",x"3752",x"b410",x"3b92",x"3261",x"3669",x"2b9b"),
(x"3acb",x"3fd8",x"3786",x"3af1",x"b04f",x"37a7",x"3637",x"331f",x"3ac4",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"3639",x"3346",x"3adb",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"361f",x"3321"),
(x"3ac4",x"3fe5",x"378d",x"3a9a",x"3440",x"37f9",x"3639",x"3346",x"3abe",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"363a",x"3356",x"3ad1",x"3fea",x"3752",x"3a66",x"3621",x"3762",x"3620",x"334e"),
(x"3ac9",x"3ff0",x"3752",x"38fd",x"390a",x"3765",x"3622",x"3363",x"3abe",x"3fea",x"378e",x"38b7",x"393a",x"3798",x"363a",x"3356",x"3ac1",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"3624",x"336f"),
(x"3adb",x"3fdb",x"3752",x"3ae6",x"a81b",x"380a",x"361f",x"3321",x"3ac5",x"3fa8",x"3752",x"3afd",x"b17a",x"3748",x"3634",x"328d",x"3acb",x"3fd8",x"3786",x"3af1",x"b04f",x"37a7",x"3637",x"331f"),
(x"3ac5",x"3fa8",x"3752",x"3afd",x"b17a",x"3748",x"3634",x"328d",x"3abd",x"3f8b",x"3752",x"3b0e",x"aeb1",x"3757",x"363e",x"323c",x"3abc",x"3fa7",x"3777",x"3b1d",x"b0f4",x"36e3",x"3643",x"3291"),
(x"3ac1",x"3ff2",x"3752",x"b21b",x"3ba5",x"332f",x"3624",x"336f",x"3aa9",x"3fea",x"378e",x"b8f8",x"3a44",x"1dd6",x"3644",x"3373",x"3aa2",x"3fe5",x"3782",x"b9d9",x"3972",x"a970",x"3645",x"3385"),
(x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3abc",x"3fa7",x"3777",x"ab80",x"ac13",x"3bf8",x"35a9",x"31f0",x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c"),
(x"3abc",x"3fa7",x"3777",x"ab80",x"ac13",x"3bf8",x"35a9",x"31f0",x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3acb",x"3fd8",x"3786",x"282c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"3ac4",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"35a5",x"327f",x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3acb",x"3fd8",x"3786",x"282c",x"ad9c",x"3bf6",x"35a0",x"327f"),
(x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ac4",x"3fe5",x"378d",x"2e28",x"ac9e",x"3bf1",x"35a6",x"32a5"),
(x"3abe",x"3fea",x"378e",x"2da8",x"257a",x"3bf7",x"35ab",x"32b3",x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ab3",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"35b3",x"32b8"),
(x"3ab3",x"3fec",x"378f",x"2231",x"267a",x"3bff",x"35b3",x"32b8",x"3ab2",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"3aa9",x"3fea",x"378e",x"ae38",x"2687",x"3bf5",x"35bc",x"32b1"),
(x"3aa9",x"3fea",x"378e",x"ae38",x"2687",x"3bf5",x"35bc",x"32b1",x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3aa0",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"35c2",x"329a"),
(x"3a9b",x"3fe0",x"378b",x"aefe",x"af3d",x"3be6",x"35c6",x"3293",x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3a9b",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"3aa0",x"3fe2",x"378c",x"ad04",x"a9d6",x"3bf7",x"35c2",x"329a",x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3a9b",x"3fe0",x"378b",x"aefe",x"af3d",x"3be6",x"35c6",x"3293"),
(x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3a9b",x"3fd4",x"3784",x"af9f",x"aede",x"3be5",x"35c6",x"3271"),
(x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3aa4",x"3faa",x"3777",x"2c2f",x"accc",x"3bf5",x"35bc",x"31f5",x"3a9b",x"3fc3",x"377f",x"a7d5",x"ad38",x"3bf8",x"35c4",x"323e"),
(x"3aa4",x"3faa",x"3777",x"2c2f",x"accc",x"3bf5",x"35bc",x"31f5",x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3a9b",x"3fa8",x"3777",x"2bc1",x"ab62",x"3bf8",x"35c2",x"31f0"),
(x"3aa4",x"3faa",x"3777",x"2c2f",x"accc",x"3bf5",x"35bc",x"31f5",x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3aa8",x"3fab",x"3775",x"3235",x"abce",x"3bd5",x"35b8",x"31f9"),
(x"3aa6",x"3fc4",x"3780",x"3042",x"adc4",x"3be5",x"35bd",x"3243",x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245"),
(x"3aa7",x"3fd5",x"3782",x"2e90",x"aed5",x"3be9",x"35bb",x"3274",x"3aa3",x"3fd5",x"3788",x"321a",x"aee2",x"3bce",x"35bf",x"3274",x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293"),
(x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293",x"3aa6",x"3fe0",x"378c",x"3200",x"b152",x"3bbe",x"35be",x"3295",x"3aaf",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"35b6",x"32a0"),
(x"3aaf",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"35b6",x"32a0",x"3aac",x"3fe7",x"378f",x"3000",x"b252",x"3bc7",x"35b9",x"32a9",x"3ab4",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"3ab2",x"3fe9",x"3790",x"9b2b",x"b31f",x"3bcc",x"35b4",x"32ae",x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ab4",x"3fe6",x"3787",x"2981",x"b812",x"3ae0",x"35b3",x"32a3"),
(x"3abb",x"3fe8",x"378f",x"ac4b",x"b2c9",x"3bcc",x"35ad",x"32ab",x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"3ac0",x"3fe3",x"378d",x"b0de",x"b193",x"3bc8",x"35a9",x"329f",x"3ac4",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"35a5",x"327f",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298"),
(x"3ac4",x"3fd8",x"3788",x"b23a",x"add2",x"3bd0",x"35a5",x"327f",x"3ab5",x"3fa9",x"3776",x"b1d8",x"aa80",x"3bda",x"35af",x"31f3",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"3aa8",x"3fab",x"3775",x"3235",x"abce",x"3bd5",x"35b8",x"31f9",x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245",x"3ab1",x"3fa9",x"3773",x"ac3e",x"aa17",x"3bf9",x"35b1",x"31f5"),
(x"3aab",x"3fc5",x"377a",x"2deb",x"ad07",x"3bf0",x"35b8",x"3245",x"3aa7",x"3fd5",x"3782",x"2e90",x"aed5",x"3be9",x"35bb",x"3274",x"3ac0",x"3fd8",x"3782",x"b118",x"ac7e",x"3be0",x"35a9",x"327d"),
(x"3aa7",x"3fd5",x"3782",x"2e90",x"aed5",x"3be9",x"35bb",x"3274",x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293",x"3abc",x"3fe1",x"3785",x"ae7b",x"afec",x"3be5",x"35ac",x"3298"),
(x"3aaa",x"3fe0",x"3787",x"32b9",x"afe5",x"3bc2",x"35ba",x"3293",x"3aaf",x"3fe4",x"3787",x"3503",x"b421",x"3b4f",x"35b6",x"32a0",x"3ab9",x"3fe5",x"3787",x"b09f",x"b24e",x"3bc1",x"35af",x"32a1"),
(x"3a98",x"3fa7",x"378a",x"3bec",x"2581",x"3053",x"35e3",x"3284",x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236",x"3a9a",x"3fa8",x"3783",x"3b1f",x"a907",x"3740",x"35e6",x"3285"),
(x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236",x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205",x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236"),
(x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205",x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203"),
(x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec",x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5"),
(x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1",x"3a93",x"3fe1",x"37b6",x"3a64",x"b8cb",x"29c5",x"35e0",x"31dc",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc",x"3a93",x"3fe1",x"37b6",x"3a64",x"b8cb",x"29c5",x"35e0",x"31dc",x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1",x"3a93",x"3fe1",x"37c1",x"3add",x"b464",x"b6f2",x"35dc",x"31dd",x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0",x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe",x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a99",x"3fc5",x"37c6",x"3af7",x"2fc0",x"b79e",x"35d2",x"322a"),
(x"3a99",x"3fc5",x"37c6",x"3af7",x"2fc0",x"b79e",x"35d2",x"322a",x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e",x"3a99",x"3f8a",x"3790",x"3bff",x"25e3",x"1e73",x"35da",x"32db",x"3a98",x"3fa8",x"37b2",x"3be6",x"a82f",x"30eb",x"35d4",x"327f"),
(x"3a98",x"3fa8",x"37b2",x"3be6",x"a82f",x"30eb",x"35d4",x"327f",x"3a99",x"3fc3",x"37d1",x"3bf3",x"a804",x"2ec5",x"35cd",x"322c",x"3a99",x"3fa8",x"37a7",x"3bb5",x"2cb2",x"b41d",x"35d8",x"327e"),
(x"3a99",x"3fc5",x"37c6",x"3af7",x"2fc0",x"b79e",x"35d2",x"322a",x"3a99",x"3fc3",x"37d1",x"3bf3",x"a804",x"2ec5",x"35cd",x"322c",x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe"),
(x"3a99",x"3fd3",x"37d4",x"3b45",x"2659",x"b6aa",x"35d0",x"31fe",x"3a98",x"3fd3",x"37de",x"3be7",x"9cea",x"30f2",x"35cc",x"31fd",x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0"),
(x"3a99",x"3fde",x"37d2",x"3b61",x"add1",x"b5fd",x"35d3",x"31e0",x"3a98",x"3fdf",x"37dc",x"3bdc",x"28a8",x"31da",x"35d0",x"31db",x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1"),
(x"3a99",x"3fe3",x"37c8",x"3b6f",x"b4b7",x"b314",x"35d9",x"31d1",x"3a99",x"3fe6",x"37cc",x"3bf2",x"2959",x"2ec5",x"35d9",x"31c8",x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"3a9a",x"3fe8",x"37b8",x"3bfd",x"2587",x"2a48",x"35e1",x"31c5",x"3a9a",x"3fe7",x"37a7",x"3bff",x"1ec2",x"2532",x"35e8",x"31ca",x"3a9a",x"3fe6",x"37b7",x"3b9f",x"b4d7",x"2439",x"35e1",x"31cc"),
(x"3a9a",x"3fe7",x"37a7",x"3bff",x"1ec2",x"2532",x"35e8",x"31ca",x"3a9a",x"3fe0",x"378e",x"3bf9",x"1818",x"2d46",x"35f0",x"31e1",x"3a9a",x"3fe4",x"37aa",x"3b36",x"b4f4",x"34d4",x"35e6",x"31d3"),
(x"3a9a",x"3fe0",x"378e",x"3bf9",x"1818",x"2d46",x"35f0",x"31e1",x"3a9b",x"3fd4",x"3784",x"3beb",x"a025",x"3083",x"35f2",x"3204",x"3a9a",x"3fde",x"3799",x"3b18",x"b180",x"36da",x"35ec",x"31e5"),
(x"3a9b",x"3fd4",x"3784",x"3beb",x"a025",x"3083",x"35f2",x"3204",x"3a9b",x"3fc3",x"377f",x"3bd2",x"a2f6",x"32b9",x"35f0",x"3237",x"3a9a",x"3fd4",x"3790",x"3ada",x"acd9",x"3814",x"35ed",x"3203"),
(x"3a9a",x"3fa8",x"3783",x"3b1f",x"a907",x"3740",x"35e6",x"3285",x"3a9a",x"3fc2",x"378b",x"3acd",x"a90b",x"3833",x"35eb",x"3236",x"3a9b",x"3fa8",x"3777",x"3bc7",x"a659",x"336e",x"35eb",x"3285"),
(x"3a97",x"3fa9",x"379f",x"3bfa",x"2c34",x"a7c1",x"35dc",x"327e",x"3a98",x"3fa7",x"378a",x"3bec",x"2581",x"3053",x"35e3",x"3284",x"3a99",x"3f8a",x"3790",x"3bff",x"25e3",x"1e73",x"35da",x"32db"),
(x"3a98",x"3fa7",x"378a",x"3bec",x"2581",x"3053",x"35e3",x"3284",x"3a97",x"3fa9",x"379f",x"3bfa",x"2c34",x"a7c1",x"35dc",x"327e",x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236"),
(x"3a94",x"3fc2",x"3794",x"3bb1",x"2446",x"345f",x"35e6",x"3236",x"3a93",x"3fc5",x"37ba",x"3be1",x"2c8e",x"b0f7",x"35d8",x"3228",x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205"),
(x"3a94",x"3fd3",x"3798",x"3bae",x"a64c",x"3470",x"35e8",x"3205",x"3a93",x"3fd3",x"37c9",x"3bcf",x"2a48",x"b2c7",x"35d6",x"3200",x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec"),
(x"3a93",x"3fdc",x"37a3",x"3bad",x"a9fd",x"346f",x"35e5",x"31ec",x"3a93",x"3fdd",x"37c7",x"3b8c",x"a673",x"b548",x"35d9",x"31e6",x"3a93",x"3fe0",x"37ac",x"3b37",x"b40b",x"359a",x"35e3",x"31e1"),
(x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a98",x"3fa8",x"37b2",x"3870",x"b1f2",x"3a7c",x"35f5",x"3500",x"3a7a",x"3f87",x"37c0",x"a48e",x"b255",x"3bd7",x"35d8",x"352f"),
(x"3a98",x"3fa8",x"37b2",x"3870",x"b1f2",x"3a7c",x"35f5",x"3500",x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a99",x"3fc3",x"37d1",x"3885",x"b324",x"3a5a",x"35f4",x"34d4"),
(x"3a99",x"3fc3",x"37d1",x"3885",x"b324",x"3a5a",x"35f4",x"34d4",x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a98",x"3fd3",x"37de",x"389a",x"ad78",x"3a82",x"35f2",x"34bc"),
(x"3a98",x"3fd3",x"37de",x"389a",x"ad78",x"3a82",x"35f2",x"34bc",x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a98",x"3fdf",x"37dc",x"3869",x"323c",x"3a7d",x"35f0",x"34aa"),
(x"3a98",x"3fdf",x"37dc",x"3869",x"323c",x"3a7d",x"35f0",x"34aa",x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a99",x"3fe6",x"37cc",x"3783",x"398b",x"385f",x"35ef",x"349c"),
(x"3a79",x"3feb",x"37e2",x"9953",x"3ada",x"3821",x"35d7",x"349e",x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495",x"3a99",x"3fe6",x"37cc",x"3783",x"398b",x"385f",x"35ef",x"349c"),
(x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495",x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e",x"3a9a",x"3fe8",x"37b8",x"35d5",x"3b70",x"2a94",x"35f1",x"3494"),
(x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e",x"3a91",x"3fe7",x"379c",x"3620",x"3a0a",x"b841",x"35ed",x"3488",x"3a9a",x"3fe7",x"37a7",x"3572",x"3a96",x"b740",x"35f3",x"348e"),
(x"3aa2",x"3fe5",x"3782",x"b9d9",x"3972",x"a970",x"3645",x"3385",x"3aa0",x"3fe2",x"378c",x"b9d1",x"382c",x"3723",x"364c",x"3387",x"3a9a",x"3fe1",x"3786",x"b88d",x"3867",x"38e2",x"364c",x"3391"),
(x"3a97",x"3fe1",x"378b",x"3994",x"399e",x"b083",x"35f6",x"3480",x"3a9a",x"3fe1",x"3786",x"381b",x"39f5",x"36cf",x"35f8",x"347e",x"3a9a",x"3fe0",x"378e",x"381d",x"395a",x"b849",x"35f9",x"3481"),
(x"3a28",x"3fd8",x"3786",x"bad9",x"b071",x"37f4",x"35c2",x"2e97",x"3a18",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"35ab",x"2e93",x"3a2f",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"35c4",x"2e47"),
(x"3a2f",x"3fe5",x"378d",x"ba9a",x"3440",x"37f9",x"35c4",x"2e47",x"3a22",x"3fea",x"3752",x"ba66",x"3621",x"3762",x"35ab",x"2e39",x"3a35",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"35c6",x"2e27"),
(x"3a40",x"3fec",x"378f",x"28ac",x"3b7d",x"3597",x"35ca",x"2e09",x"3a35",x"3fea",x"378e",x"b8b7",x"393a",x"3798",x"35c6",x"2e27",x"3a33",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"35af",x"2df7"),
(x"3a18",x"3fdb",x"3752",x"bae6",x"a81b",x"380a",x"35ab",x"2e93",x"3a28",x"3fd8",x"3786",x"bad9",x"b071",x"37f4",x"35c2",x"2e97",x"3a2e",x"3fa8",x"3752",x"badc",x"b152",x"37c7",x"35c0",x"2fbb"),
(x"3a2e",x"3fa8",x"3752",x"badc",x"b152",x"37c7",x"35c0",x"2fbb",x"3a38",x"3fa6",x"3775",x"bacd",x"b078",x"380f",x"35cf",x"2fb9",x"3a34",x"3f8b",x"3752",x"bab6",x"ad4f",x"384d",x"35c9",x"302f"),
(x"3a33",x"3ff2",x"3752",x"321b",x"3ba5",x"332f",x"35af",x"2df7",x"3a52",x"3fe5",x"3782",x"39dc",x"3971",x"a62b",x"35d1",x"2dca",x"3a4b",x"3fea",x"378e",x"38f8",x"3a44",x"1dd6",x"35cf",x"2dee"),
(x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2",x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e",x"3a38",x"3fa6",x"3775",x"ab9a",x"acf0",x"3bf6",x"3611",x"30d8"),
(x"3a2f",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"360d",x"3046",x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2",x"3a28",x"3fd8",x"3786",x"ae54",x"ae94",x"3beb",x"3607",x"3046"),
(x"3a2f",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"360d",x"3046",x"3a28",x"3fd8",x"3786",x"ae54",x"ae94",x"3beb",x"3607",x"3046",x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026"),
(x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026",x"3a2f",x"3fe5",x"378d",x"ae28",x"ac9e",x"3bf1",x"360d",x"3020",x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"3a41",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"361b",x"3016",x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a",x"3a40",x"3fec",x"378f",x"a231",x"267a",x"3bff",x"361b",x"300d"),
(x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a41",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"361b",x"3016",x"3a4b",x"3fea",x"378e",x"2e38",x"2687",x"3bf5",x"3623",x"3014"),
(x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f",x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a54",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"3a58",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"362d",x"3032",x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f",x"3a54",x"3fe2",x"378c",x"2d04",x"a9d6",x"3bf7",x"362a",x"302b"),
(x"3a59",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"362d",x"3054",x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051",x"3a58",x"3fe0",x"378b",x"2efe",x"af3d",x"3be6",x"362d",x"3032"),
(x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051",x"3a59",x"3fd4",x"3784",x"2f9f",x"aede",x"3be5",x"362d",x"3054",x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082"),
(x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082",x"3a58",x"3fc3",x"377f",x"27d5",x"ad38",x"3bf8",x"362b",x"3087",x"3a50",x"3faa",x"3777",x"ac34",x"acb0",x"3bf5",x"3623",x"30d0"),
(x"3a50",x"3faa",x"3777",x"ac34",x"acb0",x"3bf5",x"3623",x"30d0",x"3a58",x"3fa8",x"3777",x"a6fd",x"ab9a",x"3bfb",x"3629",x"30d5",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"3a50",x"3faa",x"3777",x"ac34",x"acb0",x"3bf5",x"3623",x"30d0",x"3a4b",x"3fab",x"3775",x"b227",x"ab9d",x"3bd6",x"361f",x"30cb",x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082"),
(x"3a4e",x"3fc4",x"3780",x"b042",x"adc4",x"3be5",x"3624",x"3082",x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080",x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051"),
(x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f",x"3a50",x"3fd5",x"3788",x"b21a",x"aee2",x"3bce",x"3626",x"3051",x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a4e",x"3fe0",x"378c",x"b200",x"b152",x"3bbe",x"3625",x"302f",x"3a44",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"361d",x"3025"),
(x"3a41",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"361b",x"3016",x"3a47",x"3fe7",x"378f",x"b000",x"b252",x"3bc7",x"3620",x"301c",x"3a40",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"361a",x"3022"),
(x"3a41",x"3fe9",x"3790",x"1b2b",x"b31f",x"3bcc",x"361b",x"3016",x"3a40",x"3fe6",x"3787",x"a981",x"b812",x"3ae0",x"361a",x"3022",x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a"),
(x"3a39",x"3fe8",x"378f",x"2c4b",x"b2ca",x"3bcc",x"3615",x"301a",x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026"),
(x"3a34",x"3fe3",x"378d",x"30de",x"b193",x"3bc8",x"3611",x"3026",x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a2f",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"360d",x"3046"),
(x"3a2f",x"3fd8",x"3788",x"323a",x"add2",x"3bd0",x"360d",x"3046",x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a3f",x"3fa9",x"3776",x"2ffb",x"abfc",x"3beb",x"3616",x"30d2"),
(x"3a46",x"3f89",x"376f",x"a217",x"a8a5",x"3bfe",x"3619",x"312e",x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"3a52",x"3f89",x"3770",x"ab4f",x"a8d3",x"3bfb",x"3622",x"312e"),
(x"3a4b",x"3fab",x"3775",x"b227",x"ab9d",x"3bd6",x"361f",x"30cb",x"3a42",x"3fa9",x"3773",x"2c2a",x"a9f3",x"3bf9",x"3618",x"30d0",x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080"),
(x"3a48",x"3fc5",x"377a",x"adeb",x"ad07",x"3bf0",x"361f",x"3080",x"3a33",x"3fd8",x"3782",x"3118",x"ac7e",x"3be0",x"3610",x"3048",x"3a4c",x"3fd5",x"3782",x"ae90",x"aed5",x"3be9",x"3623",x"3050"),
(x"3a4c",x"3fd5",x"3782",x"ae90",x"aed5",x"3be9",x"3623",x"3050",x"3a37",x"3fe1",x"3785",x"2e7a",x"afec",x"3be5",x"3614",x"302d",x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032"),
(x"3a4a",x"3fe0",x"3787",x"b2b9",x"afe5",x"3bc2",x"3621",x"3032",x"3a3b",x"3fe5",x"3787",x"309f",x"b24e",x"3bc1",x"3616",x"3024",x"3a44",x"3fe4",x"3787",x"b503",x"b421",x"3b4f",x"361d",x"3025"),
(x"3a5c",x"3fa8",x"378a",x"bbe0",x"2467",x"319c",x"360d",x"31c3",x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4",x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211",x"3a5a",x"3fc2",x"378b",x"ba70",x"a9d2",x"38bb",x"3615",x"3211",x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242",x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b"),
(x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b",x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263",x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268"),
(x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268",x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a5f",x"3fe2",x"37b7",x"ba93",x"b88d",x"2474",x"360a",x"326f"),
(x"3a5f",x"3fe1",x"37c3",x"bb15",x"b383",x"b669",x"3606",x"326c",x"3a5f",x"3fe2",x"37b7",x"ba93",x"b88d",x"2474",x"360a",x"326f",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277"),
(x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a5f",x"3fe1",x"37c3",x"bb15",x"b383",x"b669",x"3606",x"326c",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a5b",x"3fd3",x"37d2",x"ba75",x"2987",x"b8b5",x"35fc",x"3249"),
(x"3a60",x"3fc5",x"37be",x"bbeb",x"2c4d",x"b006",x"3601",x"321f",x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e"),
(x"3a60",x"3fc5",x"37be",x"bbeb",x"2c4d",x"b006",x"3601",x"321f",x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e",x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9"),
(x"3a5b",x"3fa9",x"37a5",x"bbef",x"2703",x"afed",x"3603",x"31c9",x"3a5b",x"3fa8",x"37b0",x"bbfa",x"a20a",x"2ca3",x"35ff",x"31c8",x"3a5a",x"3f85",x"378d",x"bbff",x"2504",x"1d87",x"3604",x"3160"),
(x"3a5b",x"3fa8",x"37b0",x"bbfa",x"a20a",x"2ca3",x"35ff",x"31c8",x"3a5b",x"3fa9",x"37a5",x"bbef",x"2703",x"afed",x"3603",x"31c9",x"3a5b",x"3fc3",x"37d0",x"bbff",x"a2f6",x"24f0",x"35f8",x"321b"),
(x"3a5b",x"3fc3",x"37d0",x"bbff",x"a2f6",x"24f0",x"35f8",x"321b",x"3a5a",x"3fc4",x"37c6",x"baf8",x"2fc1",x"b79c",x"35fc",x"321e",x"3a5a",x"3fd3",x"37dc",x"bbff",x"15bc",x"a66c",x"35f8",x"324b"),
(x"3a5a",x"3fde",x"37db",x"bbff",x"1953",x"2560",x"35fb",x"326b",x"3a5a",x"3fd3",x"37dc",x"bbff",x"15bc",x"a66c",x"35f8",x"324b",x"3a5b",x"3fdd",x"37d0",x"bb3a",x"ad9b",x"b6b6",x"35ff",x"3266"),
(x"3a5a",x"3fe6",x"37cd",x"bbf7",x"29c5",x"2d1b",x"3603",x"327f",x"3a5a",x"3fde",x"37db",x"bbff",x"1953",x"2560",x"35fb",x"326b",x"3a5a",x"3fe3",x"37c9",x"bb72",x"b453",x"b3d7",x"3604",x"3277"),
(x"3a5a",x"3fe8",x"37b8",x"bbfd",x"1ef6",x"29f0",x"360c",x"3283",x"3a5a",x"3fe6",x"37cd",x"bbf7",x"29c5",x"2d1b",x"3603",x"327f",x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b"),
(x"3a5a",x"3fe8",x"37b8",x"bbfd",x"1ef6",x"29f0",x"360c",x"3283",x"3a5a",x"3fe5",x"37b7",x"bbb2",x"b454",x"25bc",x"360b",x"327b",x"3a5a",x"3fe7",x"37a7",x"bbff",x"0a8d",x"2694",x"3612",x"327d"),
(x"3a5a",x"3fe7",x"37a7",x"bbff",x"0a8d",x"2694",x"3612",x"327d",x"3a5a",x"3fe4",x"37aa",x"bb50",x"b4c5",x"3465",x"3610",x"3274",x"3a59",x"3fe0",x"378e",x"bbf8",x"1553",x"2d82",x"361b",x"3266"),
(x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a59",x"3fd4",x"3784",x"bbea",x"a025",x"3095",x"361c",x"3243",x"3a59",x"3fde",x"3798",x"bb1d",x"b165",x"36cb",x"3617",x"3263"),
(x"3a59",x"3fd4",x"3784",x"bbea",x"a025",x"3095",x"361c",x"3243",x"3a59",x"3fd4",x"3790",x"badf",x"ac91",x"380d",x"3618",x"3244",x"3a58",x"3fc3",x"377f",x"bbce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"3a5a",x"3fc2",x"378b",x"ba70",x"a9d2",x"38bb",x"3615",x"3211",x"3a5a",x"3fa8",x"3782",x"bb3c",x"a8f7",x"36cb",x"3611",x"31c4",x"3a58",x"3fc3",x"377f",x"bbce",x"a3ef",x"32f4",x"361a",x"3210"),
(x"3a5c",x"3fa8",x"378a",x"bbe0",x"2467",x"319c",x"360d",x"31c3",x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9",x"3a5a",x"3f89",x"3770",x"bbf0",x"1d6d",x"2fcb",x"360f",x"3168"),
(x"3a60",x"3fc5",x"37be",x"bbeb",x"2c4d",x"b006",x"3601",x"321f",x"3a5c",x"3fa9",x"37a1",x"bbf1",x"2c5d",x"ae43",x"3605",x"31c9",x"3a5f",x"3fc2",x"3794",x"bbcf",x"24e3",x"32e2",x"3610",x"3211"),
(x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a60",x"3fc5",x"37be",x"bbeb",x"2c4d",x"b006",x"3601",x"321f",x"3a5f",x"3fd3",x"3798",x"bbbc",x"a0a8",x"3410",x"3612",x"3242"),
(x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a60",x"3fd3",x"37c9",x"bbd1",x"2963",x"b2aa",x"3601",x"3246",x"3a60",x"3fdc",x"37a3",x"bbc0",x"accc",x"3386",x"3610",x"325b"),
(x"3a5f",x"3fe1",x"37c3",x"bb15",x"b383",x"b669",x"3606",x"326c",x"3a5f",x"3fdd",x"37c9",x"bb95",x"ac0e",x"b4fe",x"3603",x"3262",x"3a5f",x"3fe0",x"37ac",x"bb6f",x"b421",x"3438",x"360e",x"3268"),
(x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a7a",x"3f87",x"37c0",x"a48e",x"b255",x"3bd7",x"35d8",x"352f",x"3a5b",x"3fa8",x"37b0",x"b87f",x"b1e6",x"3a73",x"35ba",x"3500"),
(x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a79",x"3fa8",x"37dc",x"a217",x"b41e",x"3bba",x"35d7",x"34fc",x"3a5b",x"3fc3",x"37d0",x"b896",x"b2c0",x"3a54",x"35bb",x"34d5"),
(x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a7a",x"3fc7",x"3800",x"a31d",x"b311",x"3bcd",x"35d8",x"34cd",x"3a5a",x"3fd3",x"37dc",x"b892",x"ade1",x"3a86",x"35bc",x"34bc"),
(x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a7a",x"3fd7",x"3804",x"a194",x"28d6",x"3bfe",x"35d8",x"34b8",x"3a5a",x"3fde",x"37db",x"b885",x"3126",x"3a79",x"35be",x"34ab"),
(x"3a79",x"3feb",x"37e2",x"9953",x"3ada",x"3821",x"35d7",x"349e",x"3a79",x"3fe6",x"37fd",x"a12b",x"36f9",x"3b33",x"35d7",x"34a8",x"3a5a",x"3fe6",x"37cd",x"b7e6",x"396d",x"385a",x"35bf",x"349d"),
(x"3a79",x"3feb",x"37e2",x"9953",x"3ada",x"3821",x"35d7",x"349e",x"3a5a",x"3fe6",x"37cd",x"b7e6",x"396d",x"385a",x"35bf",x"349d",x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495"),
(x"3a79",x"3fee",x"37c9",x"9b5f",x"3bbd",x"340d",x"35d7",x"3495",x"3a5a",x"3fe8",x"37b8",x"b61b",x"3b60",x"2bbe",x"35be",x"3495",x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e"),
(x"3a79",x"3fee",x"37b3",x"a9ed",x"3baa",x"b482",x"35d7",x"348e",x"3a5a",x"3fe7",x"37a7",x"b619",x"3a76",x"b730",x"35bb",x"348f",x"3a61",x"3fe4",x"3789",x"b646",x"3a25",x"b80b",x"35bd",x"3481"),
(x"3a52",x"3fe5",x"3782",x"39dc",x"3971",x"a62b",x"35d1",x"2dca",x"3a5b",x"3fe1",x"3782",x"38d3",x"3873",x"3892",x"35d6",x"2daa",x"3a54",x"3fe2",x"378c",x"39bb",x"383c",x"3743",x"35d7",x"2dc5"),
(x"3a5b",x"3fe1",x"3782",x"b865",x"3aa9",x"2c25",x"35b6",x"347e",x"3a5d",x"3fe1",x"378b",x"b8bd",x"3a6d",x"2c06",x"35b7",x"3482",x"3a58",x"3fe0",x"378b",x"b862",x"3a94",x"30e6",x"35b3",x"3481"),
(x"3a39",x"3f6f",x"3752",x"bae4",x"ad23",x"3802",x"35d2",x"307e",x"3a34",x"3f8b",x"3752",x"bab6",x"ad4f",x"384c",x"35c9",x"302f",x"3a3e",x"3f7e",x"376e",x"babb",x"aad9",x"384d",x"35d9",x"3052"),
(x"3a3e",x"3f7e",x"376e",x"b12d",x"203f",x"3be4",x"3613",x"314f",x"3a3f",x"3f88",x"376d",x"b03d",x"a8e0",x"3bec",x"3614",x"3130",x"3a48",x"3f83",x"3770",x"ae2b",x"280b",x"3bf5",x"361a",x"3141"),
(x"3ab9",x"3f6e",x"3752",x"3b03",x"aae6",x"37a4",x"3646",x"31e8",x"3ab3",x"3f7a",x"376e",x"3b00",x"aaa4",x"37b3",x"364e",x"320e",x"3abd",x"3f8b",x"3752",x"3b0e",x"aeb1",x"3757",x"363e",x"323c"),
(x"3aa2",x"3f8b",x"3770",x"2c6c",x"a8e0",x"3bf9",x"35bb",x"319c",x"3aae",x"3f8b",x"376f",x"0cea",x"a7e2",x"3bfe",x"35b2",x"319c",x"3aa2",x"3f7f",x"3770",x"2938",x"1b93",x"3bfe",x"35ba",x"3179"),
(x"3ab4",x"4030",x"37b3",x"348b",x"3a03",x"38c2",x"3611",x"2fda",x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9",x"3ac7",x"4030",x"3794",x"3663",x"3a38",x"37c6",x"3623",x"2fe3"),
(x"3ad7",x"4031",x"3752",x"3890",x"3a28",x"3491",x"363e",x"2fc0",x"3ad0",x"4030",x"377a",x"3864",x"3a40",x"34bc",x"3630",x"2fdb",x"3acc",x"4033",x"3752",x"324d",x"3bb2",x"31fb",x"3638",x"2fa0"),
(x"3ac4",x"4028",x"3752",x"3aa2",x"b726",x"355e",x"363e",x"341a",x"3ac4",x"402c",x"377c",x"39ed",x"b7fd",x"372e",x"364a",x"3429",x"3ad7",x"4031",x"3752",x"3a9b",x"b7a9",x"34c3",x"3635",x"3436"),
(x"3abc",x"4027",x"376e",x"38ec",x"b7ef",x"38e6",x"364a",x"3418",x"3ac4",x"402c",x"377c",x"39ed",x"b7fd",x"372e",x"364a",x"3429",x"3ac4",x"4028",x"3752",x"3aa2",x"b726",x"355e",x"363e",x"341a"),
(x"3ac4",x"402c",x"377c",x"39ed",x"b7fd",x"372e",x"364a",x"3429",x"3ab4",x"4030",x"37b3",x"389d",x"b810",x"391d",x"3662",x"3434",x"3ac7",x"4030",x"3794",x"3839",x"b89f",x"38fa",x"3650",x"3436"),
(x"3abc",x"4027",x"376e",x"38ec",x"b7ef",x"38e6",x"364a",x"3418",x"3ab4",x"4030",x"37b3",x"389d",x"b810",x"391d",x"3662",x"3434",x"3ac4",x"402c",x"377c",x"39ed",x"b7fd",x"372e",x"364a",x"3429"),
(x"3aab",x"4030",x"37ae",x"b35d",x"39d9",x"3923",x"360d",x"2fc2",x"3aa2",x"4031",x"379f",x"b54f",x"39c9",x"38d8",x"360b",x"2fa1",x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"3a94",x"4033",x"3780",x"acce",x"3bc5",x"3335",x"360d",x"2f61",x"3aae",x"4033",x"3752",x"1d38",x"3bf5",x"2e94",x"3627",x"2f61",x"3ab0",x"4032",x"37a2",x"2b55",x"3bb1",x"344c",x"3615",x"2fb9"),
(x"3a62",x"4030",x"37cd",x"b58a",x"3a1b",x"385c",x"3649",x"3358",x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349",x"3a78",x"4030",x"37da",x"b146",x"3a67",x"389c",x"3659",x"3362"),
(x"3a8a",x"4030",x"37da",x"2e09",x"3b05",x"3784",x"3667",x"3363",x"3a81",x"4031",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"3355",x"3a9b",x"4030",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"335c"),
(x"3a98",x"4021",x"3787",x"3409",x"b819",x"3a90",x"3689",x"3140",x"3a82",x"4026",x"37ad",x"23bb",x"b81b",x"3add",x"3677",x"311b",x"3a9b",x"4030",x"37d1",x"333b",x"b811",x"3aa5",x"3689",x"30d9"),
(x"3a81",x"402d",x"37cb",x"9e0a",x"b823",x"3ad8",x"3676",x"30ef",x"3a9b",x"4030",x"37d1",x"333b",x"b811",x"3aa5",x"3689",x"30d9",x"3a82",x"4026",x"37ad",x"23bb",x"b81b",x"3add",x"3677",x"311b"),
(x"3a81",x"402d",x"37cb",x"9e0a",x"b823",x"3ad8",x"3676",x"30ef",x"3a62",x"4030",x"37cd",x"b1e7",x"b81a",x"3ab5",x"365e",x"30e1",x"3a78",x"4030",x"37da",x"b24d",x"b8ad",x"3a4b",x"366f",x"30d9"),
(x"3a82",x"4026",x"37ad",x"23bb",x"b81b",x"3add",x"3677",x"311b",x"3a62",x"4030",x"37cd",x"b1e7",x"b81a",x"3ab5",x"365e",x"30e1",x"3a81",x"402d",x"37cb",x"9e0a",x"b823",x"3ad8",x"3676",x"30ef"),
(x"3a5e",x"4030",x"37ba",x"b926",x"39b7",x"3463",x"3645",x"334a",x"3a59",x"4030",x"379b",x"b825",x"3acf",x"2d30",x"3640",x"3332",x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"3a66",x"4032",x"3781",x"b1af",x"3bdf",x"1bfc",x"364b",x"331d",x"3a94",x"4033",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"331d",x"3a67",x"4032",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"3349"),
(x"3aa3",x"4030",x"37ba",x"392f",x"39d8",x"32de",x"367a",x"334c",x"3a9d",x"4032",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"3343",x"3aa2",x"4031",x"379f",x"394b",x"39eb",x"af9d",x"367a",x"3337"),
(x"3a44",x"4030",x"37b0",x"b5ad",x"b6ed",x"3aa0",x"3659",x"3502",x"3a59",x"4030",x"379b",x"365b",x"ac2a",x"3b52",x"366b",x"3506",x"3a5e",x"4021",x"378e",x"b4a7",x"b630",x"3b00",x"3668",x"3531"),
(x"3a58",x"4021",x"377f",x"b92b",x"b843",x"385f",x"3662",x"3532",x"3a3b",x"4028",x"376e",x"b92f",x"b7c9",x"38af",x"3649",x"3520",x"3a5e",x"4021",x"378e",x"b4a7",x"b630",x"3b00",x"3668",x"3531"),
(x"3a44",x"4030",x"37b0",x"b5ad",x"b6ed",x"3aa0",x"3659",x"3502",x"3a30",x"402f",x"378b",x"b815",x"b8b5",x"3904",x"3646",x"3507",x"3a32",x"4030",x"3797",x"b810",x"b8bd",x"3900",x"3649",x"3503"),
(x"3a3b",x"4028",x"376e",x"b92f",x"b7c9",x"38af",x"3649",x"3520",x"3a32",x"402c",x"377a",x"b9d4",x"b83f",x"36e9",x"3645",x"3511",x"3a44",x"4030",x"37b0",x"b5ad",x"b6ed",x"3aa0",x"3659",x"3502"),
(x"3a35",x"4029",x"3752",x"ba92",x"b7fc",x"346b",x"363e",x"3522",x"3a32",x"402c",x"377a",x"b9d4",x"b83f",x"36e9",x"3645",x"3511",x"3a3b",x"4028",x"376e",x"b92f",x"b7c9",x"38af",x"3649",x"3520"),
(x"3a21",x"4031",x"3752",x"ba84",x"b81e",x"3444",x"362e",x"350b",x"3a32",x"402c",x"377a",x"b9d4",x"b83f",x"36e9",x"3645",x"3511",x"3a35",x"4029",x"3752",x"ba92",x"b7fc",x"346b",x"363e",x"3522"),
(x"3a32",x"402c",x"377a",x"bb82",x"286d",x"b57a",x"35ac",x"20d4",x"3a32",x"4032",x"3780",x"bbd2",x"3047",x"b134",x"35bb",x"2006",x"3a30",x"402f",x"378b",x"bbd2",x"3047",x"b133",x"35b6",x"210c"),
(x"3a2a",x"4032",x"3777",x"b827",x"3037",x"3ac1",x"3628",x"31e5",x"3a32",x"4032",x"3780",x"b66c",x"ad14",x"3b4c",x"362f",x"31e1",x"3a28",x"4030",x"3775",x"b66c",x"ad14",x"3b4c",x"3626",x"31ed"),
(x"3a32",x"4032",x"3780",x"ade3",x"3bd5",x"31ce",x"3625",x"2e26",x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f",x"3a32",x"4030",x"3797",x"b553",x"3a2a",x"3858",x"361e",x"2e0a"),
(x"3a44",x"4030",x"37b0",x"9fc8",x"3964",x"39e8",x"360f",x"2e1f",x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f",x"3a59",x"4030",x"379b",x"35ee",x"392f",x"3951",x"3609",x"2e60"),
(x"3a32",x"4032",x"3780",x"ade3",x"3bd5",x"31ce",x"3625",x"2e26",x"3a55",x"4033",x"375d",x"a8bc",x"3bf3",x"2e92",x"361f",x"2e9b",x"3a49",x"4032",x"37a0",x"91bc",x"3b79",x"35b5",x"3613",x"2e3f"),
(x"3a21",x"4031",x"3752",x"b8c8",x"39c1",x"35a4",x"363b",x"2e1f",x"3a2a",x"4033",x"3752",x"b410",x"3b92",x"3261",x"3637",x"2e3f",x"3a28",x"4030",x"3775",x"b9b9",x"391a",x"348e",x"362e",x"2e0a"),
(x"3a2a",x"4033",x"3752",x"b410",x"3b92",x"3261",x"3637",x"2e3f",x"3a50",x"4033",x"3752",x"a4bc",x"3be9",x"30b5",x"3625",x"2e99",x"3a32",x"4032",x"3780",x"ade3",x"3bd5",x"31ce",x"3625",x"2e26"),
(x"3ab4",x"405b",x"37b3",x"348b",x"3a04",x"38c2",x"3648",x"33ec",x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db",x"3ac7",x"405b",x"3794",x"3663",x"3a38",x"37c6",x"3659",x"33f1"),
(x"3ad7",x"405c",x"3752",x"3890",x"3a28",x"3491",x"3673",x"33df",x"3ad0",x"405b",x"377a",x"3865",x"3a40",x"34bc",x"3665",x"33ed",x"3acc",x"405e",x"3752",x"324d",x"3bb2",x"31fb",x"366d",x"33ce"),
(x"3ac4",x"4054",x"3752",x"3a92",x"b7a6",x"34f5",x"364e",x"32d1",x"3ac4",x"4057",x"377c",x"39d5",x"b835",x"3700",x"365a",x"32ee",x"3ad7",x"405c",x"3752",x"3a92",x"b7f9",x"346d",x"3646",x"3307"),
(x"3abc",x"4053",x"376e",x"38f6",x"b815",x"38c2",x"365a",x"32ce",x"3ac4",x"4057",x"377c",x"39d5",x"b835",x"3700",x"365a",x"32ee",x"3ac4",x"4054",x"3752",x"3a92",x"b7a6",x"34f5",x"364e",x"32d1"),
(x"3ac4",x"4057",x"377c",x"39d5",x"b835",x"3700",x"365a",x"32ee",x"3ab4",x"405b",x"37b3",x"38ae",x"b826",x"38fc",x"3671",x"3303",x"3ac7",x"405b",x"3794",x"3839",x"b89f",x"38fa",x"3660",x"3309"),
(x"3abc",x"4053",x"376e",x"38f6",x"b815",x"38c2",x"365a",x"32ce",x"3ab4",x"405b",x"37b3",x"38ae",x"b826",x"38fc",x"3671",x"3303",x"3ac4",x"4057",x"377c",x"39d5",x"b835",x"3700",x"365a",x"32ee"),
(x"3aab",x"405b",x"37ae",x"b35e",x"39d9",x"3923",x"3644",x"33e0",x"3aa2",x"405b",x"379f",x"b54f",x"39c9",x"38d8",x"3642",x"33cf",x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db"),
(x"3a94",x"405d",x"3780",x"acce",x"3bc5",x"3334",x"3644",x"33ae",x"3aae",x"405e",x"3752",x"1d38",x"3bf5",x"2e94",x"365d",x"33ae",x"3ab0",x"405d",x"37a2",x"2b55",x"3bb1",x"344b",x"364b",x"33db"),
(x"3a62",x"405a",x"37cd",x"b58a",x"3a1b",x"385c",x"3649",x"253f",x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9",x"3a78",x"405b",x"37da",x"b146",x"3a67",x"389c",x"3659",x"2595"),
(x"3a8a",x"405b",x"37da",x"2e09",x"3b05",x"3784",x"3667",x"2596",x"3a81",x"405c",x"37cb",x"2393",x"3b79",x"35b2",x"3660",x"252a",x"3a9b",x"405b",x"37d1",x"31ec",x"3b16",x"36cd",x"3674",x"2563"),
(x"3a98",x"404c",x"3787",x"3409",x"b819",x"3a90",x"3600",x"2a6b",x"3a82",x"4051",x"37ad",x"23bb",x"b81b",x"3add",x"35ee",x"29d8",x"3a9b",x"405b",x"37d1",x"333b",x"b811",x"3aa5",x"3600",x"28cc"),
(x"3a81",x"4057",x"37cb",x"9e0a",x"b823",x"3ad8",x"35ed",x"2927",x"3a9b",x"405b",x"37d1",x"333b",x"b811",x"3aa5",x"3600",x"28cc",x"3a82",x"4051",x"37ad",x"23bb",x"b81b",x"3add",x"35ee",x"29d8"),
(x"3a81",x"4057",x"37cb",x"9e0a",x"b823",x"3ad8",x"35ed",x"2927",x"3a62",x"405a",x"37cd",x"b1e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"3a78",x"405b",x"37da",x"b24d",x"b8ad",x"3a4b",x"35e6",x"28d0"),
(x"3a82",x"4051",x"37ad",x"23bb",x"b81b",x"3add",x"35ee",x"29d8",x"3a62",x"405a",x"37cd",x"b1e7",x"b81a",x"3ab5",x"35d5",x"28ec",x"3a81",x"4057",x"37cb",x"9e0a",x"b823",x"3ad8",x"35ed",x"2927"),
(x"3a5e",x"405a",x"37ba",x"b926",x"39b7",x"3463",x"3645",x"24cf",x"3a59",x"405b",x"379b",x"b825",x"3acf",x"2d30",x"3640",x"2413",x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"3a66",x"405c",x"3781",x"b1af",x"3bdf",x"1c18",x"364b",x"22d3",x"3a94",x"405d",x"3780",x"16f6",x"3bfe",x"27c1",x"366e",x"22d4",x"3a67",x"405c",x"37bd",x"b0a0",x"3bd5",x"3081",x"364d",x"24c9"),
(x"3aa3",x"405b",x"37ba",x"392f",x"39d8",x"32de",x"367a",x"24e0",x"3a9d",x"405d",x"37b1",x"2f93",x"3bda",x"30c0",x"3674",x"249a",x"3aa2",x"405b",x"379f",x"394b",x"39eb",x"af9d",x"367a",x"243b"),
(x"3a59",x"405b",x"379b",x"3713",x"a8bc",x"3b2b",x"3689",x"31cb",x"3a60",x"404e",x"378f",x"367f",x"ac15",x"3b4a",x"3689",x"3214",x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"3a58",x"404c",x"377f",x"b92b",x"b843",x"385f",x"3680",x"3225",x"3a3b",x"4052",x"376e",x"b92e",x"b7c8",x"38b1",x"3668",x"3200",x"3a5e",x"404c",x"378e",x"b850",x"b763",x"39a2",x"3686",x"3221"),
(x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5",x"3a30",x"405a",x"378b",x"b815",x"b8b5",x"3904",x"3664",x"31ce",x"3a32",x"405b",x"3797",x"b810",x"b8bd",x"3900",x"3668",x"31c5"),
(x"3a3b",x"4052",x"376e",x"b92e",x"b7c8",x"38b1",x"3668",x"3200",x"3a32",x"4057",x"377a",x"b9d3",x"b83b",x"36f5",x"3663",x"31e2",x"3a44",x"405a",x"37b0",x"b564",x"b6bf",x"3abb",x"3678",x"31c5"),
(x"3a35",x"4053",x"3752",x"ba90",x"b7ee",x"348a",x"365c",x"3204",x"3a32",x"4057",x"377a",x"b9d3",x"b83b",x"36f5",x"3663",x"31e2",x"3a3b",x"4052",x"376e",x"b92e",x"b7c8",x"38b1",x"3668",x"3200"),
(x"3a21",x"405c",x"3752",x"ba86",x"b816",x"3455",x"364c",x"31d5",x"3a32",x"4057",x"377a",x"b9d3",x"b83b",x"36f5",x"3663",x"31e2",x"3a35",x"4053",x"3752",x"ba90",x"b7ee",x"348a",x"365c",x"3204"),
(x"3a32",x"4057",x"377a",x"bb82",x"286d",x"b57a",x"35aa",x"214e",x"3a32",x"405d",x"3780",x"bbd2",x"3047",x"b134",x"35a0",x"1f3a",x"3a30",x"405a",x"378b",x"bbd2",x"3048",x"b133",x"35aa",x"2000"),
(x"3a2a",x"405c",x"3777",x"b827",x"3037",x"3ac1",x"3628",x"31c1",x"3a32",x"405d",x"3780",x"b66b",x"ad14",x"3b4c",x"362f",x"31bd",x"3a28",x"405b",x"3775",x"b66b",x"ad14",x"3b4c",x"3626",x"31c9"),
(x"3a32",x"405d",x"3780",x"ade3",x"3bd5",x"31ce",x"3658",x"2b68",x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b",x"3a32",x"405b",x"3797",x"b553",x"3a2a",x"3858",x"3650",x"2b30"),
(x"3a44",x"405a",x"37b0",x"9fc8",x"3964",x"39e8",x"3641",x"2b5a",x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b",x"3a59",x"405b",x"379b",x"35ee",x"392f",x"3951",x"363c",x"2bdc"),
(x"3a32",x"405d",x"3780",x"ade3",x"3bd5",x"31ce",x"3658",x"2b68",x"3a55",x"405d",x"375d",x"a8bc",x"3bf3",x"2e92",x"3652",x"2c29",x"3a49",x"405d",x"37a0",x"91bc",x"3b79",x"35b5",x"3646",x"2b9b"),
(x"3a21",x"405c",x"3752",x"b8c8",x"39c1",x"35a4",x"366e",x"2b5b",x"3a2a",x"405d",x"3752",x"b410",x"3b92",x"3261",x"3669",x"2b9b",x"3a28",x"405b",x"3775",x"b9b9",x"391a",x"348e",x"3661",x"2b30"),
(x"3a2a",x"405d",x"3752",x"b410",x"3b92",x"3261",x"3669",x"2b9b",x"3a50",x"405e",x"3752",x"a4c2",x"3be9",x"30b5",x"3658",x"2c27",x"3a32",x"405d",x"3780",x"ade3",x"3bd5",x"31ce",x"3658",x"2b68"),
(x"3adf",x"407a",x"3752",x"375e",x"39fd",x"37a1",x"355f",x"334f",x"3a81",x"407a",x"3802",x"375e",x"39fd",x"37a1",x"34fe",x"334f",x"3a81",x"4088",x"3752",x"375e",x"39fd",x"37a1",x"352a",x"32d0"),
(x"3a50",x"4072",x"3752",x"b9fd",x"0000",x"394d",x"35ef",x"2c07",x"3a80",x"4072",x"37be",x"b9fd",x"0000",x"394d",x"3625",x"2c04",x"3a80",x"405c",x"37be",x"b9fd",x"0000",x"394d",x"3625",x"2d00"),
(x"3ab1",x"405e",x"3752",x"39ee",x"0a8d",x"395e",x"360a",x"2d16",x"3a80",x"405c",x"37be",x"39ee",x"068d",x"395e",x"3641",x"2d01",x"3a80",x"4072",x"37be",x"39ee",x"0a8d",x"395e",x"3641",x"2dfd"),
(x"3a81",x"407a",x"3802",x"3837",x"b940",x"3851",x"35b4",x"2aa4",x"3adf",x"407a",x"3752",x"37fd",x"b973",x"3847",x"3615",x"2aa4",x"3ab1",x"4071",x"3752",x"3837",x"b940",x"3851",x"35fc",x"2bb2"),
(x"3a50",x"4072",x"3752",x"b854",x"b926",x"3853",x"3516",x"34a2",x"3a23",x"407a",x"3752",x"b80d",x"b969",x"3846",x"34fe",x"3480",x"3a81",x"407a",x"3802",x"b854",x"b926",x"3853",x"355f",x"3481"),
(x"3a81",x"407a",x"3802",x"b74c",x"3a02",x"37a3",x"3537",x"2c1c",x"3a23",x"407a",x"3752",x"b74c",x"3a02",x"37a3",x"3597",x"2c08",x"3a81",x"4088",x"3752",x"b74c",x"3a02",x"37a3",x"3566",x"2d0f"),
(x"3ab7",x"3f49",x"3754",x"3ab7",x"9f2b",x"3858",x"34ae",x"259c",x"3ab6",x"3dc2",x"3752",x"3aa2",x"935f",x"3878",x"34ae",x"3122",x"3a79",x"3dc3",x"3804",x"3ab6",x"9af6",x"385a",x"345b",x"311f"),
(x"3a3b",x"3f46",x"3755",x"babd",x"9ffc",x"384e",x"34af",x"25db",x"3a77",x"3f4b",x"380f",x"bad7",x"a310",x"3824",x"3507",x"2563",x"3a79",x"3dc3",x"3804",x"babc",x"9c9b",x"3850",x"3507",x"311e"),
(x"3a53",x"3f7c",x"37bc",x"bad1",x"ab2e",x"3828",x"34d9",x"1b5d",x"3a77",x"3f4b",x"380f",x"bad7",x"a310",x"3824",x"3507",x"2563",x"3a3b",x"3f46",x"3755",x"babd",x"9ffc",x"384e",x"34af",x"25db"),
(x"3ab7",x"3f49",x"3754",x"3ab7",x"9f2b",x"3858",x"34ae",x"259c",x"3a77",x"3f4b",x"380f",x"3ac7",x"a217",x"383e",x"3455",x"2566",x"3a9e",x"3f7c",x"37bb",x"3ac2",x"abcb",x"383f",x"3483",x"1b5d"),
(x"3ade",x"3db3",x"3752",x"38d1",x"395c",x"36f1",x"348c",x"3524",x"3a78",x"3db1",x"3832",x"3904",x"38e5",x"37b5",x"350c",x"3524",x"3a79",x"3dc3",x"3804",x"38d1",x"395c",x"36f1",x"34f0",x"3544"),
(x"3a79",x"3dc3",x"3804",x"b8d0",x"395f",x"36e9",x"3493",x"3520",x"3a78",x"3db1",x"3832",x"b8f7",x"3907",x"377c",x"3477",x"3500",x"3a14",x"3db3",x"3752",x"b8d0",x"395f",x"36e9",x"34f7",x"3500"),
(x"3ade",x"3d4c",x"3752",x"3a6d",x"1c32",x"38c3",x"3512",x"263e",x"3a78",x"3d16",x"3834",x"3a6e",x"1cd0",x"38c1",x"358f",x"1ca0",x"3a78",x"3db1",x"3832",x"3a6d",x"1bfc",x"38c3",x"358f",x"2bd9"),
(x"3a78",x"3db1",x"3832",x"ba6f",x"1d6d",x"38c0",x"3587",x"3369",x"3a78",x"3d16",x"3834",x"ba6b",x"191e",x"38c5",x"3587",x"3495",x"3a11",x"3d4d",x"3752",x"ba6f",x"1d53",x"38c0",x"3505",x"3446"),
(x"3adc",x"3cfb",x"3871",x"2581",x"3a1a",x"392b",x"359d",x"2239",x"3a78",x"3d16",x"3834",x"9c67",x"3a22",x"3922",x"35eb",x"26d8",x"3ade",x"3d4c",x"3752",x"28f7",x"3a35",x"3909",x"359e",x"2b69"),
(x"3a78",x"3d16",x"3834",x"9c67",x"3a22",x"3922",x"35eb",x"26d8",x"3a14",x"3cfa",x"3872",x"a7ce",x"3a15",x"3930",x"3638",x"221d",x"3a11",x"3d4d",x"3752",x"a9e6",x"3a2c",x"3912",x"3638",x"2b6a"),
(x"3a14",x"3cfa",x"3872",x"a7ce",x"3a15",x"3930",x"3638",x"221d",x"3a78",x"3d16",x"3834",x"9c67",x"3a22",x"3922",x"35eb",x"26d8",x"3adc",x"3cfb",x"3871",x"2581",x"3a1a",x"392b",x"359d",x"2239"),
(x"3ade",x"3d4c",x"3752",x"3bff",x"1b5f",x"2393",x"3514",x"304b",x"3ae0",x"3ca2",x"3752",x"3bff",x"1b5f",x"2393",x"3514",x"323a",x"3adc",x"3cfb",x"3871",x"3bff",x"1b5f",x"2393",x"35aa",x"3137"),
(x"3a14",x"3cfa",x"3872",x"1b93",x"b9fb",x"394f",x"34fa",x"34f8",x"3adc",x"3cfb",x"3871",x"1ef6",x"b9f8",x"3952",x"345f",x"34f8",x"3ae0",x"3ca2",x"3752",x"1b93",x"b9fc",x"394f",x"345f",x"3435"),
(x"3a11",x"3d4d",x"3752",x"bbff",x"928d",x"2425",x"35a1",x"310e",x"3a14",x"3cfa",x"3872",x"bbff",x"928d",x"2425",x"350a",x"301f",x"3a11",x"3ca2",x"3752",x"bbff",x"928d",x"2425",x"35a1",x"2e3b"),
(x"3ade",x"3520",x"3752",x"3c00",x"168d",x"9a24",x"350d",x"2ff1",x"3adf",x"30ed",x"3752",x"3c00",x"168d",x"9a24",x"350e",x"2c14",x"3adf",x"3396",x"3874",x"3c00",x"168d",x"9a24",x"35a6",x"2e06"),
(x"3a12",x"351b",x"3752",x"8e8d",x"3a2a",x"3918",x"34fa",x"32b2",x"3ade",x"3520",x"3752",x"a05a",x"3a22",x"3922",x"3460",x"32b2",x"3adf",x"3396",x"3874",x"8e8d",x"3a2a",x"3918",x"3461",x"3131"),
(x"3adf",x"3396",x"3874",x"168d",x"ba26",x"391d",x"3465",x"3428",x"3adf",x"30ed",x"3752",x"991e",x"ba22",x"3922",x"3464",x"32c1",x"3a12",x"30ef",x"3752",x"16f6",x"ba26",x"391d",x"34f9",x"32bf"),
(x"3a12",x"351b",x"3752",x"bc00",x"11bc",x"205a",x"3593",x"317b",x"3a14",x"3397",x"3877",x"bc00",x"11bc",x"205a",x"34ff",x"3271",x"3a12",x"30ef",x"3752",x"bc00",x"11bc",x"205a",x"359b",x"336c"),
(x"3acd",x"401f",x"3786",x"3af9",x"ae2b",x"37ad",x"3620",x"344a",x"3ac7",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3622",x"3459",x"3ad3",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"360a",x"345b"),
(x"3ac7",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3622",x"3459",x"3ac1",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3624",x"3460",x"3acb",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"360c",x"3464"),
(x"3ac1",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3624",x"3460",x"3ab6",x"4027",x"378f",x"a731",x"3bb3",x"3450",x"3628",x"3467",x"3ac3",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"360e",x"346a"),
(x"3ac7",x"400d",x"3752",x"3ae9",x"b336",x"3733",x"361b",x"3412",x"3abe",x"400d",x"3777",x"3b0c",x"b28a",x"36d3",x"362a",x"3414",x"3acd",x"401f",x"3786",x"3af9",x"ae2b",x"37ad",x"3620",x"344a"),
(x"3abf",x"4002",x"3752",x"3b07",x"b070",x"374f",x"3623",x"33e8",x"3ab7",x"4002",x"376d",x"3af0",x"b0d8",x"3796",x"362f",x"33e9",x"3abe",x"400d",x"3777",x"3b0c",x"b28a",x"36d3",x"362a",x"3414"),
(x"3ac3",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"360e",x"346a",x"3ab6",x"4027",x"378f",x"a731",x"3bb3",x"3450",x"3628",x"3467",x"3aab",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"362c",x"346e"),
(x"3aab",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"362c",x"346e",x"3aa2",x"4023",x"378c",x"b949",x"390d",x"367c",x"3632",x"3477",x"3aa4",x"4024",x"3782",x"b904",x"3a39",x"a8ac",x"362c",x"3476"),
(x"3abe",x"400d",x"3777",x"1d6d",x"aedf",x"3bf4",x"3578",x"34f2",x"3ab7",x"4002",x"376d",x"2fac",x"ad49",x"3bea",x"357c",x"34d1",x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3acd",x"401f",x"3786",x"30fd",x"b013",x"3bd6",x"356f",x"3528",x"3abe",x"400d",x"3777",x"1d6d",x"aedf",x"3bf4",x"3578",x"34f2"),
(x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3ac7",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3575",x"3536"),
(x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3ac1",x"4026",x"378e",x"2d5c",x"a074",x"3bf8",x"357a",x"353b"),
(x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3ab6",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3582",x"353d"),
(x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3aaf",x"4025",x"378f",x"317b",x"b4aa",x"3b87",x"3587",x"3537",x"3aab",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aa2",x"4023",x"378c",x"a87a",x"ad2b",x"3bf8",x"3591",x"3531",x"3aab",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"3a9d",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3594",x"352f",x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aa6",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"358e",x"3523"),
(x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3a9e",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"3593",x"350f",x"3a9d",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"3aa6",x"400e",x"3777",x"2c2d",x"ae61",x"3bf1",x"358b",x"34f3",x"3a9d",x"400d",x"3777",x"2bbe",x"acea",x"3bf6",x"3591",x"34f1",x"3a9e",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"3593",x"350f"),
(x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3a9c",x"3fff",x"3770",x"2e76",x"a942",x"3bf3",x"3590",x"34c9",x"3a9d",x"400d",x"3777",x"2bbe",x"acea",x"3bf6",x"3591",x"34f1"),
(x"3aa6",x"400e",x"3777",x"2c2d",x"ae61",x"3bf1",x"358b",x"34f3",x"3aaa",x"400e",x"3775",x"3232",x"ad32",x"3bd2",x"3587",x"34f5",x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2"),
(x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3aae",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3586",x"3512",x"3aaa",x"400e",x"3775",x"3232",x"ad32",x"3bd2",x"3587",x"34f5"),
(x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3aa6",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"358e",x"3523",x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523"),
(x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aac",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3589",x"352f",x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523"),
(x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aaf",x"4025",x"378f",x"317b",x"b4aa",x"3b87",x"3587",x"3537",x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534"),
(x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3ab6",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3581",x"3535",x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534"),
(x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534",x"3ab6",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3581",x"3535"),
(x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534"),
(x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"3ab7",x"400d",x"3776",x"b49f",x"a9d6",x"3ba6",x"357d",x"34f3",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527"),
(x"3ab7",x"400d",x"3776",x"b49f",x"a9d6",x"3ba6",x"357d",x"34f3",x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3aaa",x"400e",x"3775",x"3232",x"ad32",x"3bd2",x"3587",x"34f5",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"3aae",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3586",x"3512",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527"),
(x"3aac",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3589",x"352f",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534",x"3ab6",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3581",x"3535",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534"),
(x"3a9c",x"3fff",x"3770",x"3be8",x"9e0a",x"30d2",x"3648",x"31cd",x"3a9a",x"400d",x"378a",x"3bec",x"2694",x"3049",x"3648",x"317b",x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b"),
(x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f",x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140",x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b"),
(x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b",x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a",x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140"),
(x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102",x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a"),
(x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff",x"3a9c",x"4024",x"37aa",x"3a49",x"b805",x"35c2",x"364a",x"30f4",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"3a95",x"4023",x"37b6",x"39d1",x"b94b",x"31cf",x"3644",x"30fb",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee",x"3a9c",x"4024",x"37aa",x"3a49",x"b805",x"35c2",x"364a",x"30f4"),
(x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a9c",x"4023",x"37c8",x"3b6a",x"b4dc",x"b301",x"363e",x"30f1",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112"),
(x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133"),
(x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a99",x"400d",x"379f",x"3bf8",x"2d3a",x"a850",x"3640",x"3175",x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"3a99",x"400d",x"379f",x"3bf8",x"2d3a",x"a850",x"3640",x"3175",x"3a9b",x"3fff",x"3790",x"3bfe",x"2874",x"9fe2",x"363d",x"31c9",x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174",x"3a9b",x"3fff",x"3790",x"3bfe",x"2874",x"9fe2",x"363d",x"31c9",x"3a9b",x"3fff",x"3798",x"3be2",x"a7a0",x"314d",x"363a",x"31c7"),
(x"3a9a",x"400d",x"37b2",x"3bee",x"a8fd",x"2fea",x"3638",x"3174",x"3a9b",x"4017",x"37d1",x"3bf6",x"a89b",x"2d99",x"3632",x"3134",x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133"),
(x"3a9b",x"4017",x"37d1",x"3bf6",x"a89b",x"2d99",x"3632",x"3134",x"3a9b",x"401d",x"37de",x"3be7",x"9e8d",x"30f1",x"3631",x"3110",x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112"),
(x"3a9b",x"401d",x"37de",x"3be7",x"9e8d",x"30f1",x"3631",x"3110",x"3a9a",x"4022",x"37dc",x"3bdb",x"2a31",x"31d8",x"3635",x"30f7",x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"3a9a",x"4022",x"37dc",x"3bdb",x"2a31",x"31d8",x"3635",x"30f7",x"3a9b",x"4024",x"37cc",x"3bf1",x"2b1d",x"2ec3",x"363d",x"30ea",x"3a9c",x"4023",x"37c8",x"3b6a",x"b4dc",x"b301",x"363e",x"30f1"),
(x"3a9b",x"4024",x"37cc",x"3bf1",x"2b1d",x"2ec3",x"363d",x"30ea",x"3a9c",x"4025",x"37b8",x"3bfc",x"2758",x"2a48",x"3645",x"30e8",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a9c",x"4025",x"37a7",x"3bff",x"21c9",x"251e",x"364c",x"30ed",x"3a9c",x"4024",x"37aa",x"3a49",x"b805",x"35c2",x"364a",x"30f4",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a9c",x"4025",x"37a7",x"3bff",x"21c9",x"251e",x"364c",x"30ed",x"3a9c",x"4022",x"378e",x"3bf3",x"a2c2",x"2edc",x"3654",x"3100",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"3a9c",x"4022",x"378e",x"3bf3",x"a2c2",x"2edc",x"3654",x"3100",x"3a9d",x"4022",x"378b",x"3afb",x"aeb0",x"37a0",x"3656",x"3100",x"3a9d",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"3656",x"311b"),
(x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102",x"3a9c",x"4022",x"378e",x"3bf3",x"a2c2",x"2edc",x"3654",x"3100"),
(x"3a9d",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"3656",x"311b",x"3a9e",x"4017",x"377f",x"3bc6",x"a573",x"337e",x"3654",x"3142",x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140"),
(x"3a9e",x"4017",x"377f",x"3bc6",x"a573",x"337e",x"3654",x"3142",x"3a9d",x"400d",x"3777",x"3bc7",x"a88e",x"3365",x"364f",x"317c",x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b"),
(x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b",x"3a9d",x"400d",x"3777",x"3bc7",x"a88e",x"3365",x"364f",x"317c",x"3a9c",x"3fff",x"3770",x"3be8",x"9e0a",x"30d2",x"3648",x"31cd"),
(x"3a9a",x"400d",x"378a",x"3bec",x"2694",x"3049",x"3648",x"317b",x"3a9c",x"3fff",x"3770",x"3be8",x"9e0a",x"30d2",x"3648",x"31cd",x"3a9b",x"3fff",x"3790",x"3bfe",x"2874",x"9fe2",x"363d",x"31c9"),
(x"3a99",x"400d",x"379f",x"3bf8",x"2d3a",x"a850",x"3640",x"3175",x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f"),
(x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b"),
(x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108"),
(x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff"),
(x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a95",x"4023",x"37b6",x"39d1",x"b94b",x"31cf",x"3644",x"30fb",x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff"),
(x"3a9a",x"400d",x"37b2",x"3866",x"b31b",x"3a70",x"35df",x"33e6",x"3a9b",x"3fff",x"3798",x"3864",x"b1fa",x"3a84",x"35df",x"341e",x"3a7c",x"3ffe",x"37c0",x"a418",x"b372",x"3bc7",x"35c2",x"341c"),
(x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a9b",x"4017",x"37d1",x"386f",x"b4aa",x"3a3c",x"35de",x"33a2"),
(x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a9b",x"401d",x"37de",x"3896",x"af43",x"3a7d",x"35db",x"337c"),
(x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a7b",x"4024",x"37fd",x"a3bb",x"3849",x"3ac0",x"35c1",x"3362",x"3a9a",x"4022",x"37dc",x"3830",x"3619",x"3a17",x"35d9",x"3360"),
(x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351",x"3a9b",x"4024",x"37cc",x"35be",x"3a7e",x"375e",x"35d9",x"334c",x"3a9a",x"4022",x"37dc",x"3830",x"3619",x"3a17",x"35d9",x"3360"),
(x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341",x"3a9c",x"4025",x"37b8",x"3483",x"3bab",x"291b",x"35da",x"333c",x"3a9b",x"4024",x"37cc",x"35be",x"3a7e",x"375e",x"35d9",x"334c"),
(x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331",x"3a9c",x"4025",x"37a7",x"3469",x"3b1b",x"b5df",x"35db",x"332f",x"3a9c",x"4025",x"37b8",x"3483",x"3bab",x"291b",x"35da",x"333c"),
(x"3a93",x"4025",x"379c",x"351a",x"3ab3",x"b716",x"35d5",x"3325",x"3a9c",x"4022",x"378e",x"3718",x"3a24",x"b764",x"35e0",x"3319",x"3a9c",x"4025",x"37a7",x"3469",x"3b1b",x"b5df",x"35db",x"332f"),
(x"3a93",x"4025",x"379c",x"351a",x"3ab3",x"b716",x"35d5",x"3325",x"3a99",x"4023",x"378b",x"38bf",x"3a5d",x"afac",x"35dc",x"3317",x"3a9c",x"4022",x"378e",x"3718",x"3a24",x"b764",x"35e0",x"3319"),
(x"3aa2",x"4023",x"378c",x"b949",x"390d",x"367c",x"3632",x"3477",x"3a9d",x"4022",x"378b",x"b842",x"3832",x"3950",x"3633",x"347b",x"3a9c",x"4022",x"3786",x"b818",x"3947",x"3865",x"3631",x"347c"),
(x"3a9c",x"4022",x"3786",x"36df",x"3aa3",x"35b1",x"35df",x"3313",x"3a9d",x"4022",x"378b",x"380b",x"3a5a",x"3567",x"35e0",x"3316",x"3a9c",x"4022",x"378e",x"3718",x"3a24",x"b764",x"35e0",x"3319"),
(x"3a2a",x"401f",x"3786",x"bae5",x"ae76",x"37f0",x"3652",x"3477",x"3a1a",x"4020",x"3752",x"bacd",x"aeb3",x"381f",x"363b",x"3478",x"3a24",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"363c",x"3466"),
(x"3a31",x"4024",x"378d",x"ba5b",x"36b9",x"3702",x"3655",x"3468",x"3a24",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"363c",x"3466",x"3a2d",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"363e",x"345e"),
(x"3a37",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3656",x"3461",x"3a2d",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"363e",x"345e",x"3a35",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"3640",x"3458"),
(x"3a2a",x"401f",x"3786",x"bae5",x"ae76",x"37f0",x"3652",x"3477",x"3a3b",x"400d",x"3775",x"babf",x"b1e9",x"3808",x"365d",x"34ae",x"3a31",x"400d",x"3752",x"baca",x"b303",x"37b2",x"364e",x"34af"),
(x"3a3b",x"400d",x"3775",x"babf",x"b1e9",x"3808",x"365d",x"34ae",x"3a41",x"4001",x"376d",x"ba5f",x"af27",x"38c0",x"3663",x"34cf",x"3a36",x"4002",x"3752",x"bab1",x"af0f",x"3849",x"3656",x"34ce"),
(x"3a42",x"4027",x"378f",x"2731",x"3bb3",x"3450",x"365a",x"345a",x"3a35",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"3640",x"3458",x"3a4d",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"365e",x"3453"),
(x"3a54",x"4024",x"3782",x"3907",x"3a38",x"a553",x"365e",x"344b",x"3a56",x"4023",x"378c",x"3932",x"391d",x"3695",x"3664",x"344a",x"3a4d",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"365e",x"3453"),
(x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0",x"3a41",x"4001",x"376d",x"b03c",x"aa80",x"3beb",x"3641",x"30bf",x"3a3b",x"400d",x"3775",x"ab97",x"ae90",x"3bf1",x"3642",x"307d"),
(x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079",x"3a3b",x"400d",x"3775",x"ab97",x"ae90",x"3bf1",x"3642",x"307d",x"3a2a",x"401f",x"3786",x"ae5c",x"b067",x"3be2",x"363e",x"300d"),
(x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e",x"3a2a",x"401f",x"3786",x"ae5c",x"b067",x"3be2",x"363e",x"300d",x"3a31",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3645",x"2fe4"),
(x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee",x"3a31",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3645",x"2fe4",x"3a37",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"364b",x"2fd2"),
(x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf",x"3a37",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"364b",x"2fd2",x"3a42",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3653",x"2fce"),
(x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd",x"3a42",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3653",x"2fce",x"3a4d",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"365b",x"2fdd"),
(x"3a4d",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"365b",x"2fdd",x"3a56",x"4023",x"378c",x"287a",x"ad2b",x"3bf8",x"3661",x"3001",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003"),
(x"3a5a",x"4022",x"378b",x"2ef6",x"b0cb",x"3bdc",x"3664",x"3007",x"3a52",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"365c",x"301d",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003"),
(x"3a5b",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3662",x"3020",x"3a5a",x"4017",x"377f",x"27ce",x"aef0",x"3bf2",x"365f",x"3047",x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040"),
(x"3a5a",x"4017",x"377f",x"27ce",x"aef0",x"3bf2",x"365f",x"3047",x"3a5a",x"400d",x"3777",x"a96a",x"ace7",x"3bf8",x"365a",x"3081",x"3a52",x"400e",x"3777",x"ac32",x"ae3d",x"3bf1",x"3654",x"307b"),
(x"3a5a",x"400d",x"3777",x"a96a",x"ace7",x"3bf8",x"365a",x"3081",x"3a5c",x"4000",x"3770",x"ac3e",x"a8a5",x"3bfa",x"3655",x"30cc",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"3a4d",x"400e",x"3775",x"b224",x"ad11",x"3bd3",x"3651",x"3077",x"3a52",x"400e",x"3777",x"ac32",x"ae3d",x"3bf1",x"3654",x"307b",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"3a4d",x"400e",x"3775",x"b224",x"ad11",x"3bd3",x"3651",x"3077",x"3a4a",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3653",x"303e",x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040"),
(x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040",x"3a4a",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3653",x"303e",x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b"),
(x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b",x"3a4c",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3658",x"3004",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003"),
(x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003",x"3a4c",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3658",x"3004",x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5",x"3a42",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd"),
(x"3a42",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf"),
(x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee"),
(x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e"),
(x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079",x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079"),
(x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0",x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079",x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079"),
(x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079",x"3a4d",x"400e",x"3775",x"b224",x"ad11",x"3bd3",x"3651",x"3077",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079",x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a4a",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3653",x"303e"),
(x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b"),
(x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a4c",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3658",x"3004"),
(x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a42",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"3a5e",x"400d",x"378a",x"bbdf",x"2581",x"319c",x"365f",x"2e8f",x"3a5c",x"4000",x"3770",x"bbe7",x"a0ea",x"30f9",x"3661",x"2df3",x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f"),
(x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03",x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03",x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50",x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50",x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f",x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74"),
(x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f",x"3a5c",x"4024",x"37aa",x"ba74",x"b7d3",x"354a",x"3662",x"2f9c",x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89"),
(x"3a5c",x"4024",x"37aa",x"ba74",x"b7d3",x"354a",x"3662",x"2f9c",x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7",x"3a61",x"4023",x"37b7",x"b9e1",x"b96b",x"23fc",x"365c",x"2f93"),
(x"3a61",x"4023",x"37b7",x"b9e1",x"b96b",x"23fc",x"365c",x"2f93",x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"3a61",x"4022",x"37c3",x"baf0",x"b4e6",x"b647",x"3658",x"2f91",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c"),
(x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e",x"3a5d",x"400d",x"37a5",x"bb77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"3a5e",x"3ffd",x"378d",x"bbfd",x"9d53",x"29ab",x"3655",x"2de8",x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a5d",x"400d",x"37a5",x"bb77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"3a5d",x"400d",x"37b0",x"bbfb",x"a724",x"2bb4",x"3651",x"2e9c",x"3a5f",x"3ffd",x"3797",x"bbe2",x"ab03",x"3118",x"3651",x"2de7",x"3a5e",x"3ffd",x"378d",x"bbfd",x"9d53",x"29ab",x"3655",x"2de8"),
(x"3a5d",x"400d",x"37b0",x"bbfb",x"a724",x"2bb4",x"3651",x"2e9c",x"3a5d",x"400d",x"37a5",x"bb77",x"2f4d",x"b571",x"3655",x"2e9c",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"3a5d",x"4017",x"37d0",x"bc00",x"9e59",x"0000",x"364a",x"2f1c",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"3a5c",x"401d",x"37dc",x"bbfd",x"135f",x"a9d9",x"364a",x"2f66",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c"),
(x"3a5d",x"4022",x"37db",x"bbff",x"1b2b",x"2560",x"364e",x"2f95",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"3a5d",x"4024",x"37cd",x"bbf5",x"2bb1",x"2d19",x"3655",x"2fb0",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4",x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7"),
(x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7",x"3a5c",x"4024",x"37aa",x"ba74",x"b7d3",x"354a",x"3662",x"2f9c",x"3a5c",x"4025",x"37a7",x"bbff",x"1fc8",x"2604",x"3664",x"2fa8"),
(x"3a5c",x"4025",x"37a7",x"bbff",x"1fc8",x"2604",x"3664",x"2fa8",x"3a5c",x"4024",x"37aa",x"ba74",x"b7d3",x"354a",x"3662",x"2f9c",x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f"),
(x"3a5a",x"4022",x"378b",x"bafb",x"aeb0",x"37a0",x"366e",x"2f82",x"3a5b",x"4022",x"378e",x"bbf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"3a5b",x"401e",x"3784",x"bbd5",x"a432",x"3275",x"366e",x"2f4e"),
(x"3a5b",x"4022",x"378e",x"bbf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f",x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50"),
(x"3a5b",x"401e",x"3784",x"bbd5",x"a432",x"3275",x"366e",x"2f4e",x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50",x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03"),
(x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"3a5a",x"400d",x"3777",x"bbc5",x"a8bf",x"3387",x"3667",x"2e8b",x"3a5a",x"4017",x"377f",x"bbc6",x"a57a",x"3387",x"366c",x"2f00"),
(x"3a5a",x"400d",x"3777",x"bbc5",x"a8bf",x"3387",x"3667",x"2e8b",x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"3a5c",x"4000",x"3770",x"bbe7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a5e",x"3ffd",x"378d",x"bbfd",x"9d53",x"29ab",x"3655",x"2de8",x"3a5c",x"4000",x"3770",x"bbe7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a5e",x"400d",x"378a",x"bbdf",x"2581",x"319c",x"365f",x"2e8f",x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05",x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e",x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74"),
(x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74",x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89"),
(x"3a61",x"4023",x"37b7",x"b9e1",x"b96b",x"23fc",x"365c",x"2f93",x"3a61",x"4022",x"37c3",x"baf0",x"b4e6",x"b647",x"3658",x"2f91",x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89"),
(x"3a7c",x"3ffe",x"37c0",x"a418",x"b372",x"3bc7",x"35c2",x"341c",x"3a5f",x"3ffd",x"3797",x"b851",x"b1da",x"3a92",x"35a6",x"3422",x"3a5d",x"400d",x"37b0",x"b883",x"b339",x"3a5a",x"35a4",x"33e7"),
(x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a5d",x"400d",x"37b0",x"b883",x"b339",x"3a5a",x"35a4",x"33e7",x"3a5d",x"4017",x"37d0",x"b883",x"b46b",x"3a39",x"35a5",x"33a3"),
(x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a5d",x"4017",x"37d0",x"b883",x"b46b",x"3a39",x"35a5",x"33a3",x"3a5c",x"401d",x"37dc",x"b88e",x"afce",x"3a80",x"35a7",x"337c"),
(x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a5c",x"401d",x"37dc",x"b88e",x"afce",x"3a80",x"35a7",x"337c",x"3a5d",x"4022",x"37db",x"b859",x"3581",x"3a1f",x"35a9",x"3362"),
(x"3a5d",x"4022",x"37db",x"b859",x"3581",x"3a1f",x"35a9",x"3362",x"3a5d",x"4024",x"37cd",x"b609",x"3a62",x"3783",x"35aa",x"334e",x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351"),
(x"3a5d",x"4024",x"37cd",x"b609",x"3a62",x"3783",x"35aa",x"334e",x"3a5c",x"4025",x"37b8",x"b4be",x"3ba1",x"2a04",x"35a8",x"333e",x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341"),
(x"3a5c",x"4025",x"37b8",x"b4be",x"3ba1",x"2a04",x"35a8",x"333e",x"3a5c",x"4025",x"37a7",x"b4f8",x"3b04",x"b5db",x"35a6",x"3332",x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331"),
(x"3a5c",x"4025",x"37a7",x"b4f8",x"3b04",x"b5db",x"35a6",x"3332",x"3a5b",x"4022",x"378e",x"b8e6",x"391d",x"b76f",x"35a1",x"331c",x"3a64",x"4024",x"3789",x"b533",x"3ac8",x"b6b3",x"35a9",x"3318"),
(x"3a5f",x"4023",x"378b",x"b7bc",x"3afd",x"2a6c",x"35a4",x"331a",x"3a64",x"4024",x"3789",x"b533",x"3ac8",x"b6b3",x"35a9",x"3318",x"3a5b",x"4022",x"378e",x"b8e6",x"391d",x"b76f",x"35a1",x"331c"),
(x"3a5d",x"4022",x"3782",x"3856",x"3952",x"381b",x"3662",x"3443",x"3a5a",x"4022",x"378b",x"3889",x"38bf",x"3890",x"3665",x"3446",x"3a56",x"4023",x"378c",x"3932",x"391d",x"3695",x"3664",x"344a"),
(x"3a5f",x"4023",x"378b",x"b7bc",x"3afd",x"2a6c",x"35a4",x"331a",x"3a5b",x"4022",x"378e",x"b8e6",x"391d",x"b76f",x"35a1",x"331c",x"3a5a",x"4022",x"378b",x"b71a",x"3b19",x"2ff1",x"35a0",x"3319"),
(x"3a36",x"4002",x"3752",x"bab1",x"af0f",x"3849",x"3656",x"34ce",x"3a41",x"4001",x"376d",x"ba5f",x"af27",x"38c0",x"3663",x"34cf",x"3a41",x"3ffb",x"376e",x"bab9",x"ac8e",x"384b",x"3665",x"34da"),
(x"3a41",x"4001",x"376d",x"b03c",x"aa80",x"3beb",x"3641",x"30bf",x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0",x"3a4a",x"3fff",x"3770",x"ad3d",x"28c9",x"3bf7",x"3647",x"30ce"),
(x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2",x"3a4a",x"3fff",x"3770",x"ad3d",x"28c9",x"3bf7",x"3647",x"30ce",x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0"),
(x"3a4a",x"3fff",x"3770",x"ad3d",x"28c9",x"3bf7",x"3647",x"30ce",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2",x"3a5c",x"4000",x"3770",x"ac3e",x"a8a5",x"3bfa",x"3655",x"30cc"),
(x"3ab5",x"3ff8",x"376e",x"3afe",x"ac6c",x"37b0",x"3633",x"33c7",x"3ab7",x"4002",x"376d",x"3af0",x"b0d8",x"3796",x"362f",x"33e9",x"3abf",x"4002",x"3752",x"3b07",x"b070",x"374f",x"3623",x"33e8"),
(x"3ab7",x"4002",x"376d",x"2fac",x"ad49",x"3bea",x"357c",x"34d1",x"3ab5",x"3ff8",x"376e",x"2d21",x"068d",x"3bf9",x"357c",x"34c0",x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"3ab5",x"3ff8",x"376e",x"2d23",x"068d",x"3bf9",x"357c",x"34c0",x"3aa4",x"3ffc",x"3770",x"2938",x"1d6d",x"3bfe",x"3589",x"34c5"),
(x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3aa4",x"3ffc",x"3770",x"2938",x"1d6d",x"3bfe",x"3589",x"34c5",x"3a9c",x"3fff",x"3770",x"2e76",x"a942",x"3bf3",x"3590",x"34c9"),
(x"3acd",x"404b",x"3786",x"3af5",x"afa5",x"37a8",x"3610",x"34de",x"3ac7",x"404f",x"378d",x"3a12",x"37f9",x"36b2",x"3613",x"34eb",x"3ad3",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35fb",x"34ec"),
(x"3ac7",x"404f",x"378d",x"3a12",x"37f9",x"36b2",x"3613",x"34eb",x"3ac1",x"4051",x"378e",x"3609",x"3ae2",x"3579",x"3615",x"34f1",x"3acb",x"4053",x"3752",x"3846",x"3a11",x"35f5",x"35fd",x"34f4"),
(x"3ac1",x"4051",x"378e",x"3609",x"3ae2",x"3579",x"3615",x"34f1",x"3ab6",x"4051",x"378f",x"a5dc",x"3bcd",x"330b",x"3619",x"34f8",x"3ac3",x"4053",x"3752",x"af98",x"3bdd",x"3078",x"35ff",x"34f9"),
(x"3ac7",x"403d",x"3752",x"3ad1",x"b46a",x"371a",x"360a",x"34b0",x"3abe",x"403d",x"3777",x"3af8",x"b403",x"36bf",x"3619",x"34b3",x"3acd",x"404b",x"3786",x"3af5",x"afa5",x"37a8",x"3610",x"34de"),
(x"3abf",x"4034",x"3752",x"3afe",x"b17b",x"3746",x"3612",x"3497",x"3ab7",x"4034",x"376d",x"3ae5",x"b1fa",x"378a",x"361e",x"3499",x"3abe",x"403d",x"3777",x"3af8",x"b403",x"36bf",x"3619",x"34b3"),
(x"3ac3",x"4053",x"3752",x"af98",x"3bdd",x"3078",x"35ff",x"34f9",x"3ab6",x"4051",x"378f",x"a5dc",x"3bcd",x"330b",x"3619",x"34f8",x"3aab",x"4051",x"378e",x"b6eb",x"3b36",x"1c18",x"361c",x"34ff"),
(x"3aab",x"4051",x"378e",x"b6eb",x"3b36",x"1c18",x"361c",x"34ff",x"3aa2",x"404e",x"378c",x"b8cb",x"39b0",x"35e1",x"3620",x"3508",x"3aa4",x"404f",x"3782",x"b85b",x"3ab4",x"a80e",x"361b",x"3507"),
(x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3abe",x"403d",x"3777",x"a53f",x"b05f",x"3bec",x"3611",x"3305",x"3ab7",x"4034",x"376d",x"25e3",x"adbf",x"3bf7",x"360e",x"333a"),
(x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3acd",x"404b",x"3786",x"30f8",x"b10a",x"3bcd",x"3619",x"32ae",x"3abe",x"403d",x"3777",x"a53f",x"b05f",x"3bec",x"3611",x"3305"),
(x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3ac7",x"404f",x"378d",x"2f46",x"b040",x"3be0",x"3613",x"3297"),
(x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3ac1",x"4051",x"378e",x"2d5b",x"a17a",x"3bf8",x"360e",x"328f"),
(x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3ab4",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3605",x"3292",x"3ab6",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3aab",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"35fe",x"3292",x"3ab6",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aa2",x"404e",x"378c",x"a877",x"ae68",x"3bf4",x"35f7",x"32a1",x"3aab",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"35fe",x"3292"),
(x"3a9d",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"35f4",x"32a5",x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aa6",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"35fb",x"32b8"),
(x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3a9e",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"35f6",x"32d9",x"3a9d",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"3aa6",x"403d",x"3777",x"2c2a",x"afe7",x"3beb",x"35fe",x"3305",x"3a9d",x"403d",x"3777",x"2bbb",x"ae16",x"3bf2",x"35f8",x"3309",x"3a9e",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"35f6",x"32d9"),
(x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b",x"3a9c",x"4032",x"3770",x"2e75",x"aa83",x"3bf2",x"35fa",x"334a",x"3a9d",x"403d",x"3777",x"2bbb",x"ae16",x"3bf2",x"35f8",x"3309"),
(x"3aa6",x"403d",x"3777",x"2c2a",x"afe7",x"3beb",x"35fe",x"3305",x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302",x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b"),
(x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3aae",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3602",x"32d4",x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3aa6",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4",x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3ab2",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3603",x"329c",x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4"),
(x"3ab4",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3605",x"3292",x"3ab6",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3606",x"329a",x"3ab2",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3603",x"329c"),
(x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b",x"3ab6",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3606",x"329a"),
(x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b"),
(x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1"),
(x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3ab4",x"403d",x"3773",x"adb8",x"ad34",x"3bf1",x"3609",x"3304",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3ab4",x"403d",x"3773",x"adb8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b",x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"3aae",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3602",x"32d4",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0",x"3ab4",x"403d",x"3773",x"adb8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1"),
(x"3ab2",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3603",x"329c",x"3ab6",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3606",x"329a",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b"),
(x"3a9c",x"4032",x"3770",x"3bc5",x"a836",x"338d",x"35a6",x"34c4",x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a9c",x"403d",x"3783",x"3b8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a97",x"4045",x"3794",x"3bbc",x"287e",x"3408",x"35a6",x"348a",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c",x"3a9c",x"404a",x"3790",x"3b17",x"ade0",x"3741",x"35ac",x"347b",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c",x"3a95",x"404d",x"37a3",x"3bd3",x"a9fd",x"3273",x"35a4",x"3474",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470",x"3a9c",x"404f",x"37aa",x"39e5",x"b8ae",x"3566",x"35a5",x"346b",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a95",x"404e",x"37b6",x"393b",x"b9e8",x"313a",x"359f",x"346f",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468",x"3a9c",x"404f",x"37aa",x"39e5",x"b8ae",x"3566",x"35a5",x"346b"),
(x"3a95",x"404e",x"37c1",x"3a55",x"b865",x"b441",x"359c",x"346e",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468"),
(x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477"),
(x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485"),
(x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a99",x"403d",x"379f",x"3bf7",x"2d6b",x"a836",x"359d",x"34a0",x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f"),
(x"3a99",x"403d",x"379f",x"3bf7",x"2d6b",x"a836",x"359d",x"34a0",x"3a99",x"4031",x"378d",x"3bfd",x"1418",x"2a73",x"359b",x"34c3",x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f"),
(x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f",x"3a99",x"4031",x"378d",x"3bfd",x"1418",x"2a73",x"359b",x"34c3",x"3a99",x"4031",x"3795",x"3be2",x"acf4",x"30cb",x"3598",x"34c3"),
(x"3a9a",x"403d",x"37b2",x"3bec",x"ac1f",x"2fcd",x"3595",x"349f",x"3a9b",x"4045",x"37d1",x"3bf6",x"a9b5",x"2d99",x"358e",x"3485",x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485"),
(x"3a9b",x"4045",x"37d1",x"3bf6",x"a9b5",x"2d99",x"358e",x"3485",x"3a9b",x"404a",x"37de",x"3be7",x"a00b",x"30f0",x"358d",x"3476",x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477"),
(x"3a9b",x"404a",x"37de",x"3be7",x"a00b",x"30f0",x"358d",x"3476",x"3a9a",x"404d",x"37dc",x"3bd6",x"2b52",x"322d",x"3590",x"346c",x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"3a9b",x"4050",x"37cc",x"3be3",x"2d8f",x"3091",x"3598",x"3466",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469",x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"3a9c",x"4050",x"37b8",x"3bf8",x"2c16",x"2b31",x"35a1",x"3466",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"3a9c",x"4050",x"37a7",x"3bff",x"232b",x"2518",x"35a7",x"3469",x"3a9c",x"404f",x"37aa",x"39e5",x"b8ae",x"3566",x"35a5",x"346b",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468"),
(x"3a9c",x"4050",x"37a7",x"3bff",x"232b",x"2518",x"35a7",x"3469",x"3a9c",x"404e",x"378e",x"3bf3",x"a432",x"2ede",x"35af",x"3471",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a9c",x"404e",x"378e",x"3bf3",x"a432",x"2ede",x"35af",x"3471",x"3a9d",x"404e",x"378b",x"3af6",x"b023",x"379a",x"35b1",x"3471",x"3a9d",x"404a",x"3784",x"3bd5",x"a532",x"3275",x"35b1",x"347c"),
(x"3a9c",x"404a",x"3790",x"3b17",x"ade0",x"3741",x"35ac",x"347b",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472",x"3a9c",x"404e",x"378e",x"3bf3",x"a432",x"2ede",x"35af",x"3471"),
(x"3a9d",x"404a",x"3784",x"3bd5",x"a532",x"3275",x"35b1",x"347c",x"3a9e",x"4045",x"377f",x"3bc6",x"a6c8",x"337e",x"35b0",x"348c",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a9e",x"4045",x"377f",x"3bc6",x"a6c8",x"337e",x"35b0",x"348c",x"3a9d",x"403d",x"3777",x"3bc6",x"a9a5",x"3364",x"35ac",x"34a4",x"3a9c",x"403d",x"3783",x"3b8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"3a9c",x"403d",x"3783",x"3b8f",x"ab5c",x"3527",x"35a7",x"34a3",x"3a9d",x"403d",x"3777",x"3bc6",x"a9a5",x"3364",x"35ac",x"34a4",x"3a9c",x"4032",x"3770",x"3bc5",x"a836",x"338d",x"35a6",x"34c4"),
(x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a9c",x"4032",x"3770",x"3bc5",x"a836",x"338d",x"35a6",x"34c4",x"3a99",x"4031",x"378d",x"3bfd",x"1418",x"2a73",x"359b",x"34c3"),
(x"3a99",x"403d",x"379f",x"3bf7",x"2d6b",x"a836",x"359d",x"34a0",x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a97",x"4045",x"3794",x"3bbc",x"287e",x"3408",x"35a6",x"348a"),
(x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c"),
(x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a95",x"404d",x"37a3",x"3bd3",x"a9fd",x"3273",x"35a4",x"3474"),
(x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a95",x"404e",x"37c1",x"3a55",x"b865",x"b441",x"359c",x"346e",x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470"),
(x"3a95",x"404e",x"37c1",x"3a55",x"b865",x"b441",x"359c",x"346e",x"3a95",x"404e",x"37b6",x"393b",x"b9e8",x"313a",x"359f",x"346f",x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470"),
(x"3a9a",x"403d",x"37b2",x"386e",x"b47a",x"3a45",x"367a",x"29b1",x"3a99",x"4031",x"3795",x"389a",x"b412",x"3a37",x"3679",x"2ae7",x"3a7c",x"4031",x"37c0",x"9bc8",x"b48d",x"3bab",x"365d",x"2ab9"),
(x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a9b",x"4045",x"37d1",x"3856",x"b5aa",x"3a18",x"3678",x"28cc"),
(x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a9b",x"404a",x"37de",x"3892",x"b07e",x"3a77",x"3675",x"284f"),
(x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a7b",x"4050",x"37fd",x"a32b",x"38f3",x"3a48",x"365b",x"2806",x"3a9a",x"404d",x"37dc",x"3809",x"374a",x"39de",x"3673",x"27ef"),
(x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e",x"3a9b",x"4050",x"37cc",x"34ee",x"3aeb",x"3653",x"3673",x"275d",x"3a9a",x"404d",x"37dc",x"3809",x"374a",x"39de",x"3673",x"27ef"),
(x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709",x"3a9c",x"4050",x"37b8",x"3361",x"3bc7",x"282c",x"3674",x"26df",x"3a9b",x"4050",x"37cc",x"34ee",x"3aeb",x"3653",x"3673",x"275d"),
(x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c",x"3a9c",x"4050",x"37a7",x"3362",x"3b62",x"b4ea",x"3676",x"2679",x"3a9c",x"4050",x"37b8",x"3361",x"3bc7",x"282c",x"3674",x"26df"),
(x"3a93",x"4050",x"379c",x"3458",x"3b15",x"b609",x"366f",x"2623",x"3a9c",x"404e",x"378e",x"362d",x"3aa4",x"b66f",x"3679",x"25cc",x"3a9c",x"4050",x"37a7",x"3362",x"3b62",x"b4ea",x"3676",x"2679"),
(x"3a93",x"4050",x"379c",x"3458",x"3b15",x"b609",x"366f",x"2623",x"3a99",x"404e",x"378b",x"3818",x"3ad2",x"ae9f",x"3676",x"25ba",x"3a9c",x"404e",x"378e",x"362d",x"3aa4",x"b66f",x"3679",x"25cc"),
(x"3aa2",x"404e",x"378c",x"b8cb",x"39b0",x"35e0",x"3620",x"3508",x"3a9d",x"404e",x"378b",x"b7f3",x"38dc",x"38f4",x"3622",x"350b",x"3a9c",x"404e",x"3786",x"b75f",x"39e5",x"37e8",x"3620",x"350c"),
(x"3a9c",x"404e",x"3786",x"35de",x"3b08",x"34dc",x"3679",x"2599",x"3a9d",x"404e",x"378b",x"36fc",x"3ace",x"34ab",x"367a",x"25b5",x"3a9c",x"404e",x"378e",x"362d",x"3aa4",x"b66f",x"3679",x"25cc"),
(x"3a2a",x"404b",x"3786",x"bae1",x"b000",x"37eb",x"35f5",x"2dd3",x"3a1a",x"404c",x"3752",x"bac8",x"b025",x"381c",x"35de",x"2dda",x"3a24",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35e0",x"2d9e"),
(x"3a31",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"35f8",x"2da1",x"3a24",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35e0",x"2d9e",x"3a2d",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35e2",x"2d7f"),
(x"3a37",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"35fa",x"2d8a",x"3a2d",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35e2",x"2d7f",x"3a35",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35e4",x"2d68"),
(x"3a2a",x"404b",x"3786",x"bae1",x"b000",x"37eb",x"35f5",x"2dd3",x"3a3b",x"403c",x"3775",x"bab0",x"b345",x"37fd",x"35ff",x"2e87",x"3a31",x"403d",x"3752",x"bab4",x"b44c",x"3799",x"35f0",x"2e8e"),
(x"3a3b",x"403c",x"3775",x"bab0",x"b345",x"37fd",x"35ff",x"2e87",x"3a41",x"4033",x"376d",x"ba5a",x"b06c",x"38bc",x"3604",x"2ef0",x"3a36",x"4034",x"3752",x"baac",x"b05e",x"3846",x"35f7",x"2ef0"),
(x"3a42",x"4051",x"378f",x"25dc",x"3bcd",x"330b",x"35fe",x"2d6c",x"3a35",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35e4",x"2d68",x"3a4d",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"3601",x"2d50"),
(x"3a54",x"404f",x"3782",x"385d",x"3ab3",x"a49b",x"3600",x"2d31",x"3a56",x"404e",x"378c",x"38b4",x"39be",x"35f4",x"3605",x"2d2d",x"3a4d",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"3601",x"2d50"),
(x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a41",x"4033",x"376d",x"b03b",x"ac08",x"3be9",x"3668",x"2c64",x"3a3b",x"403c",x"3775",x"adad",x"b0c1",x"3be1",x"3667",x"2cd0"),
(x"3a3b",x"403c",x"3775",x"adad",x"b0c1",x"3be1",x"3667",x"2cd0",x"3a2a",x"404b",x"3786",x"b0f0",x"b193",x"3bc7",x"366a",x"2d86",x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83",x"3a2a",x"404b",x"3786",x"b0f0",x"b193",x"3bc7",x"366a",x"2d86",x"3a31",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3663",x"2db2"),
(x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8",x"3a31",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3663",x"2db2",x"3a37",x"4051",x"378e",x"ad5b",x"a17a",x"3bf8",x"365d",x"2dbf"),
(x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4",x"3a37",x"4051",x"378e",x"ad5b",x"a17a",x"3bf8",x"365d",x"2dbf",x"3a42",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3655",x"2dc0"),
(x"3a42",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3655",x"2dc0",x"3a4d",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"364d",x"2db2",x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"3a4d",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"364d",x"2db2",x"3a56",x"404e",x"378c",x"2877",x"ae68",x"3bf4",x"3647",x"2d91",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"3a5a",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"3645",x"2d87",x"3a52",x"404a",x"3788",x"ac6d",x"b1f6",x"3bd7",x"364c",x"2d65",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"3a5b",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"3a5a",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"364a",x"2d20",x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"3a5a",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"364a",x"2d20",x"3a5a",x"403d",x"3777",x"aa04",x"ae02",x"3bf4",x"364f",x"2cc3",x"3a52",x"403d",x"3777",x"ac2f",x"afb9",x"3bec",x"3655",x"2cce"),
(x"3a5a",x"403d",x"3777",x"aa04",x"ae02",x"3bf4",x"364f",x"2cc3",x"3a5c",x"4032",x"3770",x"aca2",x"a97a",x"3bf8",x"3655",x"2c46",x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"3a52",x"403d",x"3777",x"ac2f",x"afb9",x"3bec",x"3655",x"2cce",x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"3a4a",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3656",x"2d31",x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c",x"3a4a",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3656",x"2d31",x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68"),
(x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68",x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d",x"3a46",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3654",x"2d9f",x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"3a46",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3654",x"2d9f",x"3a42",x"4050",x"3787",x"270a",x"b98f",x"39bf",x"3656",x"2da5",x"3a43",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3654",x"2db4"),
(x"3a42",x"4050",x"3787",x"270a",x"b98f",x"39bf",x"3656",x"2da5",x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4"),
(x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8"),
(x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a44",x"403d",x"3773",x"2dae",x"ad20",x"3bf1",x"3660",x"2cd4",x"3a41",x"403d",x"3776",x"331d",x"aca2",x"3bc7",x"3662",x"2cd4"),
(x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a41",x"403d",x"3776",x"331d",x"aca2",x"3bc7",x"3662",x"2cd4",x"3a44",x"403d",x"3773",x"2dae",x"ad20",x"3bf1",x"3660",x"2cd4"),
(x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a44",x"403d",x"3773",x"2dae",x"ad20",x"3bf1",x"3660",x"2cd4",x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5"),
(x"3a44",x"403d",x"3773",x"2dae",x"ad20",x"3bf1",x"3660",x"2cd4",x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a4a",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3656",x"2d31"),
(x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68"),
(x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d"),
(x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a42",x"4050",x"3787",x"270a",x"b98f",x"39bf",x"3656",x"2da5",x"3a46",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3654",x"2d9f"),
(x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8",x"3a5c",x"4032",x"3770",x"bbe2",x"a025",x"3161",x"35f6",x"340d",x"3a5c",x"403d",x"3782",x"bb88",x"abb1",x"354b",x"35f4",x"33d9"),
(x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8",x"3a5c",x"403d",x"3782",x"bb88",x"abb1",x"354b",x"35f4",x"33d9",x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa",x"3a5c",x"404a",x"3790",x"bb10",x"ad8c",x"3760",x"35ed",x"338b",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b"),
(x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b",x"3a5c",x"404a",x"3790",x"bb10",x"ad8c",x"3760",x"35ed",x"338b",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377",x"3a5c",x"404f",x"37aa",x"ba13",x"b891",x"34fa",x"35f4",x"336a",x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"3a5c",x"404f",x"37aa",x"ba13",x"b891",x"34fa",x"35f4",x"336a",x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a61",x"404f",x"37b7",x"b977",x"b9c7",x"2ebe",x"35fa",x"336e"),
(x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a5c",x"404f",x"37c9",x"bb31",x"b5e3",x"b398",x"3600",x"3366",x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e"),
(x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e",x"3a5c",x"404f",x"37c9",x"bb31",x"b5e3",x"b398",x"3600",x"3366",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b"),
(x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b",x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1"),
(x"3a5c",x"4030",x"378d",x"bbfe",x"28c2",x"2138",x"3602",x"340f",x"3a5f",x"403d",x"37a1",x"bbf5",x"2dc9",x"aa2e",x"3600",x"33d2",x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1"),
(x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1",x"3a5d",x"403d",x"37b0",x"bbff",x"a3ef",x"2511",x"3606",x"33d1",x"3a5d",x"4030",x"3797",x"bbf6",x"a3bb",x"2e0a",x"3606",x"340f"),
(x"3a5d",x"403d",x"37b0",x"bbff",x"a3ef",x"2511",x"3606",x"33d1",x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b"),
(x"3a5d",x"4045",x"37d0",x"bc00",x"9fe2",x"8000",x"360b",x"339c",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"3a5c",x"404a",x"37dc",x"bbfd",x"14ea",x"a9d6",x"360c",x"337d",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f",x"3a5c",x"404f",x"37c9",x"bb31",x"b5e3",x"b398",x"3600",x"3366",x"3a5d",x"4050",x"37cd",x"bbfa",x"2874",x"2c13",x"3601",x"3360"),
(x"3a5c",x"404f",x"37c9",x"bb31",x"b5e3",x"b398",x"3600",x"3366",x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a5c",x"4050",x"37b8",x"bbfa",x"2a69",x"2a66",x"35f8",x"3360"),
(x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a5c",x"404f",x"37aa",x"ba13",x"b891",x"34fa",x"35f4",x"336a",x"3a5c",x"4050",x"37a7",x"bbff",x"20dd",x"2604",x"35f2",x"3366"),
(x"3a5c",x"4050",x"37a7",x"bbff",x"20dd",x"2604",x"35f2",x"3366",x"3a5c",x"404f",x"37aa",x"ba13",x"b891",x"34fa",x"35f4",x"336a",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"3a5a",x"404e",x"378b",x"baf6",x"b023",x"379a",x"35e8",x"3377",x"3a5b",x"404e",x"378e",x"bbf3",x"a432",x"2f1d",x"35ea",x"3376",x"3a5b",x"404a",x"3784",x"bbd5",x"a532",x"3275",x"35e9",x"338d"),
(x"3a5b",x"404e",x"378e",x"bbf3",x"a432",x"2f1d",x"35ea",x"3376",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377",x"3a5c",x"404a",x"3790",x"bb10",x"ad8c",x"3760",x"35ed",x"338b"),
(x"3a5b",x"404a",x"3784",x"bbd5",x"a532",x"3275",x"35e9",x"338d",x"3a5c",x"404a",x"3790",x"bb10",x"ad8c",x"3760",x"35ed",x"338b",x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"3a5c",x"403d",x"3782",x"bb88",x"abb1",x"354b",x"35f4",x"33d9",x"3a5a",x"403d",x"3777",x"bbc4",x"a9cf",x"3386",x"35ef",x"33db",x"3a5a",x"4045",x"377f",x"bbc5",x"a6cf",x"3387",x"35eb",x"33ac"),
(x"3a5a",x"403d",x"3777",x"bbc4",x"a9cf",x"3386",x"35ef",x"33db",x"3a5c",x"403d",x"3782",x"bb88",x"abb1",x"354b",x"35f4",x"33d9",x"3a5c",x"4032",x"3770",x"bbe2",x"a025",x"3161",x"35f6",x"340d"),
(x"3a5c",x"4030",x"378d",x"bbfe",x"28c2",x"2138",x"3602",x"340f",x"3a5c",x"4032",x"3770",x"bbe2",x"a025",x"3161",x"35f6",x"340d",x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8"),
(x"3a5f",x"403d",x"37a1",x"bbf5",x"2dc9",x"aa2e",x"3600",x"33d2",x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8",x"3a61",x"4045",x"3794",x"bbd9",x"292f",x"3209",x"35f5",x"33a8"),
(x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a61",x"4045",x"3794",x"bbd9",x"292f",x"3209",x"35f5",x"33a8",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b"),
(x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b",x"3a62",x"404d",x"37a3",x"bbda",x"aea9",x"311c",x"35f5",x"337c"),
(x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a62",x"404d",x"37a3",x"bbda",x"aea9",x"311c",x"35f5",x"337c",x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"3a61",x"404f",x"37b7",x"b977",x"b9c7",x"2ebe",x"35fa",x"336e",x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e",x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"3a7c",x"4031",x"37c0",x"9bc8",x"b48d",x"3bab",x"365d",x"2ab9",x"3a5d",x"4030",x"3797",x"b813",x"b281",x"3ab0",x"3640",x"2b01",x"3a5d",x"403d",x"37b0",x"b860",x"b445",x"3a59",x"363e",x"29b6"),
(x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a5d",x"403d",x"37b0",x"b860",x"b445",x"3a59",x"363e",x"29b6",x"3a5d",x"4045",x"37d0",x"b86c",x"b560",x"3a19",x"3640",x"28d0"),
(x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a5d",x"4045",x"37d0",x"b86c",x"b560",x"3a19",x"3640",x"28d0",x"3a5c",x"404a",x"37dc",x"b889",x"b0d3",x"3a7a",x"3643",x"2852"),
(x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a5c",x"404a",x"37dc",x"b889",x"b0d3",x"3a7a",x"3643",x"2852",x"3a5d",x"404d",x"37db",x"b837",x"36a0",x"39ef",x"3644",x"2800"),
(x"3a5d",x"404d",x"37db",x"b837",x"36a0",x"39ef",x"3644",x"2800",x"3a5d",x"4050",x"37cd",x"b534",x"3ad5",x"367a",x"3644",x"2773",x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e"),
(x"3a5d",x"4050",x"37cd",x"b534",x"3ad5",x"367a",x"3644",x"2773",x"3a5c",x"4050",x"37b8",x"b3c4",x"3bc1",x"28ed",x"3642",x"26f2",x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709"),
(x"3a5c",x"4050",x"37b8",x"b3c4",x"3bc1",x"28ed",x"3642",x"26f2",x"3a5c",x"4050",x"37a7",x"b42d",x"3b51",x"b4ec",x"3641",x"268d",x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c"),
(x"3a5c",x"4050",x"37a7",x"b42d",x"3b51",x"b4ec",x"3641",x"268d",x"3a5b",x"404e",x"378e",x"b86f",x"39bf",x"b6ba",x"363c",x"25e5",x"3a64",x"404f",x"3789",x"b469",x"3b25",x"b5af",x"3644",x"25c3"),
(x"3a5f",x"404e",x"378b",x"b682",x"3b4c",x"297d",x"363f",x"25d0",x"3a64",x"404f",x"3789",x"b469",x"3b25",x"b5af",x"3644",x"25c3",x"3a5b",x"404e",x"378e",x"b86f",x"39bf",x"b6ba",x"363c",x"25e5"),
(x"3a5d",x"404e",x"3782",x"37ca",x"39ef",x"375f",x"3603",x"2d14",x"3a5a",x"404e",x"378b",x"3828",x"3967",x"382f",x"3606",x"2d1e",x"3a56",x"404e",x"378c",x"38b4",x"39be",x"35f4",x"3605",x"2d2d"),
(x"3a5f",x"404e",x"378b",x"b682",x"3b4c",x"297d",x"363f",x"25d0",x"3a5b",x"404e",x"378e",x"b86f",x"39bf",x"b6ba",x"363c",x"25e5",x"3a5a",x"404e",x"378b",x"b5f3",x"3b61",x"2ea6",x"363c",x"25cf"),
(x"3a36",x"4034",x"3752",x"baac",x"b05e",x"3846",x"35f7",x"2ef0",x"3a41",x"4033",x"376d",x"ba5a",x"b06c",x"38bc",x"3604",x"2ef0",x"3a41",x"4030",x"376e",x"bab7",x"ada6",x"384a",x"3606",x"2f15"),
(x"3a41",x"4033",x"376d",x"b03b",x"ac08",x"3be9",x"3668",x"2c64",x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a4a",x"4032",x"3770",x"acfa",x"29bc",x"3bf7",x"3663",x"2c4b"),
(x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c",x"3a4a",x"4032",x"3770",x"acfa",x"29bc",x"3bf7",x"3663",x"2c4b",x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62"),
(x"3a4a",x"4032",x"3770",x"acfa",x"29bc",x"3bf7",x"3663",x"2c4b",x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c",x"3a5c",x"4032",x"3770",x"aca2",x"a97a",x"3bf8",x"3655",x"2c46"),
(x"3ab5",x"402f",x"376e",x"3afb",x"ad7c",x"37ae",x"3622",x"348b",x"3ab7",x"4034",x"376d",x"3ae5",x"b1fa",x"378a",x"361e",x"3499",x"3abf",x"4034",x"3752",x"3afe",x"b17b",x"3746",x"3612",x"3497"),
(x"3ab7",x"4034",x"376d",x"25e3",x"adbf",x"3bf7",x"360e",x"333a",x"3ab5",x"402f",x"376e",x"2d21",x"068d",x"3bf9",x"360e",x"3357",x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a"),
(x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3ab5",x"402f",x"376e",x"2d21",x"068d",x"3bf9",x"360e",x"3357",x"3aa4",x"4031",x"3770",x"2935",x"1ec2",x"3bfe",x"3601",x"3350"),
(x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b",x"3aa4",x"4031",x"3770",x"2935",x"1ec2",x"3bfe",x"3601",x"3350",x"3a9c",x"4032",x"3770",x"2e75",x"aa83",x"3bf2",x"35fa",x"334a"),
(x"3a50",x"405c",x"3752",x"b9fd",x"0000",x"394d",x"35ef",x"2cfe",x"3a50",x"4072",x"3752",x"b9fd",x"0000",x"394d",x"35ef",x"2c07",x"3a80",x"405c",x"37be",x"b9fd",x"0000",x"394d",x"3625",x"2d00"),
(x"3ab1",x"4071",x"3752",x"39ee",x"0cea",x"395e",x"360a",x"2df8",x"3ab1",x"405e",x"3752",x"39ee",x"0a8d",x"395e",x"360a",x"2d16",x"3a80",x"4072",x"37be",x"39ee",x"0a8d",x"395e",x"3641",x"2dfd"),
(x"3a80",x"4072",x"37be",x"38a6",x"b8cf",x"3862",x"35c5",x"2b97",x"3a81",x"407a",x"3802",x"3837",x"b940",x"3851",x"35b4",x"2aa4",x"3ab1",x"4071",x"3752",x"3837",x"b940",x"3851",x"35fc",x"2bb2"),
(x"3a80",x"4072",x"37be",x"b8df",x"b892",x"3866",x"354c",x"349f",x"3a50",x"4072",x"3752",x"b854",x"b926",x"3853",x"3516",x"34a2",x"3a81",x"407a",x"3802",x"b854",x"b926",x"3853",x"355f",x"3481"),
(x"3a77",x"3f4b",x"380f",x"3ac7",x"a224",x"383e",x"3455",x"2566",x"3ab7",x"3f49",x"3754",x"3ab7",x"9f2b",x"3858",x"34ae",x"259c",x"3a79",x"3dc3",x"3804",x"3ab6",x"9af6",x"385a",x"345b",x"311f"),
(x"3a3b",x"3dc2",x"3752",x"ba9d",x"90ea",x"3880",x"34b4",x"3123",x"3a3b",x"3f46",x"3755",x"babd",x"9ffc",x"384e",x"34af",x"25db",x"3a79",x"3dc3",x"3804",x"babc",x"9c9b",x"3850",x"3507",x"311e"),
(x"3ab6",x"3dc2",x"3752",x"3873",x"3a03",x"35ad",x"349d",x"3544",x"3ade",x"3db3",x"3752",x"38d1",x"395c",x"36f1",x"348c",x"3524",x"3a79",x"3dc3",x"3804",x"38d1",x"395c",x"36f1",x"34f0",x"3544"),
(x"3a3b",x"3dc2",x"3752",x"b88b",x"39de",x"35f7",x"34e6",x"3520",x"3a79",x"3dc3",x"3804",x"b8d0",x"395f",x"36e9",x"3493",x"3520",x"3a14",x"3db3",x"3752",x"b8d0",x"395f",x"36e9",x"34f7",x"3500"),
(x"3ade",x"3db3",x"3752",x"3a6b",x"19bc",x"38c5",x"3513",x"2bf1",x"3ade",x"3d4c",x"3752",x"3a6d",x"1c32",x"38c3",x"3512",x"263e",x"3a78",x"3db1",x"3832",x"3a6d",x"1bfc",x"38c3",x"358f",x"2bd9"),
(x"3a14",x"3db3",x"3752",x"ba75",x"20ea",x"38b8",x"3507",x"3363",x"3a78",x"3db1",x"3832",x"ba6f",x"1d6d",x"38c0",x"3587",x"3369",x"3a11",x"3d4d",x"3752",x"ba6f",x"1d53",x"38c0",x"3505",x"3446"),
(x"3a11",x"3ca2",x"3752",x"128d",x"b9fe",x"394b",x"34fa",x"3435",x"3a14",x"3cfa",x"3872",x"1bc8",x"b9fb",x"394f",x"34fa",x"34f8",x"3ae0",x"3ca2",x"3752",x"1b93",x"b9fc",x"394f",x"345f",x"3435"),
(x"3a14",x"3397",x"3877",x"1ffc",x"3a32",x"390e",x"34fa",x"3130",x"3a12",x"351b",x"3752",x"8e8d",x"3a2a",x"3918",x"34fa",x"32b2",x"3adf",x"3396",x"3874",x"8e8d",x"3a2a",x"3918",x"3461",x"3131"),
(x"3a14",x"3397",x"3877",x"1dd6",x"ba2a",x"3918",x"34f9",x"3428",x"3adf",x"3396",x"3874",x"168d",x"ba26",x"391d",x"3465",x"3428",x"3a12",x"30ef",x"3752",x"16f6",x"ba26",x"391d",x"34f9",x"32bf"),
(x"3ade",x"4020",x"3752",x"3acd",x"aeb3",x"381f",x"3609",x"344a",x"3acd",x"401f",x"3786",x"3af9",x"ae2b",x"37ad",x"3620",x"344a",x"3ad3",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"360a",x"345b"),
(x"3ad3",x"4026",x"3752",x"3a59",x"35e6",x"37bd",x"360a",x"345b",x"3ac7",x"4024",x"378d",x"3a5b",x"36b9",x"3703",x"3622",x"3459",x"3acb",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"360c",x"3464"),
(x"3acb",x"4028",x"3752",x"38c9",x"3979",x"36ab",x"360c",x"3464",x"3ac1",x"4026",x"378e",x"3704",x"3a72",x"365d",x"3624",x"3460",x"3ac3",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"360e",x"346a"),
(x"3ade",x"4020",x"3752",x"3acd",x"aeb3",x"381f",x"3609",x"344a",x"3ac7",x"400d",x"3752",x"3ae9",x"b336",x"3733",x"361b",x"3412",x"3acd",x"401f",x"3786",x"3af9",x"ae2b",x"37ad",x"3620",x"344a"),
(x"3ac7",x"400d",x"3752",x"3ae9",x"b336",x"3733",x"361b",x"3412",x"3abf",x"4002",x"3752",x"3b07",x"b070",x"374f",x"3623",x"33e8",x"3abe",x"400d",x"3777",x"3b0c",x"b28a",x"36d3",x"362a",x"3414"),
(x"3ac3",x"4029",x"3752",x"b0ac",x"3bcb",x"3180",x"360e",x"346a",x"3aab",x"4026",x"378e",x"b817",x"3adf",x"1c67",x"362c",x"346e",x"3aa4",x"4024",x"3782",x"b904",x"3a39",x"a8ac",x"362c",x"3476"),
(x"3ab7",x"400d",x"3776",x"b49f",x"a9d6",x"3ba6",x"357d",x"34f3",x"3abe",x"400d",x"3777",x"1d6d",x"aedf",x"3bf4",x"3578",x"34f2",x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2"),
(x"3ab7",x"400d",x"3776",x"b49f",x"a9d6",x"3ba6",x"357d",x"34f3",x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3abe",x"400d",x"3777",x"1d6d",x"aedf",x"3bf4",x"3578",x"34f2"),
(x"3acd",x"401f",x"3786",x"30fd",x"b013",x"3bd6",x"356f",x"3528",x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3ac7",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3575",x"3536"),
(x"3ac7",x"4024",x"378d",x"2f4b",x"aede",x"3be6",x"3575",x"3536",x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3ac1",x"4026",x"378e",x"2d5c",x"a074",x"3bf8",x"357a",x"353b"),
(x"3ac1",x"4026",x"378e",x"2d5c",x"a074",x"3bf8",x"357a",x"353b",x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3ab6",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3582",x"353d"),
(x"3ab6",x"4027",x"378f",x"2231",x"2850",x"3bfe",x"3582",x"353d",x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3aab",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"3aaf",x"4025",x"378f",x"317b",x"b4aa",x"3b87",x"3587",x"3537",x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aab",x"4026",x"378e",x"ad20",x"a16d",x"3bf9",x"358a",x"353a"),
(x"3a9d",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3594",x"352f",x"3aa6",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"358e",x"3523",x"3a9d",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"3aa2",x"4023",x"378c",x"a87a",x"ad2b",x"3bf8",x"3591",x"3531",x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3a9d",x"4022",x"378b",x"aef6",x"b0cc",x"3bdc",x"3594",x"352f"),
(x"3aa6",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"358e",x"3523",x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3a9d",x"401e",x"3784",x"af97",x"b08d",x"3bdc",x"3594",x"3522"),
(x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3aa6",x"400e",x"3777",x"2c2d",x"ae61",x"3bf1",x"358b",x"34f3",x"3a9e",x"4017",x"377f",x"a7ce",x"aef0",x"3bf2",x"3593",x"350f"),
(x"3aa6",x"400e",x"3777",x"2c2d",x"ae61",x"3bf1",x"358b",x"34f3",x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3a9d",x"400d",x"3777",x"2bbe",x"acea",x"3bf6",x"3591",x"34f1"),
(x"3aa6",x"400e",x"3777",x"2c2d",x"ae61",x"3bf1",x"358b",x"34f3",x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3aaa",x"400e",x"3775",x"3232",x"ad32",x"3bd2",x"3587",x"34f5"),
(x"3aae",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3586",x"3512",x"3aa8",x"4018",x"3780",x"316d",x"af52",x"3bd4",x"358b",x"3511",x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523"),
(x"3aa6",x"401e",x"3788",x"2c75",x"b0d4",x"3be3",x"358e",x"3523",x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523"),
(x"3aac",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3589",x"352f",x"3aa8",x"4022",x"378c",x"327a",x"b214",x"3baf",x"358c",x"3530",x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534"),
(x"3aaf",x"4025",x"378f",x"317b",x"b4aa",x"3b87",x"3587",x"3537",x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534"),
(x"3ab4",x"4025",x"3790",x"274b",x"b568",x"3b86",x"3583",x"3539",x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3ab6",x"4024",x"3787",x"a7bb",x"b8ea",x"3a4e",x"3581",x"3535"),
(x"3abd",x"4025",x"378f",x"ad99",x"b52b",x"3b89",x"357c",x"3538",x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534"),
(x"3ac2",x"4023",x"378d",x"b3c6",x"b397",x"3b86",x"3578",x"3534",x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"3ac6",x"401f",x"3788",x"b0d4",x"aed9",x"3bdc",x"3574",x"3528",x"3ab7",x"400d",x"3776",x"b49f",x"a9d6",x"3ba6",x"357d",x"34f3",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527"),
(x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"3aaa",x"400e",x"3775",x"3232",x"ad32",x"3bd2",x"3587",x"34f5",x"3aae",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3586",x"3512",x"3ab4",x"400e",x"3773",x"ac3c",x"ac0d",x"3bf7",x"3580",x"34f3"),
(x"3aae",x"4018",x"377a",x"2c36",x"aec3",x"3bf0",x"3586",x"3512",x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523",x"3ac2",x"401f",x"3782",x"b116",x"adfa",x"3bdc",x"3578",x"3527"),
(x"3aaa",x"401e",x"3782",x"315c",x"b078",x"3bce",x"358a",x"3523",x"3aac",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3589",x"352f",x"3abf",x"4023",x"3785",x"ae71",x"b13e",x"3bd9",x"357b",x"3531"),
(x"3aac",x"4022",x"3787",x"30b8",x"b106",x"3bcf",x"3589",x"352f",x"3ab2",x"4024",x"3787",x"34c3",x"b626",x"3afd",x"3585",x"3534",x"3abb",x"4024",x"3787",x"b08d",x"b423",x"3ba4",x"357e",x"3534"),
(x"3a9a",x"400d",x"378a",x"3bec",x"2694",x"3049",x"3648",x"317b",x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f",x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b"),
(x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f",x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b",x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140"),
(x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b",x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108",x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a"),
(x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108",x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff",x"3a95",x"4023",x"37b6",x"39d1",x"b94b",x"31cf",x"3644",x"30fb",x"3a9c",x"4024",x"37aa",x"3a49",x"b805",x"35c2",x"364a",x"30f4"),
(x"3a95",x"4023",x"37b6",x"39d1",x"b94b",x"31cf",x"3644",x"30fb",x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a9c",x"4023",x"37c8",x"3b6a",x"b4dc",x"b301",x"363e",x"30f1",x"3a95",x"4022",x"37c1",x"3a68",x"b74a",x"b638",x"3640",x"30fb",x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb",x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112"),
(x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112",x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133"),
(x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133",x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174"),
(x"3a9a",x"400d",x"37b2",x"3bee",x"a8fd",x"2fea",x"3638",x"3174",x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174",x"3a9b",x"3fff",x"3798",x"3be2",x"a7a0",x"314d",x"363a",x"31c7"),
(x"3a9b",x"400d",x"37a7",x"3bb8",x"2e24",x"b3c9",x"363c",x"3174",x"3a9a",x"400d",x"37b2",x"3bee",x"a8fd",x"2fea",x"3638",x"3174",x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133"),
(x"3a9b",x"4018",x"37c6",x"3b58",x"3009",x"b604",x"3636",x"3133",x"3a9b",x"4017",x"37d1",x"3bf6",x"a89b",x"2d99",x"3632",x"3134",x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112"),
(x"3a9b",x"401d",x"37d4",x"3b44",x"2867",x"b6a9",x"3635",x"3112",x"3a9b",x"401d",x"37de",x"3be7",x"9e8d",x"30f1",x"3631",x"3110",x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb"),
(x"3a9b",x"4021",x"37d2",x"3b5b",x"afb9",x"b5f8",x"3638",x"30fb",x"3a9a",x"4022",x"37dc",x"3bdb",x"2a31",x"31d8",x"3635",x"30f7",x"3a9c",x"4023",x"37c8",x"3b6a",x"b4dc",x"b301",x"363e",x"30f1"),
(x"3a9c",x"4023",x"37c8",x"3b6a",x"b4dc",x"b301",x"363e",x"30f1",x"3a9b",x"4024",x"37cc",x"3bf1",x"2b1d",x"2ec3",x"363d",x"30ea",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a9c",x"4025",x"37b8",x"3bfc",x"2758",x"2a48",x"3645",x"30e8",x"3a9c",x"4025",x"37a7",x"3bff",x"21c9",x"251e",x"364c",x"30ed",x"3a9c",x"4024",x"37b7",x"3b1c",x"b755",x"a280",x"3645",x"30ee"),
(x"3a9c",x"4024",x"37aa",x"3a49",x"b805",x"35c2",x"364a",x"30f4",x"3a9c",x"4025",x"37a7",x"3bff",x"21c9",x"251e",x"364c",x"30ed",x"3a9c",x"4021",x"3799",x"3afb",x"b3ae",x"36ce",x"3650",x"3102"),
(x"3a9d",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"3656",x"311b",x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a",x"3a9c",x"4022",x"378e",x"3bf3",x"a2c2",x"2edc",x"3654",x"3100"),
(x"3a9c",x"401e",x"3790",x"3ad6",x"aec0",x"3811",x"3651",x"311a",x"3a9d",x"401e",x"3784",x"3bd5",x"a432",x"3276",x"3656",x"311b",x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140"),
(x"3a9c",x"4017",x"378b",x"3aba",x"aa69",x"384e",x"364f",x"3140",x"3a9e",x"4017",x"377f",x"3bc6",x"a573",x"337e",x"3654",x"3142",x"3a9c",x"400d",x"3783",x"3b43",x"aa24",x"36a7",x"364a",x"317b"),
(x"3a99",x"400d",x"379f",x"3bf8",x"2d3a",x"a850",x"3640",x"3175",x"3a9a",x"400d",x"378a",x"3bec",x"2694",x"3049",x"3648",x"317b",x"3a9b",x"3fff",x"3790",x"3bfe",x"2874",x"9fe2",x"363d",x"31c9"),
(x"3a9a",x"400d",x"378a",x"3bec",x"2694",x"3049",x"3648",x"317b",x"3a99",x"400d",x"379f",x"3bf8",x"2d3a",x"a850",x"3640",x"3175",x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f"),
(x"3a97",x"4017",x"3794",x"3bb1",x"25b5",x"345f",x"364a",x"313f",x"3a95",x"4018",x"37ba",x"3bde",x"2e0d",x"b0f4",x"363d",x"3133",x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b"),
(x"3a96",x"401d",x"3798",x"3bae",x"a832",x"3470",x"364c",x"311b",x"3a95",x"401d",x"37c9",x"3bcd",x"2c2d",x"b2c6",x"363b",x"3114",x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108"),
(x"3a95",x"4021",x"37a3",x"3bab",x"abf9",x"346d",x"3649",x"3108",x"3a95",x"4021",x"37c7",x"3b8c",x"a849",x"b547",x"363e",x"3102",x"3a95",x"4022",x"37ac",x"3b0b",x"b542",x"3578",x"3647",x"30ff"),
(x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a9a",x"400d",x"37b2",x"3866",x"b31b",x"3a70",x"35df",x"33e6",x"3a7c",x"3ffe",x"37c0",x"a418",x"b372",x"3bc7",x"35c2",x"341c"),
(x"3a9a",x"400d",x"37b2",x"3866",x"b31b",x"3a70",x"35df",x"33e6",x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a9b",x"4017",x"37d1",x"386f",x"b4aa",x"3a3c",x"35de",x"33a2"),
(x"3a9b",x"4017",x"37d1",x"386f",x"b4aa",x"3a3c",x"35de",x"33a2",x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a9b",x"401d",x"37de",x"3896",x"af43",x"3a7d",x"35db",x"337c"),
(x"3a9b",x"401d",x"37de",x"3896",x"af43",x"3a7d",x"35db",x"337c",x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a9a",x"4022",x"37dc",x"3830",x"3619",x"3a17",x"35d9",x"3360"),
(x"3a7b",x"4024",x"37fd",x"a3bb",x"3849",x"3ac0",x"35c1",x"3362",x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351",x"3a9a",x"4022",x"37dc",x"3830",x"3619",x"3a17",x"35d9",x"3360"),
(x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351",x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341",x"3a9b",x"4024",x"37cc",x"35be",x"3a7e",x"375e",x"35d9",x"334c"),
(x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341",x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331",x"3a9c",x"4025",x"37b8",x"3483",x"3bab",x"291b",x"35da",x"333c"),
(x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331",x"3a93",x"4025",x"379c",x"351a",x"3ab3",x"b716",x"35d5",x"3325",x"3a9c",x"4025",x"37a7",x"3469",x"3b1b",x"b5df",x"35db",x"332f"),
(x"3aa4",x"4024",x"3782",x"b904",x"3a39",x"a8ac",x"362c",x"3476",x"3aa2",x"4023",x"378c",x"b949",x"390d",x"367c",x"3632",x"3477",x"3a9c",x"4022",x"3786",x"b818",x"3947",x"3865",x"3631",x"347c"),
(x"3a99",x"4023",x"378b",x"38bf",x"3a5d",x"afac",x"35dc",x"3317",x"3a9c",x"4022",x"3786",x"36df",x"3aa3",x"35b1",x"35df",x"3313",x"3a9c",x"4022",x"378e",x"3718",x"3a24",x"b764",x"35e0",x"3319"),
(x"3a31",x"4024",x"378d",x"ba5b",x"36b9",x"3702",x"3655",x"3468",x"3a2a",x"401f",x"3786",x"bae5",x"ae76",x"37f0",x"3652",x"3477",x"3a24",x"4026",x"3752",x"ba59",x"35e6",x"37bd",x"363c",x"3466"),
(x"3a37",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3656",x"3461",x"3a31",x"4024",x"378d",x"ba5b",x"36b9",x"3702",x"3655",x"3468",x"3a2d",x"4028",x"3752",x"b8c9",x"3979",x"36ab",x"363e",x"345e"),
(x"3a42",x"4027",x"378f",x"2731",x"3bb3",x"3450",x"365a",x"345a",x"3a37",x"4026",x"378e",x"b704",x"3a72",x"365d",x"3656",x"3461",x"3a35",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"3640",x"3458"),
(x"3a1a",x"4020",x"3752",x"bacd",x"aeb3",x"381f",x"363b",x"3478",x"3a2a",x"401f",x"3786",x"bae5",x"ae76",x"37f0",x"3652",x"3477",x"3a31",x"400d",x"3752",x"baca",x"b303",x"37b2",x"364e",x"34af"),
(x"3a31",x"400d",x"3752",x"baca",x"b303",x"37b2",x"364e",x"34af",x"3a3b",x"400d",x"3775",x"babf",x"b1e9",x"3808",x"365d",x"34ae",x"3a36",x"4002",x"3752",x"bab1",x"af0f",x"3849",x"3656",x"34ce"),
(x"3a35",x"4029",x"3752",x"30ac",x"3bcb",x"3180",x"3640",x"3458",x"3a54",x"4024",x"3782",x"3907",x"3a38",x"a553",x"365e",x"344b",x"3a4d",x"4026",x"378e",x"3817",x"3adf",x"1cd0",x"365e",x"3453"),
(x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079",x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0",x"3a3b",x"400d",x"3775",x"ab97",x"ae90",x"3bf1",x"3642",x"307d"),
(x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e",x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079",x"3a2a",x"401f",x"3786",x"ae5c",x"b067",x"3be2",x"363e",x"300d"),
(x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee",x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e",x"3a31",x"4024",x"378d",x"af4b",x"aede",x"3be6",x"3645",x"2fe4"),
(x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf",x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee",x"3a37",x"4026",x"378e",x"ad5c",x"a067",x"3bf8",x"364b",x"2fd2"),
(x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd",x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf",x"3a42",x"4027",x"378f",x"a231",x"2850",x"3bfe",x"3653",x"2fce"),
(x"3a49",x"4025",x"378f",x"b17c",x"b4aa",x"3b87",x"3658",x"2fe7",x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd",x"3a4d",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"365b",x"2fdd"),
(x"3a49",x"4025",x"378f",x"b17c",x"b4aa",x"3b87",x"3658",x"2fe7",x"3a4d",x"4026",x"378e",x"2d20",x"a16d",x"3bf9",x"365b",x"2fdd",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003"),
(x"3a5a",x"4022",x"378b",x"2ef6",x"b0cb",x"3bdc",x"3664",x"3007",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003",x"3a56",x"4023",x"378c",x"287a",x"ad2b",x"3bf8",x"3661",x"3001"),
(x"3a5b",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3662",x"3020",x"3a52",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"365c",x"301d",x"3a5a",x"4022",x"378b",x"2ef6",x"b0cb",x"3bdc",x"3664",x"3007"),
(x"3a52",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"365c",x"301d",x"3a5b",x"401e",x"3784",x"2f97",x"b08d",x"3bdc",x"3662",x"3020",x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040"),
(x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040",x"3a5a",x"4017",x"377f",x"27ce",x"aef0",x"3bf2",x"365f",x"3047",x"3a52",x"400e",x"3777",x"ac32",x"ae3d",x"3bf1",x"3654",x"307b"),
(x"3a52",x"400e",x"3777",x"ac32",x"ae3d",x"3bf1",x"3654",x"307b",x"3a5a",x"400d",x"3777",x"a96a",x"ace7",x"3bf8",x"365a",x"3081",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"3a52",x"400e",x"3777",x"ac32",x"ae3d",x"3bf1",x"3654",x"307b",x"3a4d",x"400e",x"3775",x"b224",x"ad11",x"3bd3",x"3651",x"3077",x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040"),
(x"3a52",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"365c",x"301d",x"3a50",x"4018",x"3780",x"b16d",x"af52",x"3bd4",x"3658",x"3040",x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b"),
(x"3a52",x"401e",x"3788",x"ac75",x"b0d4",x"3be3",x"365c",x"301d",x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003"),
(x"3a49",x"4025",x"378f",x"b17c",x"b4aa",x"3b87",x"3658",x"2fe7",x"3a50",x"4022",x"378c",x"b27a",x"b213",x"3baf",x"365c",x"3003",x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"3a49",x"4025",x"378f",x"b17c",x"b4aa",x"3b87",x"3658",x"2fe7",x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5",x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd"),
(x"3a43",x"4025",x"3790",x"a74b",x"b568",x"3b86",x"3654",x"2fdd",x"3a42",x"4024",x"3787",x"27bb",x"b8ea",x"3a4e",x"3652",x"2fee",x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf"),
(x"3a3b",x"4025",x"378f",x"2d99",x"b52b",x"3b89",x"364d",x"2fdf",x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee"),
(x"3a36",x"4023",x"378d",x"33c6",x"b397",x"3b86",x"3648",x"2fee",x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e"),
(x"3a31",x"401f",x"3788",x"3153",x"afe4",x"3bd3",x"3643",x"300e",x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a41",x"400d",x"3776",x"2ff7",x"ad4e",x"3be9",x"3647",x"3079"),
(x"3a48",x"4001",x"376f",x"a217",x"aa2e",x"3bfd",x"3646",x"30c0",x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079",x"3a54",x"4002",x"3770",x"abef",x"aa2e",x"3bf9",x"364f",x"30c2"),
(x"3a4d",x"400e",x"3775",x"b224",x"ad11",x"3bd3",x"3651",x"3077",x"3a44",x"400e",x"3773",x"2c28",x"abec",x"3bf7",x"3649",x"3079",x"3a4a",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3653",x"303e"),
(x"3a4a",x"4018",x"377a",x"ac36",x"aec3",x"3bf0",x"3653",x"303e",x"3a35",x"401f",x"3782",x"3115",x"adfa",x"3bdc",x"3647",x"3011",x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b"),
(x"3a4e",x"401e",x"3782",x"b15c",x"b078",x"3bce",x"3658",x"301b",x"3a39",x"4023",x"3785",x"2e71",x"b13e",x"3bd9",x"364b",x"2ffc",x"3a4c",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3658",x"3004"),
(x"3a4c",x"4022",x"3787",x"b0b8",x"b106",x"3bcf",x"3658",x"3004",x"3a3d",x"4024",x"3787",x"308d",x"b423",x"3ba4",x"364e",x"2ff0",x"3a46",x"4024",x"3787",x"b4c3",x"b626",x"3afd",x"3655",x"2ff5"),
(x"3a5e",x"400d",x"378a",x"bbdf",x"2581",x"319c",x"365f",x"2e8f",x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05",x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03",x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e",x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50",x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74"),
(x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74",x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f",x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89"),
(x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89",x"3a5c",x"4024",x"37aa",x"ba74",x"b7d3",x"354a",x"3662",x"2f9c",x"3a61",x"4023",x"37b7",x"b9e1",x"b96b",x"23fc",x"365c",x"2f93"),
(x"3a61",x"4022",x"37c3",x"baf0",x"b4e6",x"b647",x"3658",x"2f91",x"3a61",x"4023",x"37b7",x"b9e1",x"b96b",x"23fc",x"365c",x"2f93",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a61",x"4022",x"37c3",x"baf0",x"b4e6",x"b647",x"3658",x"2f91",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c"),
(x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a5d",x"400d",x"37a5",x"bb77",x"2f4d",x"b571",x"3655",x"2e9c"),
(x"3a5d",x"400d",x"37a5",x"bb77",x"2f4d",x"b571",x"3655",x"2e9c",x"3a5d",x"400d",x"37b0",x"bbfb",x"a724",x"2bb4",x"3651",x"2e9c",x"3a5e",x"3ffd",x"378d",x"bbfd",x"9d53",x"29ab",x"3655",x"2de8"),
(x"3a5d",x"4017",x"37d0",x"bc00",x"9e59",x"0000",x"364a",x"2f1c",x"3a5d",x"400d",x"37b0",x"bbfb",x"a724",x"2bb4",x"3651",x"2e9c",x"3a5d",x"4018",x"37c6",x"bb32",x"3043",x"b6a8",x"364e",x"2f1e"),
(x"3a5c",x"401d",x"37dc",x"bbfd",x"135f",x"a9d9",x"364a",x"2f66",x"3a5d",x"4017",x"37d0",x"bc00",x"9e59",x"0000",x"364a",x"2f1c",x"3a5d",x"401d",x"37d2",x"bafe",x"29bc",x"b7b9",x"364e",x"2f61"),
(x"3a5d",x"4022",x"37db",x"bbff",x"1b2b",x"2560",x"364e",x"2f95",x"3a5c",x"401d",x"37dc",x"bbfd",x"135f",x"a9d9",x"364a",x"2f66",x"3a5d",x"4021",x"37d0",x"bb35",x"af71",x"b6b1",x"3651",x"2f8c"),
(x"3a5d",x"4024",x"37cd",x"bbf5",x"2bb1",x"2d19",x"3655",x"2fb0",x"3a5d",x"4022",x"37db",x"bbff",x"1b2b",x"2560",x"364e",x"2f95",x"3a5c",x"4023",x"37c9",x"bb3e",x"b59b",x"b3a1",x"3656",x"2fa4"),
(x"3a5c",x"4025",x"37b8",x"bbfd",x"208e",x"29e9",x"365e",x"2fb3",x"3a5d",x"4024",x"37cd",x"bbf5",x"2bb1",x"2d19",x"3655",x"2fb0",x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7"),
(x"3a5c",x"4025",x"37b8",x"bbfd",x"208e",x"29e9",x"365e",x"2fb3",x"3a5c",x"4024",x"37b7",x"bb7d",x"b59c",x"2594",x"365e",x"2fa7",x"3a5c",x"4025",x"37a7",x"bbff",x"1fc8",x"2604",x"3664",x"2fa8"),
(x"3a5b",x"4022",x"378e",x"bbf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"3a5c",x"4025",x"37a7",x"bbff",x"1fc8",x"2604",x"3664",x"2fa8",x"3a5b",x"4021",x"3798",x"baff",x"b392",x"36c4",x"3668",x"2f7f"),
(x"3a5b",x"401e",x"3784",x"bbd5",x"a432",x"3275",x"366e",x"2f4e",x"3a5b",x"4022",x"378e",x"bbf3",x"a2c2",x"2f1d",x"366c",x"2f83",x"3a5c",x"401e",x"3790",x"bad4",x"ae75",x"3815",x"3669",x"2f50"),
(x"3a5a",x"4017",x"377f",x"bbc6",x"a57a",x"3387",x"366c",x"2f00",x"3a5b",x"401e",x"3784",x"bbd5",x"a432",x"3275",x"366e",x"2f4e",x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03"),
(x"3a5c",x"4017",x"378b",x"baba",x"aab1",x"384d",x"3667",x"2f03",x"3a5c",x"400d",x"3782",x"bb3d",x"aa5f",x"36c0",x"3663",x"2e8f",x"3a5a",x"4017",x"377f",x"bbc6",x"a57a",x"3387",x"366c",x"2f00"),
(x"3a5e",x"400d",x"378a",x"bbdf",x"2581",x"319c",x"365f",x"2e8f",x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a5c",x"4000",x"3770",x"bbe7",x"a0ea",x"30f9",x"3661",x"2df3"),
(x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a5f",x"400d",x"37a1",x"bbfd",x"2a97",x"9553",x"3657",x"2e9c",x"3a61",x"4017",x"3794",x"bbcf",x"2680",x"32e2",x"3662",x"2f05"),
(x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a62",x"4018",x"37be",x"bbe0",x"2e19",x"b0b1",x"3654",x"2f20",x"3a61",x"401d",x"3798",x"bbbc",x"a231",x"3410",x"3664",x"2f4e"),
(x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a63",x"401d",x"37c9",x"bbcf",x"2b2e",x"b2a9",x"3653",x"2f5a",x"3a62",x"4021",x"37a3",x"bbbc",x"ae5c",x"3383",x"3662",x"2f74"),
(x"3a61",x"4022",x"37c3",x"baf0",x"b4e6",x"b647",x"3658",x"2f91",x"3a62",x"4021",x"37c9",x"bb92",x"ad66",x"b4fc",x"3655",x"2f83",x"3a62",x"4022",x"37ac",x"bb40",x"b55d",x"341d",x"3660",x"2f89"),
(x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a7c",x"3ffe",x"37c0",x"a418",x"b372",x"3bc7",x"35c2",x"341c",x"3a5d",x"400d",x"37b0",x"b883",x"b339",x"3a5a",x"35a4",x"33e7"),
(x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a7b",x"400d",x"37dc",x"a1fd",x"b51b",x"3b94",x"35c1",x"33de",x"3a5d",x"4017",x"37d0",x"b883",x"b46b",x"3a39",x"35a5",x"33a3"),
(x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a7d",x"4019",x"3800",x"a2f6",x"b49e",x"3ba8",x"35c2",x"3397",x"3a5c",x"401d",x"37dc",x"b88e",x"afce",x"3a80",x"35a7",x"337c"),
(x"3a7b",x"4024",x"37fd",x"a3bb",x"3849",x"3ac0",x"35c1",x"3362",x"3a7c",x"401f",x"3804",x"a194",x"2a70",x"3bfd",x"35c2",x"3379",x"3a5d",x"4022",x"37db",x"b859",x"3581",x"3a1f",x"35a9",x"3362"),
(x"3a7b",x"4024",x"37fd",x"a3bb",x"3849",x"3ac0",x"35c1",x"3362",x"3a5d",x"4022",x"37db",x"b859",x"3581",x"3a1f",x"35a9",x"3362",x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351"),
(x"3a7b",x"4026",x"37e2",x"9c81",x"3a99",x"3885",x"35c1",x"3351",x"3a5d",x"4024",x"37cd",x"b609",x"3a62",x"3783",x"35aa",x"334e",x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341"),
(x"3a7b",x"4027",x"37c9",x"9987",x"3bd9",x"322d",x"35c1",x"3341",x"3a5c",x"4025",x"37b8",x"b4be",x"3ba1",x"2a04",x"35a8",x"333e",x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331"),
(x"3a7b",x"4027",x"37b3",x"a887",x"3bce",x"b2e4",x"35c0",x"3331",x"3a5c",x"4025",x"37a7",x"b4f8",x"3b04",x"b5db",x"35a6",x"3332",x"3a64",x"4024",x"3789",x"b533",x"3ac8",x"b6b3",x"35a9",x"3318"),
(x"3a54",x"4024",x"3782",x"3907",x"3a38",x"a553",x"365e",x"344b",x"3a5d",x"4022",x"3782",x"3856",x"3952",x"381b",x"3662",x"3443",x"3a56",x"4023",x"378c",x"3932",x"391d",x"3695",x"3664",x"344a"),
(x"3a5d",x"4022",x"3782",x"b718",x"3b28",x"2aae",x"35a3",x"3313",x"3a5f",x"4023",x"378b",x"b7bc",x"3afd",x"2a6c",x"35a4",x"331a",x"3a5a",x"4022",x"378b",x"b71a",x"3b19",x"2ff1",x"35a0",x"3319"),
(x"3a3b",x"3ff0",x"3752",x"bae0",x"aed4",x"37ff",x"365d",x"34ec",x"3a36",x"4002",x"3752",x"bab1",x"af0f",x"3849",x"3656",x"34ce",x"3a41",x"3ffb",x"376e",x"bab9",x"ac8e",x"384b",x"3665",x"34da"),
(x"3a41",x"3ffb",x"376e",x"b12d",x"21ae",x"3be4",x"363f",x"30d7",x"3a41",x"4001",x"376d",x"b03c",x"aa80",x"3beb",x"3641",x"30bf",x"3a4a",x"3fff",x"3770",x"ad3d",x"28c9",x"3bf7",x"3647",x"30ce"),
(x"3abb",x"3fef",x"3752",x"3b01",x"ac96",x"37a2",x"362b",x"33a9",x"3ab5",x"3ff8",x"376e",x"3afe",x"ac6c",x"37b0",x"3633",x"33c7",x"3abf",x"4002",x"3752",x"3b07",x"b070",x"374f",x"3623",x"33e8"),
(x"3aa4",x"4002",x"3770",x"2c6a",x"aa7d",x"3bf8",x"358a",x"34d2",x"3ab0",x"4002",x"376f",x"0e8d",x"a93f",x"3bfe",x"3581",x"34d2",x"3aa4",x"3ffc",x"3770",x"2938",x"1d6d",x"3bfe",x"3589",x"34c5"),
(x"3ade",x"404c",x"3752",x"3ac8",x"b025",x"381c",x"35f9",x"34dd",x"3acd",x"404b",x"3786",x"3af5",x"afa5",x"37a8",x"3610",x"34de",x"3ad3",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35fb",x"34ec"),
(x"3ad3",x"4051",x"3752",x"3a20",x"3711",x"3778",x"35fb",x"34ec",x"3ac7",x"404f",x"378d",x"3a12",x"37f9",x"36b2",x"3613",x"34eb",x"3acb",x"4053",x"3752",x"3846",x"3a11",x"35f5",x"35fd",x"34f4"),
(x"3acb",x"4053",x"3752",x"3846",x"3a11",x"35f5",x"35fd",x"34f4",x"3ac1",x"4051",x"378e",x"3609",x"3ae2",x"3579",x"3615",x"34f1",x"3ac3",x"4053",x"3752",x"af98",x"3bdd",x"3078",x"35ff",x"34f9"),
(x"3ade",x"404c",x"3752",x"3ac8",x"b025",x"381c",x"35f9",x"34dd",x"3ac7",x"403d",x"3752",x"3ad1",x"b46a",x"371a",x"360a",x"34b0",x"3acd",x"404b",x"3786",x"3af5",x"afa5",x"37a8",x"3610",x"34de"),
(x"3ac7",x"403d",x"3752",x"3ad1",x"b46a",x"371a",x"360a",x"34b0",x"3abf",x"4034",x"3752",x"3afe",x"b17b",x"3746",x"3612",x"3497",x"3abe",x"403d",x"3777",x"3af8",x"b403",x"36bf",x"3619",x"34b3"),
(x"3ac3",x"4053",x"3752",x"af98",x"3bdd",x"3078",x"35ff",x"34f9",x"3aab",x"4051",x"378e",x"b6eb",x"3b36",x"1c18",x"361c",x"34ff",x"3aa4",x"404f",x"3782",x"b85b",x"3ab4",x"a80e",x"361b",x"3507"),
(x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3ab7",x"4034",x"376d",x"25e3",x"adbf",x"3bf7",x"360e",x"333a"),
(x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3abe",x"403d",x"3777",x"a53f",x"b05f",x"3bec",x"3611",x"3305"),
(x"3acd",x"404b",x"3786",x"30f8",x"b10a",x"3bcd",x"3619",x"32ae",x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3ac7",x"404f",x"378d",x"2f46",x"b040",x"3be0",x"3613",x"3297"),
(x"3ac7",x"404f",x"378d",x"2f46",x"b040",x"3be0",x"3613",x"3297",x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3ac1",x"4051",x"378e",x"2d5b",x"a17a",x"3bf8",x"360e",x"328f"),
(x"3ac1",x"4051",x"378e",x"2d5b",x"a17a",x"3bf8",x"360e",x"328f",x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3ab6",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"3ab4",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3605",x"3292",x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3ab6",x"4051",x"378f",x"9da1",x"29fd",x"3bfd",x"3606",x"328c"),
(x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aab",x"4051",x"378e",x"ad32",x"a525",x"3bf8",x"35fe",x"3292"),
(x"3a9d",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"35f4",x"32a5",x"3aa6",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"3a9d",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"3aa2",x"404e",x"378c",x"a877",x"ae68",x"3bf4",x"35f7",x"32a1",x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3a9d",x"404e",x"378b",x"aeec",x"b1eb",x"3bd0",x"35f4",x"32a5"),
(x"3aa6",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3a9d",x"404a",x"3784",x"af8b",x"b19e",x"3bd1",x"35f4",x"32ba"),
(x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3aa6",x"403d",x"3777",x"2c2a",x"afe7",x"3beb",x"35fe",x"3305",x"3a9e",x"4045",x"377f",x"a7ce",x"b04a",x"3bec",x"35f6",x"32d9"),
(x"3aa6",x"403d",x"3777",x"2c2a",x"afe7",x"3beb",x"35fe",x"3305",x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b",x"3a9d",x"403d",x"3777",x"2bbb",x"ae16",x"3bf2",x"35f8",x"3309"),
(x"3aa6",x"403d",x"3777",x"2c2a",x"afe7",x"3beb",x"35fe",x"3305",x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"3aae",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3602",x"32d4",x"3aa8",x"4045",x"3780",x"3168",x"b087",x"3bcd",x"35fd",x"32d5",x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"3aa6",x"404a",x"3788",x"2c6f",x"b1f6",x"3bd7",x"35fb",x"32b8",x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7"),
(x"3aa8",x"404e",x"378c",x"3169",x"b278",x"3bb7",x"35fc",x"32a3",x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4"),
(x"3aaf",x"4050",x"378f",x"31a5",x"b517",x"3b73",x"3601",x"3296",x"3ab4",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3605",x"3292",x"3ab2",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3603",x"329c"),
(x"3ab4",x"4051",x"3790",x"2b8d",x"b837",x"3ac8",x"3605",x"3292",x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3ab6",x"4050",x"3787",x"a710",x"b98f",x"39bf",x"3606",x"329a"),
(x"3abd",x"4050",x"378f",x"ad72",x"b63e",x"3b55",x"360c",x"3294",x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b"),
(x"3ac2",x"404f",x"378d",x"b3a9",x"b4a4",x"3b69",x"3610",x"329a",x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1"),
(x"3ac6",x"404c",x"3788",x"b0d0",x"b03c",x"3bd6",x"3614",x"32ae",x"3ab7",x"403d",x"3776",x"b339",x"accc",x"3bc5",x"360c",x"3304",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"3ab4",x"403d",x"3773",x"adb8",x"ad34",x"3bf1",x"3609",x"3304",x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302"),
(x"3aaa",x"403e",x"3775",x"30b9",x"adbc",x"3be1",x"3602",x"3302",x"3aae",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3602",x"32d4",x"3ab4",x"403d",x"3773",x"adb8",x"ad34",x"3bf1",x"3609",x"3304"),
(x"3aae",x"4046",x"377a",x"2c32",x"b02f",x"3be9",x"3602",x"32d4",x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7",x"3ac2",x"404b",x"3782",x"b113",x"af65",x"3bd8",x"3610",x"32b0"),
(x"3aaa",x"404b",x"3782",x"3155",x"b185",x"3bc4",x"35fe",x"32b7",x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4",x"3abf",x"404e",x"3785",x"ae66",x"b276",x"3bcb",x"360d",x"32a1"),
(x"3aac",x"404e",x"3787",x"3200",x"b38a",x"3ba0",x"35ff",x"32a4",x"3ab2",x"404f",x"3787",x"3370",x"b70b",x"3af0",x"3603",x"329c",x"3abb",x"404f",x"3787",x"b079",x"b50b",x"3b82",x"360a",x"329b"),
(x"3a9c",x"403d",x"3783",x"3b8f",x"ab5c",x"3527",x"35a7",x"34a3",x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a97",x"4045",x"3794",x"3bbc",x"287e",x"3408",x"35a6",x"348a",x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a9c",x"404a",x"3790",x"3b17",x"ade0",x"3741",x"35ac",x"347b",x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a95",x"404d",x"37a3",x"3bd3",x"a9fd",x"3273",x"35a4",x"3474",x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470",x"3a95",x"404e",x"37b6",x"393b",x"b9e8",x"313a",x"359f",x"346f",x"3a9c",x"404f",x"37aa",x"39e5",x"b8ae",x"3566",x"35a5",x"346b"),
(x"3a95",x"404e",x"37b6",x"393b",x"b9e8",x"313a",x"359f",x"346f",x"3a95",x"404e",x"37c1",x"3a55",x"b865",x"b441",x"359c",x"346e",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468"),
(x"3a95",x"404e",x"37c1",x"3a55",x"b865",x"b441",x"359c",x"346e",x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e",x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477"),
(x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477",x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485"),
(x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485",x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f"),
(x"3a9a",x"403d",x"37b2",x"3bec",x"ac1f",x"2fcd",x"3595",x"349f",x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f",x"3a99",x"4031",x"3795",x"3be2",x"acf4",x"30cb",x"3598",x"34c3"),
(x"3a9b",x"403d",x"37a7",x"3bbc",x"2e00",x"b38d",x"3599",x"349f",x"3a9a",x"403d",x"37b2",x"3bec",x"ac1f",x"2fcd",x"3595",x"349f",x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485"),
(x"3a9b",x"4046",x"37c6",x"3b50",x"30fc",x"b5fd",x"3592",x"3485",x"3a9b",x"4045",x"37d1",x"3bf6",x"a9b5",x"2d99",x"358e",x"3485",x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477"),
(x"3a9b",x"404a",x"37d4",x"3b43",x"293f",x"b6a9",x"3590",x"3477",x"3a9b",x"404a",x"37de",x"3be7",x"a00b",x"30f0",x"358d",x"3476",x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"3a9a",x"404d",x"37dc",x"3bd6",x"2b52",x"322d",x"3590",x"346c",x"3a9b",x"4050",x"37cc",x"3be3",x"2d8f",x"3091",x"3598",x"3466",x"3a9b",x"404d",x"37d2",x"3bb1",x"ad7d",x"b42c",x"3594",x"346e"),
(x"3a9b",x"4050",x"37cc",x"3be3",x"2d8f",x"3091",x"3598",x"3466",x"3a9c",x"4050",x"37b8",x"3bf8",x"2c16",x"2b31",x"35a1",x"3466",x"3a9c",x"404f",x"37c8",x"3aa6",x"b6d3",x"b5b4",x"3599",x"3469"),
(x"3a9c",x"4050",x"37b8",x"3bf8",x"2c16",x"2b31",x"35a1",x"3466",x"3a9c",x"4050",x"37a7",x"3bff",x"232b",x"2518",x"35a7",x"3469",x"3a9c",x"4050",x"37b7",x"3a3a",x"b904",x"a765",x"35a0",x"3468"),
(x"3a9c",x"404f",x"37aa",x"39e5",x"b8ae",x"3566",x"35a5",x"346b",x"3a9c",x"4050",x"37a7",x"3bff",x"232b",x"2518",x"35a7",x"3469",x"3a9c",x"404d",x"3799",x"3a98",x"b4d2",x"37a9",x"35ab",x"3472"),
(x"3a9d",x"404a",x"3784",x"3bd5",x"a532",x"3275",x"35b1",x"347c",x"3a9c",x"404a",x"3790",x"3b17",x"ade0",x"3741",x"35ac",x"347b",x"3a9c",x"404e",x"378e",x"3bf3",x"a432",x"2ede",x"35af",x"3471"),
(x"3a9c",x"404a",x"3790",x"3b17",x"ade0",x"3741",x"35ac",x"347b",x"3a9d",x"404a",x"3784",x"3bd5",x"a532",x"3275",x"35b1",x"347c",x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b"),
(x"3a9c",x"4045",x"378b",x"3aba",x"ab10",x"384d",x"35ab",x"348b",x"3a9e",x"4045",x"377f",x"3bc6",x"a6c8",x"337e",x"35b0",x"348c",x"3a9c",x"403d",x"3783",x"3b8f",x"ab5c",x"3527",x"35a7",x"34a3"),
(x"3a99",x"403d",x"379f",x"3bf7",x"2d6b",x"a836",x"359d",x"34a0",x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a99",x"4031",x"378d",x"3bfd",x"1418",x"2a73",x"359b",x"34c3"),
(x"3a9a",x"403d",x"378a",x"3bb7",x"a074",x"3436",x"35a4",x"34a2",x"3a99",x"403d",x"379f",x"3bf7",x"2d6b",x"a836",x"359d",x"34a0",x"3a97",x"4045",x"3794",x"3bbc",x"287e",x"3408",x"35a6",x"348a"),
(x"3a97",x"4045",x"3794",x"3bbc",x"287e",x"3408",x"35a6",x"348a",x"3a95",x"4046",x"37ba",x"3bd9",x"2f80",x"b0f2",x"3599",x"3485",x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c"),
(x"3a96",x"404a",x"3798",x"3b91",x"abb4",x"3517",x"35a7",x"347c",x"3a95",x"404a",x"37c9",x"3bca",x"2d2f",x"b2c3",x"3597",x"3478",x"3a95",x"404d",x"37a3",x"3bd3",x"a9fd",x"3273",x"35a4",x"3474"),
(x"3a95",x"404d",x"37a3",x"3bd3",x"a9fd",x"3273",x"35a4",x"3474",x"3a95",x"404d",x"37c7",x"3b5f",x"ae12",x"b605",x"3599",x"3471",x"3a95",x"404e",x"37ac",x"3ad8",x"b658",x"3550",x"35a2",x"3470"),
(x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a9a",x"403d",x"37b2",x"386e",x"b47a",x"3a45",x"367a",x"29b1",x"3a7c",x"4031",x"37c0",x"9bc8",x"b48d",x"3bab",x"365d",x"2ab9"),
(x"3a9a",x"403d",x"37b2",x"386e",x"b47a",x"3a45",x"367a",x"29b1",x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a9b",x"4045",x"37d1",x"3856",x"b5aa",x"3a18",x"3678",x"28cc"),
(x"3a9b",x"4045",x"37d1",x"3856",x"b5aa",x"3a18",x"3678",x"28cc",x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a9b",x"404a",x"37de",x"3892",x"b07e",x"3a77",x"3675",x"284f"),
(x"3a9b",x"404a",x"37de",x"3892",x"b07e",x"3a77",x"3675",x"284f",x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a9a",x"404d",x"37dc",x"3809",x"374a",x"39de",x"3673",x"27ef"),
(x"3a7b",x"4050",x"37fd",x"a32b",x"38f3",x"3a48",x"365b",x"2806",x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e",x"3a9a",x"404d",x"37dc",x"3809",x"374a",x"39de",x"3673",x"27ef"),
(x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e",x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709",x"3a9b",x"4050",x"37cc",x"34ee",x"3aeb",x"3653",x"3673",x"275d"),
(x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709",x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c",x"3a9c",x"4050",x"37b8",x"3361",x"3bc7",x"282c",x"3674",x"26df"),
(x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c",x"3a93",x"4050",x"379c",x"3458",x"3b15",x"b609",x"366f",x"2623",x"3a9c",x"4050",x"37a7",x"3362",x"3b62",x"b4ea",x"3676",x"2679"),
(x"3aa4",x"404f",x"3782",x"b85b",x"3ab4",x"a80e",x"361b",x"3507",x"3aa2",x"404e",x"378c",x"b8cb",x"39b0",x"35e1",x"3620",x"3508",x"3a9c",x"404e",x"3786",x"b75f",x"39e5",x"37e9",x"3620",x"350c"),
(x"3a99",x"404e",x"378b",x"3818",x"3ad2",x"ae9f",x"3676",x"25ba",x"3a9c",x"404e",x"3786",x"35de",x"3b08",x"34dc",x"3679",x"2599",x"3a9c",x"404e",x"378e",x"362d",x"3aa4",x"b66f",x"3679",x"25cc"),
(x"3a31",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"35f8",x"2da1",x"3a2a",x"404b",x"3786",x"bae1",x"b000",x"37eb",x"35f5",x"2dd3",x"3a24",x"4051",x"3752",x"ba20",x"3711",x"3778",x"35e0",x"2d9e"),
(x"3a37",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"35fa",x"2d8a",x"3a31",x"404f",x"378d",x"ba12",x"37fa",x"36b2",x"35f8",x"2da1",x"3a2d",x"4053",x"3752",x"b846",x"3a11",x"35f5",x"35e2",x"2d7f"),
(x"3a42",x"4051",x"378f",x"25dc",x"3bcd",x"330b",x"35fe",x"2d6c",x"3a37",x"4051",x"378e",x"b609",x"3ae2",x"3579",x"35fa",x"2d8a",x"3a35",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35e4",x"2d68"),
(x"3a1a",x"404c",x"3752",x"bac8",x"b025",x"381c",x"35de",x"2dda",x"3a2a",x"404b",x"3786",x"bae1",x"b000",x"37eb",x"35f5",x"2dd3",x"3a31",x"403d",x"3752",x"bab4",x"b44c",x"3799",x"35f0",x"2e8e"),
(x"3a31",x"403d",x"3752",x"bab4",x"b44c",x"3799",x"35f0",x"2e8e",x"3a3b",x"403c",x"3775",x"bab0",x"b345",x"37fd",x"35ff",x"2e87",x"3a36",x"4034",x"3752",x"baac",x"b05e",x"3846",x"35f7",x"2ef0"),
(x"3a35",x"4053",x"3752",x"2f98",x"3bdd",x"3078",x"35e4",x"2d68",x"3a54",x"404f",x"3782",x"385d",x"3ab3",x"a49b",x"3600",x"2d31",x"3a4d",x"4051",x"378e",x"36eb",x"3b36",x"1c18",x"3601",x"2d50"),
(x"3a41",x"403d",x"3776",x"331d",x"aca2",x"3bc7",x"3662",x"2cd4",x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a3b",x"403c",x"3775",x"adad",x"b0c1",x"3be1",x"3667",x"2cd0"),
(x"3a41",x"403d",x"3776",x"331d",x"aca2",x"3bc7",x"3662",x"2cd4",x"3a3b",x"403c",x"3775",x"adad",x"b0c1",x"3be1",x"3667",x"2cd0",x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8",x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83",x"3a31",x"404f",x"378d",x"af46",x"b040",x"3be0",x"3663",x"2db2"),
(x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4",x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8",x"3a37",x"4051",x"378e",x"ad5b",x"a17a",x"3bf8",x"365d",x"2dbf"),
(x"3a43",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3654",x"2db4",x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4",x"3a42",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3655",x"2dc0"),
(x"3a43",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3654",x"2db4",x"3a42",x"4051",x"378f",x"1da1",x"29fd",x"3bfd",x"3655",x"2dc0",x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa",x"3a4d",x"4051",x"378e",x"2d32",x"a525",x"3bf8",x"364d",x"2db2",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"3a5a",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"3645",x"2d87",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f",x"3a56",x"404e",x"378c",x"2877",x"ae68",x"3bf4",x"3647",x"2d91"),
(x"3a5b",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"3a52",x"404a",x"3788",x"ac6d",x"b1f6",x"3bd7",x"364c",x"2d65",x"3a5a",x"404e",x"378b",x"2eec",x"b1eb",x"3bd0",x"3645",x"2d87"),
(x"3a52",x"404a",x"3788",x"ac6d",x"b1f6",x"3bd7",x"364c",x"2d65",x"3a5b",x"404a",x"3784",x"2f8b",x"b19e",x"3bd1",x"3646",x"2d5e",x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c",x"3a5a",x"4045",x"377f",x"27ce",x"b04a",x"3bec",x"364a",x"2d20",x"3a52",x"403d",x"3777",x"ac2f",x"afb9",x"3bec",x"3655",x"2cce"),
(x"3a52",x"403d",x"3777",x"ac2f",x"afb9",x"3bec",x"3655",x"2cce",x"3a5a",x"403d",x"3777",x"aa04",x"ae02",x"3bf4",x"364f",x"2cc3",x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c"),
(x"3a52",x"403d",x"3777",x"ac2f",x"afb9",x"3bec",x"3655",x"2cce",x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c"),
(x"3a52",x"404a",x"3788",x"ac6d",x"b1f6",x"3bd7",x"364c",x"2d65",x"3a50",x"4045",x"3780",x"b168",x"b087",x"3bcd",x"3651",x"2d2c",x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68"),
(x"3a52",x"404a",x"3788",x"ac6d",x"b1f6",x"3bd7",x"364c",x"2d65",x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68",x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f"),
(x"3a50",x"404e",x"378c",x"b169",x"b278",x"3bb7",x"364c",x"2d8f",x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d",x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa"),
(x"3a49",x"4050",x"378f",x"b1a5",x"b517",x"3b73",x"3650",x"2daa",x"3a46",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3654",x"2d9f",x"3a43",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3654",x"2db4"),
(x"3a43",x"4051",x"3790",x"ab8d",x"b837",x"3ac8",x"3654",x"2db4",x"3a42",x"4050",x"3787",x"270a",x"b98f",x"39bf",x"3656",x"2da5",x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4"),
(x"3a3b",x"4050",x"378f",x"2d73",x"b63f",x"3b55",x"365b",x"2db4",x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8"),
(x"3a36",x"404f",x"378d",x"33a9",x"b4a4",x"3b69",x"3660",x"2da8",x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83"),
(x"3a31",x"404c",x"3788",x"2ed7",x"b0dc",x"3bdc",x"3665",x"2d83",x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a41",x"403d",x"3776",x"331d",x"aca2",x"3bc7",x"3662",x"2cd4"),
(x"3a54",x"4034",x"3770",x"ac25",x"ab90",x"3bf8",x"365a",x"2c5c",x"3a48",x"4034",x"376f",x"a5ae",x"abef",x"3bfb",x"3663",x"2c62",x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5"),
(x"3a4d",x"403e",x"3775",x"b0a6",x"ad8a",x"3be2",x"3658",x"2cd5",x"3a44",x"403d",x"3773",x"2dae",x"ad20",x"3bf1",x"3660",x"2cd4",x"3a4a",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3656",x"2d31"),
(x"3a4a",x"4046",x"377a",x"ac32",x"b02f",x"3be9",x"3656",x"2d31",x"3a35",x"404b",x"3782",x"3113",x"af65",x"3bd8",x"3661",x"2d7d",x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68"),
(x"3a4e",x"404b",x"3782",x"b154",x"b185",x"3bc4",x"3650",x"2d68",x"3a39",x"404e",x"3785",x"2e64",x"b275",x"3bcb",x"365d",x"2d9b",x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d"),
(x"3a4c",x"404e",x"3787",x"b200",x"b38a",x"3ba0",x"3650",x"2d8d",x"3a3d",x"404f",x"3787",x"3079",x"b50b",x"3b82",x"365a",x"2da4",x"3a46",x"404f",x"3787",x"b370",x"b70b",x"3af0",x"3654",x"2d9f"),
(x"3a61",x"4045",x"3794",x"bbd9",x"292f",x"3209",x"35f5",x"33a8",x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8",x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"3a61",x"4045",x"3794",x"bbd9",x"292f",x"3209",x"35f5",x"33a8",x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b"),
(x"3a62",x"404d",x"37a3",x"bbda",x"aea9",x"311c",x"35f5",x"337c",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"3a62",x"404d",x"37a3",x"bbda",x"aea9",x"311c",x"35f5",x"337c",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377",x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373",x"3a5c",x"404f",x"37aa",x"ba13",x"b891",x"34fa",x"35f4",x"336a",x"3a61",x"404f",x"37b7",x"b977",x"b9c7",x"2ebe",x"35fa",x"336e"),
(x"3a61",x"404f",x"37b7",x"b977",x"b9c7",x"2ebe",x"35fa",x"336e",x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e"),
(x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b"),
(x"3a5f",x"403d",x"37a1",x"bbf5",x"2dc9",x"aa2e",x"3600",x"33d2",x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1"),
(x"3a5c",x"4030",x"378d",x"bbfe",x"28c2",x"2138",x"3602",x"340f",x"3a5d",x"403d",x"37a5",x"bbc3",x"2ec2",x"b2f6",x"3601",x"33d1",x"3a5d",x"4030",x"3797",x"bbf6",x"a3bb",x"2e0a",x"3606",x"340f"),
(x"3a5d",x"4045",x"37d0",x"bc00",x"9fe2",x"8000",x"360b",x"339c",x"3a5d",x"403d",x"37b0",x"bbff",x"a3ef",x"2511",x"3606",x"33d1",x"3a5d",x"4046",x"37c6",x"bb29",x"3144",x"b6a0",x"3608",x"339b"),
(x"3a5c",x"404a",x"37dc",x"bbfd",x"14ea",x"a9d6",x"360c",x"337d",x"3a5d",x"4045",x"37d0",x"bc00",x"9fe2",x"8000",x"360b",x"339c",x"3a5d",x"404a",x"37d2",x"bafe",x"2b1d",x"b7b8",x"3608",x"3380"),
(x"3a5d",x"404d",x"37db",x"bbff",x"9018",x"a31d",x"3608",x"336a",x"3a5c",x"404a",x"37dc",x"bbfd",x"14ea",x"a9d6",x"360c",x"337d",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f"),
(x"3a5d",x"404d",x"37db",x"bbff",x"9018",x"a31d",x"3608",x"336a",x"3a5d",x"404d",x"37d0",x"bb62",x"afb4",x"b5d8",x"3604",x"336f",x"3a5d",x"4050",x"37cd",x"bbfa",x"2874",x"2c13",x"3601",x"3360"),
(x"3a5d",x"4050",x"37cd",x"bbfa",x"2874",x"2c13",x"3601",x"3360",x"3a5c",x"404f",x"37c9",x"bb31",x"b5e3",x"b398",x"3600",x"3366",x"3a5c",x"4050",x"37b8",x"bbfa",x"2a69",x"2a66",x"35f8",x"3360"),
(x"3a5c",x"4050",x"37b8",x"bbfa",x"2a69",x"2a66",x"35f8",x"3360",x"3a5c",x"404f",x"37b7",x"ba7d",x"b8a9",x"a953",x"35f9",x"3365",x"3a5c",x"4050",x"37a7",x"bbff",x"20dd",x"2604",x"35f2",x"3366"),
(x"3a5b",x"404e",x"378e",x"bbf3",x"a432",x"2f1d",x"35ea",x"3376",x"3a5c",x"4050",x"37a7",x"bbff",x"20dd",x"2604",x"35f2",x"3366",x"3a5b",x"404d",x"3798",x"ba9c",x"b4c1",x"37a5",x"35ee",x"3377"),
(x"3a5b",x"404a",x"3784",x"bbd5",x"a532",x"3275",x"35e9",x"338d",x"3a5b",x"404e",x"378e",x"bbf3",x"a432",x"2f1d",x"35ea",x"3376",x"3a5c",x"404a",x"3790",x"bb10",x"ad8c",x"3760",x"35ed",x"338b"),
(x"3a5a",x"4045",x"377f",x"bbc5",x"a6cf",x"3387",x"35eb",x"33ac",x"3a5b",x"404a",x"3784",x"bbd5",x"a532",x"3275",x"35e9",x"338d",x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa"),
(x"3a5c",x"4045",x"378b",x"babf",x"ab14",x"3846",x"35ef",x"33aa",x"3a5c",x"403d",x"3782",x"bb88",x"abb1",x"354b",x"35f4",x"33d9",x"3a5a",x"4045",x"377f",x"bbc5",x"a6cf",x"3387",x"35eb",x"33ac"),
(x"3a5f",x"403d",x"37a1",x"bbf5",x"2dc9",x"aa2e",x"3600",x"33d2",x"3a5c",x"4030",x"378d",x"bbfe",x"28c2",x"2138",x"3602",x"340f",x"3a5e",x"403d",x"378a",x"bbd9",x"243f",x"3220",x"35f7",x"33d8"),
(x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a5f",x"403d",x"37a1",x"bbf5",x"2dc9",x"aa2e",x"3600",x"33d2",x"3a61",x"4045",x"3794",x"bbd9",x"292f",x"3209",x"35f5",x"33a8"),
(x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a62",x"4046",x"37be",x"bbdb",x"2f8d",x"b0af",x"3602",x"339b",x"3a61",x"404a",x"3798",x"bba3",x"a84d",x"34bc",x"35f2",x"338b"),
(x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a63",x"404a",x"37c9",x"bbce",x"2c74",x"b2a7",x"3603",x"3383",x"3a62",x"404d",x"37a3",x"bbda",x"aea9",x"311c",x"35f5",x"337c"),
(x"3a61",x"404e",x"37c3",x"ba5f",x"b7e4",x"b595",x"35fe",x"336e",x"3a62",x"404d",x"37c9",x"bb8e",x"aeb0",x"b4f9",x"3601",x"3374",x"3a62",x"404e",x"37ac",x"bb0a",x"b677",x"33fe",x"35f6",x"3373"),
(x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a7c",x"4031",x"37c0",x"9bc8",x"b48d",x"3bab",x"365d",x"2ab9",x"3a5d",x"403d",x"37b0",x"b860",x"b445",x"3a59",x"363e",x"29b6"),
(x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a7b",x"403d",x"37dc",x"a1d6",x"b62a",x"3b61",x"365c",x"298f",x"3a5d",x"4045",x"37d0",x"b86c",x"b560",x"3a19",x"3640",x"28d0"),
(x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a7d",x"4046",x"3800",x"a2cf",x"b59c",x"3b7d",x"365c",x"28a9",x"3a5c",x"404a",x"37dc",x"b889",x"b0d3",x"3a7a",x"3643",x"2852"),
(x"3a7b",x"4050",x"37fd",x"a32b",x"38f3",x"3a48",x"365b",x"2806",x"3a7c",x"404b",x"3804",x"a194",x"2bfc",x"3bfb",x"365c",x"284f",x"3a5d",x"404d",x"37db",x"b837",x"36a0",x"39ef",x"3644",x"2800"),
(x"3a7b",x"4050",x"37fd",x"a32b",x"38f3",x"3a48",x"365b",x"2806",x"3a5d",x"404d",x"37db",x"b837",x"36a0",x"39ef",x"3644",x"2800",x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e"),
(x"3a7b",x"4051",x"37e2",x"9bc8",x"3b01",x"37bb",x"365b",x"278e",x"3a5d",x"4050",x"37cd",x"b534",x"3ad5",x"367a",x"3644",x"2773",x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709"),
(x"3a7b",x"4052",x"37c9",x"9881",x"3be6",x"3102",x"365b",x"2709",x"3a5c",x"4050",x"37b8",x"b3c4",x"3bc1",x"28ed",x"3642",x"26f2",x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c"),
(x"3a7b",x"4052",x"37b3",x"a75f",x"3bdf",x"b19a",x"365b",x"268c",x"3a5c",x"4050",x"37a7",x"b42d",x"3b51",x"b4ec",x"3641",x"268d",x"3a64",x"404f",x"3789",x"b469",x"3b25",x"b5af",x"3644",x"25c3"),
(x"3a54",x"404f",x"3782",x"385d",x"3ab3",x"a49b",x"3600",x"2d31",x"3a5d",x"404e",x"3782",x"37ca",x"39ef",x"375f",x"3603",x"2d14",x"3a56",x"404e",x"378c",x"38b4",x"39be",x"35f4",x"3605",x"2d2d"),
(x"3a5d",x"404e",x"3782",x"b5ed",x"3b6c",x"2997",x"363e",x"2598",x"3a5f",x"404e",x"378b",x"b682",x"3b4c",x"297d",x"363f",x"25d0",x"3a5a",x"404e",x"378b",x"b5f3",x"3b61",x"2ea6",x"363c",x"25cf"),
(x"3a3b",x"402c",x"3752",x"bada",x"b039",x"37f8",x"35fe",x"2f4f",x"3a36",x"4034",x"3752",x"baac",x"b05e",x"3846",x"35f7",x"2ef0",x"3a41",x"4030",x"376e",x"bab7",x"ada6",x"384a",x"3606",x"2f15"),
(x"3a41",x"4030",x"376e",x"b12d",x"2310",x"3be4",x"366a",x"2c3f",x"3a41",x"4033",x"376d",x"b03b",x"ac08",x"3be9",x"3668",x"2c64",x"3a4a",x"4032",x"3770",x"acfa",x"29bc",x"3bf7",x"3663",x"2c4b"),
(x"3abb",x"402b",x"3752",x"3aff",x"adb0",x"379f",x"3619",x"347e",x"3ab5",x"402f",x"376e",x"3afb",x"ad7c",x"37ae",x"3622",x"348b",x"3abf",x"4034",x"3752",x"3afe",x"b17b",x"3746",x"3612",x"3497"),
(x"3aa4",x"4034",x"3770",x"2c95",x"ac08",x"3bf6",x"3600",x"333b",x"3ab0",x"4034",x"376f",x"27bb",x"a9c9",x"3bfc",x"3609",x"333a",x"3aa4",x"4031",x"3770",x"2935",x"1ec2",x"3bfe",x"3601",x"3350"),
(x"3a4e",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"3a40",x"3f95",x"37cf",x"bafd",x"36b2",x"b3e9",x"3562",x"3530",x"3a2b",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518"),
(x"3a4e",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"3a40",x"3f95",x"37cf",x"b33d",x"35ac",x"3b41",x"3604",x"30cf"),
(x"3aa0",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4",x"3ab1",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce",x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"3abe",x"3f47",x"3752",x"0000",x"0000",x"3c00",x"35b6",x"2b4f",x"3ab4",x"3f46",x"3752",x"330f",x"b68f",x"3b14",x"35af",x"2b2d",x"3ac8",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88"),
(x"3ab1",x"3f95",x"37ce",x"373e",x"b495",x"3ac1",x"358b",x"2d70",x"3ad7",x"3f58",x"3752",x"374a",x"b488",x"3ac0",x"35c3",x"2c17",x"3a9c",x"3f77",x"37bd",x"367e",x"b50c",x"3adc",x"3585",x"2cb9"),
(x"3ad7",x"3f58",x"3752",x"3b2b",x"3633",x"b2e4",x"35e5",x"2c0c",x"3ab1",x"3f95",x"37ce",x"3af6",x"36ac",x"b42c",x"359e",x"2d3c",x"3ac4",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91"),
(x"3a54",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"3a3a",x"3f46",x"3752",x"b179",x"b6cc",x"3b1c",x"350b",x"349a",x"3a31",x"3f48",x"3752",x"b5a1",x"b590",x"3af3",x"3506",x"349f"),
(x"3a40",x"3f95",x"37cf",x"ba59",x"b59a",x"37f3",x"353f",x"350c",x"3a54",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"3a17",x"3f58",x"3752",x"b6ba",x"b4d8",x"3ad7",x"34fb",x"34bd"),
(x"3a7a",x"3f4b",x"380b",x"3b6a",x"b5fa",x"a853",x"35e2",x"2e9e",x"3a78",x"3f49",x"380d",x"3ac4",x"b843",x"a386",x"35e1",x"2e92",x"3a7c",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1"),
(x"3a78",x"3f49",x"382e",x"b94b",x"b9fe",x"2025",x"3582",x"3498",x"3a78",x"3f49",x"380d",x"ba6f",x"b8c0",x"a6fd",x"356a",x"3496",x"3a75",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c"),
(x"3a7a",x"3f4b",x"380b",x"3b6a",x"b5fa",x"a853",x"35e2",x"2e9e",x"3a7c",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1",x"3a9c",x"3f77",x"37bd",x"3b7c",x"b5a3",x"a1ae",x"3602",x"2fb5"),
(x"3a7c",x"3f4b",x"382c",x"38c7",x"30be",x"3a4d",x"35d2",x"31ac",x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"3ab1",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce"),
(x"3a40",x"3f95",x"37cf",x"ba59",x"b59a",x"37f3",x"353f",x"350c",x"3a75",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c",x"3a54",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd"),
(x"3a75",x"3f4b",x"382c",x"b89c",x"310b",x"3a6a",x"35d7",x"31ad",x"3a40",x"3f95",x"37cf",x"b33d",x"35ac",x"3b41",x"3604",x"30cf",x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad"),
(x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"3a7c",x"3f4b",x"382c",x"38c7",x"30be",x"3a4d",x"35d2",x"31ac",x"3a78",x"3f49",x"382e",x"2467",x"b509",x"3b97",x"35d4",x"31b1"),
(x"3a75",x"3f4b",x"382c",x"b89c",x"310b",x"3a6a",x"35d7",x"31ad",x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"3a78",x"3f49",x"382e",x"2467",x"b509",x"3b97",x"35d4",x"31b1"),
(x"3a4e",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"3a78",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"3aa0",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4",x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"3a78",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1"),
(x"3a78",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"3a4e",x"3fa2",x"37bf",x"32c1",x"37e3",x"3ac0",x"35fa",x"30a7",x"3a6b",x"3fa3",x"37a0",x"363d",x"3811",x"3a24",x"35e2",x"3096"),
(x"3a78",x"3f91",x"37c3",x"a24c",x"38b9",x"3a74",x"35d6",x"30d1",x"3a8d",x"3fa2",x"379c",x"b829",x"38f7",x"38b1",x"35c6",x"3094",x"3aa0",x"3fa2",x"37c0",x"b2af",x"3812",x"3aae",x"35b3",x"30a4"),
(x"3a8d",x"3fa2",x"379c",x"38d4",x"376b",x"b92f",x"35ad",x"2dca",x"3a96",x"3f82",x"3752",x"381e",x"3818",x"b980",x"35d8",x"2d45",x"3aa0",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a"),
(x"3a6b",x"3fa3",x"37a0",x"b70f",x"36eb",x"ba4a",x"3560",x"355b",x"3a4e",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"3a4f",x"3f71",x"3752",x"b43c",x"3773",x"bac1",x"3517",x"3533"),
(x"3a40",x"3f95",x"37cf",x"bafd",x"36b2",x"b3e9",x"3562",x"3530",x"3a17",x"3f58",x"3752",x"bb05",x"36a0",x"b3ae",x"3504",x"34fb",x"3a2b",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518"),
(x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151",x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"3a40",x"3f95",x"37cf",x"b33d",x"35ac",x"3b41",x"3604",x"30cf"),
(x"3ab1",x"3f95",x"37ce",x"336a",x"35ac",x"3b3f",x"35a7",x"30ce",x"3a78",x"3f4b",x"382f",x"1481",x"35aa",x"3b7b",x"35d4",x"31ad",x"3a77",x"3f6d",x"3814",x"2138",x"3720",x"3b29",x"35d6",x"3151"),
(x"3ab4",x"3f46",x"3752",x"330f",x"b68f",x"3b14",x"35af",x"2b2d",x"3a9c",x"3f77",x"37bd",x"367e",x"b50c",x"3adc",x"3585",x"2cb9",x"3ac8",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88"),
(x"3ad7",x"3f58",x"3752",x"374a",x"b488",x"3ac0",x"35c3",x"2c17",x"3ac8",x"3f4b",x"3752",x"35a3",x"b57a",x"3af7",x"35bb",x"2b88",x"3a9c",x"3f77",x"37bd",x"367e",x"b50c",x"3adc",x"3585",x"2cb9"),
(x"3ab1",x"3f95",x"37ce",x"3af6",x"36ac",x"b42c",x"359e",x"2d3c",x"3aa0",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a",x"3ac4",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91"),
(x"3a54",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd",x"3a31",x"3f48",x"3752",x"b5a1",x"b590",x"3af3",x"3506",x"349f",x"3a17",x"3f58",x"3752",x"b6ba",x"b4d8",x"3ad7",x"34fb",x"34bd"),
(x"3a78",x"3f49",x"380d",x"3ac4",x"b843",x"a386",x"35e1",x"2e92",x"3a78",x"3f49",x"382e",x"3a6c",x"b8c3",x"9624",x"35c9",x"2e91",x"3a7c",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1"),
(x"3a78",x"3f49",x"380d",x"ba6f",x"b8bf",x"a6fd",x"356a",x"3496",x"3a77",x"3f4b",x"380c",x"bb52",x"b656",x"ac81",x"3569",x"3499",x"3a75",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c"),
(x"3a7c",x"3f4b",x"382c",x"3b77",x"b5bd",x"a1bc",x"35ca",x"2ea1",x"3ab1",x"3f95",x"37ce",x"3b84",x"b57a",x"175f",x"35fa",x"3035",x"3a9c",x"3f77",x"37bd",x"3b7c",x"b5a3",x"a1ae",x"3602",x"2fb5"),
(x"3a75",x"3f4b",x"382c",x"bb77",x"b5bc",x"a018",x"3580",x"349c",x"3a77",x"3f4b",x"380c",x"bb52",x"b656",x"ac81",x"3569",x"3499",x"3a54",x"3f78",x"37bb",x"b9f0",x"b62d",x"3862",x"353e",x"34dd"),
(x"3a96",x"3f82",x"3752",x"381e",x"3818",x"b980",x"35d8",x"2d45",x"3ac4",x"3f6e",x"3752",x"39c9",x"37db",x"b7c2",x"35db",x"2c91",x"3aa0",x"3fa2",x"37c0",x"38f9",x"380e",x"b8c6",x"359d",x"2d9a"),
(x"3a4e",x"3fa2",x"37bf",x"b724",x"37d3",x"b9fe",x"3569",x"3545",x"3a2b",x"3f6d",x"3752",x"b8ff",x"3817",x"b8b8",x"3518",x"3518",x"3a4f",x"3f71",x"3752",x"b43c",x"3773",x"bac1",x"3517",x"3533"),
(x"3a2c",x"34b8",x"36fb",x"3c00",x"0000",x"0000",x"35f8",x"38f3",x"3a2c",x"3cc1",x"36fb",x"3c00",x"0000",x"0000",x"35f8",x"3a68",x"3a2c",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"360d",x"38f3"),
(x"2c34",x"34b8",x"368e",x"bc00",x"8000",x"0000",x"383c",x"1cef",x"2c34",x"3cc1",x"368e",x"bc00",x"8000",x"0000",x"383c",x"3508",x"2c34",x"34b8",x"36fb",x"bc00",x"8000",x"0000",x"385a",x"1cef"),
(x"3193",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3a04",x"3838",x"394e",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3af7",x"3838",x"3193",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3a04",x"3832"),
(x"3a2c",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"39b1",x"3bdb",x"2c34",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"38eb",x"3bdb",x"3a2c",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"39b1",x"3bf4"),
(x"2c34",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"38ea",x"3bd3",x"3a2c",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"39b0",x"3bd3",x"2c34",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"38ea",x"3bb9"),
(x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93",x"3a2c",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"397d",x"3962",x"376a",x"36fb",x"0000",x"0000",x"3c00",x"3aa3",x"39b1"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"3009",x"39cc",x"36fb",x"0000",x"0000",x"3c00",x"39f1",x"3a03",x"3004",x"39d4",x"36fb",x"868d",x"0000",x"3c00",x"39f1",x"3a04"),
(x"394e",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"39a2",x"3a2c",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"397d",x"3193",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"39a2"),
(x"394e",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"3a6d",x"3193",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"3a6d",x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93"),
(x"3193",x"36aa",x"36d0",x"0000",x"0000",x"3c00",x"31b2",x"3adb",x"3193",x"3c44",x"36d0",x"0000",x"0000",x"3c00",x"31b2",x"3bf9",x"394e",x"36aa",x"36d0",x"0000",x"0000",x"3c00",x"3468",x"3adb"),
(x"3193",x"36e5",x"36fb",x"3c00",x"0000",x"0000",x"3a31",x"34c6",x"3193",x"370d",x"36e5",x"3c00",x"0000",x"0000",x"3a26",x"34d1",x"3193",x"36aa",x"36d0",x"3c00",x"0000",x"0000",x"3a40",x"34db"),
(x"394e",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3b7d",x"35b9",x"3193",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3af4",x"35b9",x"394e",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3b7d",x"35cd"),
(x"3141",x"3c25",x"36fb",x"396d",x"9af6",x"39e0",x"355f",x"3742",x"316f",x"3c38",x"36fb",x"39bc",x"b304",x"394a",x"355b",x"372f",x"3193",x"3c28",x"36d7",x"394c",x"a074",x"39fd",x"3552",x"373f"),
(x"3193",x"36e5",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"39a7",x"3193",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"39a2",x"3160",x"3716",x"36fb",x"0000",x"0000",x"3c00",x"39ff",x"39ab"),
(x"3193",x"3c37",x"36e4",x"3a1e",x"b322",x"38d5",x"3554",x"3730",x"316f",x"3c38",x"36fb",x"39bc",x"b304",x"394a",x"355b",x"372f",x"3193",x"3c41",x"36fb",x"39d6",x"b5ae",x"38ac",x"3558",x"3725"),
(x"3193",x"36aa",x"36d0",x"3c00",x"0000",x"0000",x"3a40",x"34db",x"3193",x"3743",x"36d4",x"3c00",x"0000",x"0000",x"3a18",x"34d9",x"3193",x"3c44",x"36d0",x"3c00",x"0000",x"0000",x"3a07",x"34db"),
(x"3193",x"3c37",x"36e4",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c41",x"36fb",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c44",x"36d0",x"3c00",x"0000",x"0000",x"3a07",x"34db"),
(x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d",x"3143",x"374d",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"39af",x"3160",x"3716",x"36fb",x"0000",x"0000",x"3c00",x"39ff",x"39ab"),
(x"3143",x"374d",x"36fb",x"3993",x"1c9b",x"39bd",x"355f",x"38c8",x"3141",x"3c25",x"36fb",x"396d",x"9af6",x"39e0",x"355f",x"3742",x"3193",x"3743",x"36d4",x"396e",x"1b2b",x"39df",x"3552",x"38ca"),
(x"3143",x"374d",x"36fb",x"3993",x"1c9b",x"39bd",x"355f",x"38c8",x"3193",x"3743",x"36d4",x"396e",x"1b2b",x"39df",x"3552",x"38ca",x"3160",x"3716",x"36fb",x"3988",x"33a7",x"3973",x"355d",x"38cf"),
(x"3193",x"370d",x"36e5",x"396c",x"347c",x"396f",x"3555",x"38d1",x"3193",x"36e5",x"36fb",x"3969",x"359e",x"392e",x"3559",x"38d6",x"3160",x"3716",x"36fb",x"3988",x"33a7",x"3973",x"355d",x"38cf"),
(x"394e",x"3c44",x"36d0",x"ba68",x"217a",x"b8c9",x"3a8e",x"34d4",x"394e",x"3c44",x"36fb",x"bbf4",x"2eb8",x"0000",x"3a8e",x"34e8",x"394d",x"3c42",x"36fb",x"bbfe",x"276c",x"a4f7",x"3a91",x"34e8"),
(x"394d",x"3709",x"36dd",x"bbff",x"a074",x"a60a",x"3b14",x"34d8",x"394d",x"36db",x"36fb",x"bbff",x"a3a0",x"a0d0",x"3b17",x"34da",x"394e",x"36aa",x"36d0",x"3b8d",x"a187",x"b543",x"3b19",x"34d4"),
(x"394d",x"3709",x"36dd",x"ba1a",x"3321",x"38da",x"3569",x"372e",x"3959",x"3709",x"36fb",x"ba1d",x"31d2",x"38f2",x"3572",x"372e",x"394d",x"36db",x"36fb",x"b9d1",x"35ef",x"389f",x"356f",x"3722"),
(x"394d",x"3c28",x"36d8",x"bbf1",x"15bc",x"afa2",x"3aab",x"34d9",x"394d",x"3761",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b0f",x"34d8",x"394e",x"3c44",x"36d0",x"ba68",x"217a",x"b8c9",x"3a8e",x"34d4"),
(x"3962",x"376a",x"36fb",x"b9b6",x"128d",x"3999",x"3575",x"3747",x"3959",x"3709",x"36fb",x"ba1d",x"31d2",x"38f2",x"3572",x"372e",x"394d",x"3761",x"36ca",x"ba14",x"1cd0",x"3932",x"3566",x"3744"),
(x"3961",x"3c28",x"36fb",x"b935",x"9d6d",x"3a12",x"3572",x"38c9",x"3962",x"376a",x"36fb",x"b9b6",x"128d",x"3999",x"3575",x"3747",x"394d",x"3c28",x"36d8",x"b9b2",x"9dbc",x"399d",x"3566",x"38c9"),
(x"3961",x"3c28",x"36fb",x"b935",x"9d6d",x"3a12",x"3572",x"38c9",x"394d",x"3c28",x"36d8",x"b9b2",x"9dbc",x"399d",x"3566",x"38c9",x"3958",x"3c37",x"36fb",x"b94f",x"b2e4",x"39ba",x"356f",x"38d0"),
(x"394d",x"3c37",x"36e5",x"b97e",x"b36f",x"3983",x"3567",x"38d0",x"394d",x"3c42",x"36fb",x"b958",x"b562",x"394e",x"356b",x"38d6",x"3958",x"3c37",x"36fb",x"b94f",x"b2e4",x"39ba",x"356f",x"38d0"),
(x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d",x"2edb",x"39cd",x"36fb",x"0000",x"0000",x"3c00",x"39eb",x"3a03",x"2ef7",x"397e",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"39f7"),
(x"2c34",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3b36",x"30cd",x"3a2c",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3a7a",x"30cd",x"2c34",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3b36",x"3420"),
(x"2fe5",x"39c1",x"36fb",x"bb7d",x"359e",x"0000",x"3b31",x"3a08",x"2fe5",x"39c1",x"36b4",x"bb3f",x"36c6",x"0000",x"3b31",x"3a10",x"3009",x"39cc",x"36fb",x"bb8f",x"3538",x"0000",x"3b34",x"3a08"),
(x"2ef7",x"397e",x"36fb",x"a439",x"3bff",x"91bc",x"3b77",x"3a39",x"2f02",x"397e",x"36b4",x"a44d",x"3bff",x"8e8d",x"3b6d",x"3a39",x"3025",x"397f",x"36fb",x"a44d",x"3bff",x"8cea",x"3b77",x"3a43"),
(x"2f19",x"39d7",x"36fb",x"36f3",x"bb34",x"0000",x"3b3f",x"3a08",x"2f19",x"39d7",x"36b4",x"3917",x"ba2b",x"2153",x"3b3f",x"3a10",x"2edb",x"39cd",x"36fb",x"3bbb",x"b413",x"26dc",x"3b42",x"3a08"),
(x"3009",x"39cc",x"36fb",x"bb8f",x"3538",x"0000",x"3b34",x"3a08",x"3009",x"39cc",x"36b4",x"bbef",x"3012",x"0000",x"3b34",x"3a10",x"3004",x"39d4",x"36fb",x"baa8",x"b870",x"0000",x"3b36",x"3a08"),
(x"3025",x"397f",x"36fb",x"bbcb",x"b335",x"0000",x"3b1f",x"3a08",x"3025",x"397f",x"36b4",x"bbcb",x"b335",x"0000",x"3b1f",x"3a10",x"2fda",x"39bb",x"36fb",x"bbd4",x"b28e",x"0000",x"3b2f",x"3a08"),
(x"2edb",x"39cd",x"36fb",x"3bbb",x"b413",x"26dc",x"3b42",x"3a08",x"2ee6",x"39cd",x"36b4",x"3bf0",x"2f65",x"2911",x"3b42",x"3a10",x"2f05",x"39c0",x"36fb",x"3bf5",x"2e12",x"2918",x"3b45",x"3a08"),
(x"3004",x"39d4",x"36fb",x"baa8",x"b870",x"0000",x"3b36",x"3a08",x"3004",x"39d4",x"36b4",x"b8fa",x"ba42",x"0000",x"3b36",x"3a10",x"2f99",x"39db",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a08"),
(x"2fda",x"39bb",x"36fb",x"bbd4",x"b28e",x"0000",x"3b2f",x"3a08",x"2fda",x"39bb",x"36b4",x"bbe8",x"b0e3",x"0000",x"3b2f",x"3a10",x"2fe5",x"39c1",x"36fb",x"bb7d",x"359e",x"0000",x"3b31",x"3a08"),
(x"2f05",x"39c0",x"36fb",x"3bf5",x"2e12",x"2918",x"3b45",x"3a08",x"2f10",x"39c0",x"36b4",x"3bfe",x"2231",x"291b",x"3b45",x"3a10",x"2ef7",x"397e",x"36fb",x"3bfd",x"a6cf",x"291b",x"3b57",x"3a08"),
(x"2f99",x"39db",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a08",x"2f99",x"39db",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a10",x"2f19",x"39d7",x"36fb",x"36f3",x"bb34",x"0000",x"3b3f",x"3a08"),
(x"2da5",x"3cbe",x"36fa",x"0000",x"8000",x"bc00",x"350f",x"3ab5",x"2a34",x"3cbe",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"3ab5",x"2da5",x"34c1",x"36fa",x"0000",x"8000",x"bc00",x"350f",x"38f4"),
(x"2a34",x"3cbe",x"36fa",x"baf4",x"0000",x"37e6",x"35a4",x"3a80",x"2af5",x"3cb6",x"3725",x"baf4",x"0000",x"37e6",x"35b0",x"3a7b",x"2a34",x"34c1",x"36fa",x"baf4",x"0000",x"37e6",x"35a4",x"38f4"),
(x"2d44",x"34e1",x"3725",x"0000",x"0000",x"3c00",x"358a",x"38f4",x"2af5",x"34e1",x"3725",x"0000",x"0000",x"3c00",x"3571",x"38f4",x"2d44",x"3cb6",x"3725",x"0000",x"0000",x"3c00",x"358a",x"3aad"),
(x"2d44",x"3cb6",x"3725",x"0000",x"3a66",x"38cc",x"3b15",x"3ba0",x"2af5",x"3cb6",x"3725",x"0000",x"3a66",x"38cc",x"3b06",x"3ba0",x"2da5",x"3cbe",x"36fa",x"0000",x"3a66",x"38cc",x"3b19",x"3ba8"),
(x"2a34",x"34c1",x"36fa",x"0000",x"ba66",x"38cc",x"3b02",x"3bb1",x"2af5",x"34e1",x"3725",x"0000",x"ba66",x"38cc",x"3b06",x"3bb9",x"2da5",x"34c1",x"36fa",x"0000",x"ba66",x"38cc",x"3b19",x"3bb1"),
(x"2da5",x"3cbe",x"36fa",x"3af4",x"0000",x"37e6",x"3597",x"3a7f",x"2da5",x"34c1",x"36fa",x"3af4",x"0000",x"37e6",x"3597",x"38f4",x"2d44",x"3cb6",x"3725",x"3af4",x"0000",x"37e6",x"358b",x"3a7c"),
(x"3a2c",x"3cc1",x"36fb",x"3c00",x"0000",x"0000",x"35f8",x"3a68",x"3a2c",x"3cc1",x"368e",x"3c00",x"0000",x"0000",x"360d",x"3a68",x"3a2c",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"360d",x"38f3"),
(x"2c34",x"3cc1",x"368e",x"bc00",x"8000",x"0000",x"383c",x"3508",x"2c34",x"3cc1",x"36fb",x"bc00",x"8000",x"0000",x"385a",x"3508",x"2c34",x"34b8",x"36fb",x"bc00",x"8000",x"0000",x"385a",x"1cef"),
(x"394e",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3af7",x"3838",x"394e",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3af7",x"3832",x"3193",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3a04",x"3832"),
(x"2c34",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"38eb",x"3bdb",x"2c34",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"38eb",x"3bf4",x"3a2c",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"39b1",x"3bf4"),
(x"3a2c",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"39b0",x"3bd3",x"3a2c",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"39b0",x"3bb9",x"2c34",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"38ea",x"3bb9"),
(x"3959",x"3709",x"36fb",x"0000",x"0000",x"3c00",x"3aa2",x"39aa",x"394e",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"39a2",x"394d",x"36db",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"39a6"),
(x"3959",x"3709",x"36fb",x"0000",x"0000",x"3c00",x"3aa2",x"39aa",x"3a2c",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"397d",x"394e",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"39a2"),
(x"3958",x"3c37",x"36fb",x"0000",x"0000",x"3c00",x"3aa1",x"3a69",x"394e",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"3a6d",x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93"),
(x"3958",x"3c37",x"36fb",x"0000",x"0000",x"3c00",x"3aa1",x"3a69",x"394d",x"3c42",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"3a6d",x"394e",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3aa0",x"3a6d"),
(x"3a2c",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"397d",x"3959",x"3709",x"36fb",x"0000",x"0000",x"3c00",x"3aa2",x"39aa",x"3962",x"376a",x"36fb",x"0000",x"0000",x"3c00",x"3aa3",x"39b1"),
(x"3961",x"3c28",x"36fb",x"0000",x"0000",x"3c00",x"3aa3",x"3a65",x"3958",x"3c37",x"36fb",x"0000",x"0000",x"3c00",x"3aa1",x"3a69",x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93"),
(x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93",x"3962",x"376a",x"36fb",x"0000",x"0000",x"3c00",x"3aa3",x"39b1",x"3961",x"3c28",x"36fb",x"0000",x"0000",x"3c00",x"3aa3",x"3a65"),
(x"316f",x"3c38",x"36fb",x"0000",x"0000",x"3c00",x"3a00",x"3a6a",x"3193",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"3a6d",x"3193",x"3c41",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"3a6c"),
(x"316f",x"3c38",x"36fb",x"0000",x"0000",x"3c00",x"3a00",x"3a6a",x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93",x"3193",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"3a6d"),
(x"2edb",x"39cd",x"36fb",x"0000",x"0000",x"3c00",x"39eb",x"3a03",x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d",x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93"),
(x"2f19",x"39d7",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"3a04",x"2edb",x"39cd",x"36fb",x"0000",x"0000",x"3c00",x"39eb",x"3a03",x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"3143",x"374d",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"39af",x"3025",x"397f",x"36fb",x"0000",x"0000",x"3c00",x"39f3",x"39f7"),
(x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93",x"316f",x"3c38",x"36fb",x"0000",x"0000",x"3c00",x"3a00",x"3a6a",x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"2f19",x"39d7",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"3a04",x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"2f99",x"39db",x"36fb",x"0000",x"0000",x"3c00",x"39ef",x"3a05",x"2f19",x"39d7",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"3a04"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"3004",x"39d4",x"36fb",x"868d",x"0000",x"3c00",x"39f1",x"3a04",x"2f99",x"39db",x"36fb",x"0000",x"0000",x"3c00",x"39ef",x"3a05"),
(x"3009",x"39cc",x"36fb",x"0000",x"0000",x"3c00",x"39f1",x"3a03",x"2fda",x"39bb",x"36fb",x"0000",x"0000",x"3c00",x"39f0",x"3a00",x"2fe5",x"39c1",x"36fb",x"0000",x"0000",x"3c00",x"39f1",x"3a01"),
(x"3009",x"39cc",x"36fb",x"0000",x"0000",x"3c00",x"39f1",x"3a03",x"3025",x"397f",x"36fb",x"0000",x"0000",x"3c00",x"39f3",x"39f7",x"2fda",x"39bb",x"36fb",x"0000",x"0000",x"3c00",x"39f0",x"3a00"),
(x"3141",x"3c25",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"3a64",x"3025",x"397f",x"36fb",x"0000",x"0000",x"3c00",x"39f3",x"39f7",x"3009",x"39cc",x"36fb",x"0000",x"0000",x"3c00",x"39f1",x"3a03"),
(x"3a2c",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"397d",x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d",x"3193",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"39a2"),
(x"3193",x"3c44",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"3a6d",x"2c34",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"3a93",x"3a2c",x"3cc1",x"36fb",x"0000",x"0000",x"3c00",x"3ac3",x"3a93"),
(x"3193",x"3c44",x"36d0",x"0000",x"0000",x"3c00",x"31b2",x"3bf9",x"394e",x"3c44",x"36d0",x"0000",x"0000",x"3c00",x"3468",x"3bf9",x"394e",x"36aa",x"36d0",x"0000",x"0000",x"3c00",x"3468",x"3adb"),
(x"3193",x"36aa",x"36d0",x"3c00",x"0000",x"0000",x"3a40",x"34db",x"3193",x"36aa",x"36fb",x"3c00",x"0000",x"0000",x"3a40",x"34c6",x"3193",x"36e5",x"36fb",x"3c00",x"0000",x"0000",x"3a31",x"34c6"),
(x"3193",x"370d",x"36e5",x"3c00",x"0000",x"0000",x"3a26",x"34d1",x"3193",x"3743",x"36d4",x"3c00",x"0000",x"0000",x"3a18",x"34d9",x"3193",x"36aa",x"36d0",x"3c00",x"0000",x"0000",x"3a40",x"34db"),
(x"3193",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3af4",x"35b9",x"3193",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3af4",x"35cd",x"394e",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3b7d",x"35cd"),
(x"316f",x"3c38",x"36fb",x"39bc",x"b304",x"394a",x"355b",x"372f",x"3193",x"3c37",x"36e4",x"3a1e",x"b322",x"38d5",x"3554",x"3730",x"3193",x"3c28",x"36d7",x"394c",x"a074",x"39fd",x"3552",x"373f"),
(x"3193",x"36aa",x"36fb",x"0000",x"0000",x"3c00",x"3a01",x"39a2",x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d",x"3160",x"3716",x"36fb",x"0000",x"0000",x"3c00",x"39ff",x"39ab"),
(x"3193",x"3743",x"36d4",x"3c00",x"0000",x"0000",x"3a18",x"34d9",x"3193",x"3c28",x"36d7",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c44",x"36d0",x"3c00",x"0000",x"0000",x"3a07",x"34db"),
(x"3193",x"3c41",x"36fb",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c44",x"36fb",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c44",x"36d0",x"3c00",x"0000",x"0000",x"3a07",x"34db"),
(x"3193",x"3c44",x"36d0",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c28",x"36d7",x"3c00",x"0000",x"0000",x"3a07",x"34db",x"3193",x"3c37",x"36e4",x"3c00",x"0000",x"0000",x"3a07",x"34db"),
(x"3141",x"3c25",x"36fb",x"396d",x"9af6",x"39e0",x"355f",x"3742",x"3193",x"3c28",x"36d7",x"394c",x"a074",x"39fd",x"3552",x"373f",x"3193",x"3743",x"36d4",x"396e",x"1b2b",x"39df",x"3552",x"38ca"),
(x"3193",x"3743",x"36d4",x"396e",x"1b2b",x"39df",x"3552",x"38ca",x"3193",x"370d",x"36e5",x"396c",x"347c",x"396f",x"3555",x"38d1",x"3160",x"3716",x"36fb",x"3988",x"33a7",x"3973",x"355d",x"38cf"),
(x"394d",x"3c37",x"36e5",x"bbfe",x"2111",x"a779",x"3a9c",x"34de",x"394d",x"3c28",x"36d8",x"bbf1",x"15bc",x"afa2",x"3aab",x"34d9",x"394e",x"3c44",x"36d0",x"ba68",x"217a",x"b8c9",x"3a8e",x"34d4"),
(x"394e",x"3c44",x"36d0",x"ba68",x"217a",x"b8c9",x"3a8e",x"34d4",x"394d",x"3c42",x"36fb",x"bbfe",x"276c",x"a4f7",x"3a91",x"34e8",x"394d",x"3c37",x"36e5",x"bbfe",x"2111",x"a779",x"3a9c",x"34de"),
(x"394d",x"36db",x"36fb",x"bbff",x"a3a0",x"a0d0",x"3b17",x"34da",x"394e",x"36aa",x"36fb",x"bbff",x"a5e9",x"0000",x"3b19",x"34d8",x"394e",x"36aa",x"36d0",x"3b8d",x"a187",x"b543",x"3b19",x"34d4"),
(x"394e",x"36aa",x"36d0",x"3b8d",x"a187",x"b543",x"3b19",x"34d4",x"394d",x"3761",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b0f",x"34d8",x"394d",x"3709",x"36dd",x"bbff",x"a074",x"a60a",x"3b14",x"34d8"),
(x"394d",x"3761",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b0f",x"34d8",x"394e",x"36aa",x"36d0",x"3b8d",x"a187",x"b543",x"3b19",x"34d4",x"394e",x"3c44",x"36d0",x"ba68",x"217a",x"b8c9",x"3a8e",x"34d4"),
(x"3959",x"3709",x"36fb",x"ba1d",x"31d2",x"38f2",x"3572",x"372e",x"394d",x"3709",x"36dd",x"ba1a",x"3321",x"38da",x"3569",x"372e",x"394d",x"3761",x"36ca",x"ba14",x"1cd0",x"3932",x"3566",x"3744"),
(x"3962",x"376a",x"36fb",x"b9b6",x"128d",x"3999",x"3575",x"3747",x"394d",x"3761",x"36ca",x"ba14",x"1cd0",x"3932",x"3566",x"3744",x"394d",x"3c28",x"36d8",x"b9b2",x"9dbc",x"399d",x"3566",x"38c9"),
(x"394d",x"3c28",x"36d8",x"b9b2",x"9dbc",x"399d",x"3566",x"38c9",x"394d",x"3c37",x"36e5",x"b97e",x"b36f",x"3983",x"3567",x"38d0",x"3958",x"3c37",x"36fb",x"b94f",x"b2e4",x"39ba",x"356f",x"38d0"),
(x"2ef7",x"397e",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"39f7",x"3143",x"374d",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"39af",x"2c34",x"34b8",x"36fb",x"0000",x"0000",x"3c00",x"39de",x"397d"),
(x"2ef7",x"397e",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"39f7",x"3025",x"397f",x"36fb",x"0000",x"0000",x"3c00",x"39f3",x"39f7",x"3143",x"374d",x"36fb",x"0000",x"0000",x"3c00",x"39fe",x"39af"),
(x"2edb",x"39cd",x"36fb",x"0000",x"0000",x"3c00",x"39eb",x"3a03",x"2f05",x"39c0",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"3a01",x"2ef7",x"397e",x"36fb",x"0000",x"0000",x"3c00",x"39ec",x"39f7"),
(x"3a2c",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3a7a",x"30cd",x"3a2c",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3a7a",x"3420",x"2c34",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3b36",x"3420"),
(x"2fe5",x"39c1",x"36b4",x"bb3f",x"36c6",x"0000",x"3b31",x"3a10",x"3009",x"39cc",x"36b4",x"bbef",x"3012",x"0000",x"3b34",x"3a10",x"3009",x"39cc",x"36fb",x"bb8f",x"3538",x"0000",x"3b34",x"3a08"),
(x"2f02",x"397e",x"36b4",x"a44d",x"3bff",x"8e8d",x"3b6d",x"3a39",x"3025",x"397f",x"36b4",x"a460",x"3bff",x"0000",x"3b6d",x"3a43",x"3025",x"397f",x"36fb",x"a44d",x"3bff",x"8cea",x"3b77",x"3a43"),
(x"2f19",x"39d7",x"36b4",x"3917",x"ba2b",x"2153",x"3b3f",x"3a10",x"2ee6",x"39cd",x"36b4",x"3bf0",x"2f65",x"2911",x"3b42",x"3a10",x"2edb",x"39cd",x"36fb",x"3bbb",x"b413",x"26dc",x"3b42",x"3a08"),
(x"3009",x"39cc",x"36b4",x"bbef",x"3012",x"0000",x"3b34",x"3a10",x"3004",x"39d4",x"36b4",x"b8fa",x"ba42",x"0000",x"3b36",x"3a10",x"3004",x"39d4",x"36fb",x"baa8",x"b870",x"0000",x"3b36",x"3a08"),
(x"3025",x"397f",x"36b4",x"bbcb",x"b335",x"0000",x"3b1f",x"3a10",x"2fda",x"39bb",x"36b4",x"bbe8",x"b0e3",x"0000",x"3b2f",x"3a10",x"2fda",x"39bb",x"36fb",x"bbd4",x"b28e",x"0000",x"3b2f",x"3a08"),
(x"2ee6",x"39cd",x"36b4",x"3bf0",x"2f65",x"2911",x"3b42",x"3a10",x"2f10",x"39c0",x"36b4",x"3bfe",x"2231",x"291b",x"3b45",x"3a10",x"2f05",x"39c0",x"36fb",x"3bf5",x"2e12",x"2918",x"3b45",x"3a08"),
(x"3004",x"39d4",x"36b4",x"b8fa",x"ba42",x"0000",x"3b36",x"3a10",x"2f99",x"39db",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a10",x"2f99",x"39db",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a08"),
(x"2fda",x"39bb",x"36b4",x"bbe8",x"b0e3",x"0000",x"3b2f",x"3a10",x"2fe5",x"39c1",x"36b4",x"bb3f",x"36c6",x"0000",x"3b31",x"3a10",x"2fe5",x"39c1",x"36fb",x"bb7d",x"359e",x"0000",x"3b31",x"3a08"),
(x"2f10",x"39c0",x"36b4",x"3bfe",x"2231",x"291b",x"3b45",x"3a10",x"2f02",x"397e",x"36b4",x"3bfd",x"a6cf",x"291b",x"3b57",x"3a10",x"2ef7",x"397e",x"36fb",x"3bfd",x"a6cf",x"291b",x"3b57",x"3a08"),
(x"2f99",x"39db",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a10",x"2f19",x"39d7",x"36b4",x"3917",x"ba2b",x"2153",x"3b3f",x"3a10",x"2f19",x"39d7",x"36fb",x"36f3",x"bb34",x"0000",x"3b3f",x"3a08"),
(x"2a34",x"3cbe",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"3ab5",x"2a34",x"34c1",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"38f4",x"2da5",x"34c1",x"36fa",x"0000",x"8000",x"bc00",x"350f",x"38f4"),
(x"2af5",x"3cb6",x"3725",x"baf4",x"0000",x"37e6",x"35b0",x"3a7b",x"2af5",x"34e1",x"3725",x"baf4",x"0000",x"37e6",x"35b0",x"38f7",x"2a34",x"34c1",x"36fa",x"baf4",x"0000",x"37e6",x"35a4",x"38f4"),
(x"2af5",x"34e1",x"3725",x"0000",x"0000",x"3c00",x"3571",x"38f4",x"2af5",x"3cb6",x"3725",x"0000",x"0000",x"3c00",x"3571",x"3aad",x"2d44",x"3cb6",x"3725",x"0000",x"0000",x"3c00",x"358a",x"3aad"),
(x"2af5",x"3cb6",x"3725",x"0000",x"3a66",x"38cc",x"3b06",x"3ba0",x"2a34",x"3cbe",x"36fa",x"0000",x"3a66",x"38cc",x"3b02",x"3ba8",x"2da5",x"3cbe",x"36fa",x"0000",x"3a66",x"38cc",x"3b19",x"3ba8"),
(x"2af5",x"34e1",x"3725",x"0000",x"ba66",x"38cc",x"3b06",x"3bb9",x"2d44",x"34e1",x"3725",x"0000",x"ba66",x"38cc",x"3b15",x"3bb9",x"2da5",x"34c1",x"36fa",x"0000",x"ba66",x"38cc",x"3b19",x"3bb1"),
(x"2da5",x"34c1",x"36fa",x"3af4",x"0000",x"37e6",x"3597",x"38f4",x"2d44",x"34e1",x"3725",x"3af4",x"0000",x"37e6",x"358a",x"38f8",x"2d44",x"3cb6",x"3725",x"3af4",x"0000",x"37e6",x"358b",x"3a7c"),
(x"2f10",x"39c0",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"350c",x"2fe5",x"39c1",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"351a",x"2fda",x"39bb",x"36b4",x"0000",x"0000",x"3c00",x"3a96",x"3519"),
(x"303e",x"39c2",x"3718",x"3bb8",x"b22d",x"31b0",x"3934",x"3040",x"304f",x"39c2",x"36eb",x"3ba3",x"b452",x"2fdf",x"393f",x"3031",x"3033",x"39b8",x"3715",x"3bf4",x"2da3",x"2b3e",x"3933",x"302a"),
(x"303e",x"39c2",x"3718",x"3bb8",x"b22d",x"31b0",x"3934",x"3040",x"3048",x"39d2",x"3715",x"3bda",x"2e4f",x"312f",x"3937",x"305f",x"304f",x"39c2",x"36eb",x"3ba3",x"b452",x"2fdf",x"393f",x"3031"),
(x"3048",x"39d2",x"3715",x"3bda",x"2e4f",x"312f",x"3937",x"305f",x"3027",x"39e1",x"3714",x"3a0a",x"3915",x"3126",x"393a",x"3083",x"3054",x"39d2",x"36eb",x"3b7a",x"3531",x"30a8",x"3942",x"3052"),
(x"3027",x"39e1",x"3714",x"3a0a",x"3915",x"3126",x"393a",x"3083",x"2fca",x"39e9",x"3714",x"3235",x"3bc0",x"30e0",x"393b",x"30aa",x"302b",x"39e5",x"36eb",x"38c7",x"3a49",x"310b",x"3944",x"307f"),
(x"2fca",x"39e9",x"3714",x"3235",x"3bc0",x"30e0",x"393b",x"30aa",x"2ef2",x"39e6",x"3714",x"b35f",x"3baf",x"30fd",x"393c",x"30e4",x"2fcc",x"39ec",x"36eb",x"23ae",x"3bec",x"306c",x"3945",x"30a6"),
(x"2ef2",x"39e6",x"3714",x"b35f",x"3baf",x"30fd",x"393c",x"30e4",x"2e86",x"39db",x"3715",x"ba37",x"38de",x"311d",x"393b",x"310a",x"2ed8",x"39e9",x"36eb",x"b6e0",x"3b1c",x"3118",x"3946",x"30e8"),
(x"2e86",x"39db",x"3715",x"ba37",x"38de",x"311d",x"393b",x"310a",x"2e63",x"39cc",x"3715",x"bbf2",x"2495",x"2f43",x"393a",x"312b",x"2e6e",x"39db",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3945",x"3110"),
(x"2e80",x"39be",x"3715",x"bb87",x"b537",x"2d81",x"3938",x"3149",x"2e6b",x"39be",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3943",x"3150",x"2e63",x"39cc",x"3715",x"bbf2",x"2495",x"2f43",x"393a",x"312b"),
(x"2e96",x"39b5",x"3717",x"bbff",x"2481",x"2487",x"3937",x"315d",x"2e93",x"39b4",x"36eb",x"bbfd",x"212b",x"29e6",x"3942",x"3166",x"2e80",x"39be",x"3715",x"bb87",x"b537",x"2d81",x"3938",x"3149"),
(x"2e34",x"397f",x"36eb",x"bb76",x"3593",x"2dee",x"393d",x"31e3",x"2e6c",x"3981",x"36eb",x"bb9b",x"34d2",x"2ca7",x"393d",x"31d3",x"2e3f",x"397d",x"3714",x"bb74",x"35a7",x"2d5e",x"3933",x"31dc"),
(x"2f2c",x"39c2",x"36eb",x"3b82",x"350f",x"3071",x"38af",x"31f1",x"2f22",x"39b7",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38af",x"3208",x"2f16",x"39c0",x"3716",x"3ba5",x"3473",x"2e24",x"38ba",x"31f3"),
(x"2f22",x"39b7",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38af",x"3208",x"2f2a",x"3983",x"36eb",x"3a79",x"3840",x"3401",x"38b0",x"3278",x"2f13",x"39b7",x"3718",x"3bf1",x"95bc",x"2fb6",x"38bb",x"3207"),
(x"3072",x"3969",x"3715",x"33c8",x"bbc2",x"235f",x"3921",x"2f0d",x"306e",x"397f",x"3715",x"3bb4",x"33e8",x"2ed7",x"3926",x"2f62",x"3079",x"3969",x"36eb",x"3409",x"bbbc",x"27db",x"392b",x"2ee7"),
(x"2e32",x"396a",x"3714",x"af03",x"bbf3",x"23ef",x"3930",x"3204",x"2e24",x"3969",x"36eb",x"b6d0",x"bb39",x"2ab1",x"393a",x"3210",x"2e3f",x"397d",x"3714",x"bb74",x"35a7",x"2d5e",x"3933",x"31dc"),
(x"2fd9",x"39b7",x"3716",x"bbce",x"b2bb",x"2b41",x"38bc",x"313e",x"2fc8",x"39b8",x"36eb",x"bbd3",x"b208",x"2da6",x"38b1",x"313c",x"2fd7",x"39bf",x"3715",x"bb88",x"3531",x"2dc2",x"38bb",x"314f"),
(x"2fc7",x"39c0",x"36ee",x"bb70",x"358e",x"2fc0",x"38b1",x"314f",x"2ffa",x"39c8",x"36ee",x"bb20",x"3725",x"2d51",x"38b2",x"3164",x"2fd7",x"39bf",x"3715",x"bb88",x"3531",x"2dc2",x"38bb",x"314f"),
(x"2ffa",x"39c8",x"36ee",x"bb20",x"3725",x"2d51",x"38b2",x"3164",x"2fff",x"39d0",x"36ee",x"bb1d",x"b747",x"2911",x"38b1",x"3176",x"3005",x"39ca",x"3717",x"bbd6",x"323b",x"2a8a",x"38bc",x"3169"),
(x"2f3e",x"39d9",x"36ee",x"3123",x"bbe4",x"a874",x"38b1",x"31b1",x"2ef6",x"39d0",x"36ee",x"3a41",x"b8fc",x"243f",x"38b0",x"31cc",x"2f3a",x"39d8",x"3715",x"3670",x"bb52",x"9df0",x"38ba",x"31b4"),
(x"2fc8",x"39b8",x"36eb",x"bbd3",x"b208",x"2da6",x"38b1",x"313c",x"2fd9",x"39b7",x"3716",x"bbce",x"b2bb",x"2b41",x"38bc",x"313e",x"3016",x"3985",x"36eb",x"bbe6",x"2cac",x"3077",x"38b3",x"30cc"),
(x"2e77",x"3981",x"3717",x"a984",x"a0c2",x"3bfd",x"3963",x"31ac",x"2e32",x"396a",x"3714",x"a73e",x"ad9b",x"3bf7",x"3961",x"318d",x"2e3f",x"397d",x"3714",x"b3e6",x"2587",x"3bc0",x"3961",x"31a7"),
(x"3056",x"3980",x"3718",x"26a1",x"97c8",x"3bff",x"3977",x"31ab",x"306e",x"397f",x"3715",x"33f4",x"1d38",x"3bbf",x"3979",x"31aa",x"3072",x"3969",x"3715",x"2081",x"ad9e",x"3bf8",x"3979",x"318d"),
(x"303e",x"39c2",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3975",x"3203",x"3033",x"39b8",x"3715",x"21a1",x"23fc",x"3bff",x"3974",x"31f5",x"2fd7",x"39bf",x"3715",x"a8d3",x"a80e",x"3bfd",x"396f",x"31ff"),
(x"3048",x"39d2",x"3715",x"1e59",x"2bec",x"3bfc",x"3976",x"3218",x"303e",x"39c2",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3975",x"3203",x"3005",x"39ca",x"3717",x"a511",x"281b",x"3bfe",x"3971",x"320c"),
(x"3027",x"39e1",x"3714",x"a63f",x"27c1",x"3bfe",x"3973",x"322b",x"3048",x"39d2",x"3715",x"1e59",x"2bec",x"3bfc",x"3976",x"3218",x"2fff",x"39d2",x"3716",x"a52b",x"2c98",x"3bfa",x"3971",x"3218"),
(x"2fca",x"39e9",x"3714",x"217a",x"a0ea",x"3bff",x"396f",x"3236",x"3027",x"39e1",x"3714",x"a63f",x"27c1",x"3bfe",x"3973",x"322b",x"2fc2",x"39d7",x"3713",x"991e",x"9cd0",x"3c00",x"396f",x"321e"),
(x"2ef2",x"39e6",x"3714",x"9dbc",x"247a",x"3bff",x"3967",x"3232",x"2fca",x"39e9",x"3714",x"217a",x"a0ea",x"3bff",x"396f",x"3236",x"2f3a",x"39d8",x"3715",x"1c81",x"1953",x"3c00",x"396a",x"3220"),
(x"2e86",x"39db",x"3715",x"2793",x"184d",x"3bff",x"3963",x"3223",x"2ef2",x"39e6",x"3714",x"9dbc",x"247a",x"3bff",x"3967",x"3232",x"2ef1",x"39d0",x"3714",x"1da1",x"252b",x"3bff",x"3967",x"3215"),
(x"2e86",x"39db",x"3715",x"2793",x"184d",x"3bff",x"3963",x"3223",x"2ef1",x"39d0",x"3714",x"1da1",x"252b",x"3bff",x"3967",x"3215",x"2e63",x"39cc",x"3715",x"1818",x"26bb",x"3bff",x"3962",x"320f"),
(x"2e63",x"39cc",x"3715",x"1818",x"26bb",x"3bff",x"3962",x"320f",x"2eed",x"39c9",x"3716",x"a338",x"267a",x"3bff",x"3967",x"320c",x"2e80",x"39be",x"3715",x"a64c",x"29dc",x"3bfd",x"3963",x"31fd"),
(x"2e96",x"39b5",x"3717",x"a7d5",x"236c",x"3bfe",x"3964",x"31f0",x"2e80",x"39be",x"3715",x"a64c",x"29dc",x"3bfd",x"3963",x"31fd",x"2f13",x"39b7",x"3718",x"a793",x"2439",x"3bfe",x"3968",x"31f3"),
(x"2f0c",x"397d",x"3718",x"a3ae",x"ac2d",x"3bfb",x"3968",x"31a7",x"2e77",x"3981",x"3717",x"a984",x"a0c2",x"3bfd",x"3963",x"31ac",x"2f13",x"39b7",x"3718",x"a793",x"2439",x"3bfe",x"3968",x"31f3"),
(x"2ef6",x"39d0",x"36ee",x"3a41",x"b8fc",x"243f",x"38b0",x"31cc",x"2ef0",x"39c9",x"36ee",x"3b71",x"35c6",x"2c00",x"38b0",x"31db",x"2ef1",x"39d0",x"3714",x"3b3d",x"b6cc",x"26f6",x"38ba",x"31ce"),
(x"3056",x"3980",x"3718",x"3ba4",x"33dc",x"313d",x"3926",x"2f7d",x"3033",x"39b8",x"3715",x"3bf4",x"2da3",x"2b3e",x"3933",x"302a",x"3065",x"3981",x"36eb",x"3baa",x"3479",x"2b93",x"3930",x"2f54"),
(x"3077",x"3981",x"36eb",x"3bc6",x"328d",x"2f71",x"3930",x"2f41",x"306e",x"397f",x"3715",x"3bb4",x"33e8",x"2ed7",x"3926",x"2f62",x"3065",x"3981",x"36eb",x"3baa",x"3479",x"2b93",x"3930",x"2f54"),
(x"2f0c",x"397d",x"3718",x"a3ae",x"ac2d",x"3bfb",x"3968",x"31a7",x"2e32",x"396a",x"3714",x"a73e",x"ad9b",x"3bf7",x"3961",x"318d",x"2e77",x"3981",x"3717",x"a984",x"a0c2",x"3bfd",x"3963",x"31ac"),
(x"2e32",x"396a",x"3714",x"a73e",x"ad9b",x"3bf7",x"3961",x"318d",x"2f0c",x"397d",x"3718",x"a3ae",x"ac2d",x"3bfb",x"3968",x"31a7",x"3072",x"3969",x"3715",x"2081",x"ad9e",x"3bf8",x"3979",x"318d"),
(x"301e",x"397e",x"3718",x"224c",x"a379",x"3bff",x"3973",x"31a9",x"3056",x"3980",x"3718",x"26a1",x"97c8",x"3bff",x"3977",x"31ab",x"3072",x"3969",x"3715",x"2081",x"ad9e",x"3bf8",x"3979",x"318d"),
(x"2fff",x"39d2",x"3716",x"baa5",x"b86c",x"2baa",x"38bb",x"317d",x"2fff",x"39d0",x"36ee",x"bb1d",x"b747",x"2911",x"38b1",x"3176",x"2fc2",x"39d7",x"3713",x"b46c",x"bbaf",x"a5f6",x"38ba",x"318f"),
(x"2e96",x"39b5",x"3717",x"bbff",x"2481",x"2487",x"3937",x"315d",x"2e77",x"3981",x"3717",x"bbe8",x"30a2",x"2973",x"3932",x"31ca",x"2e93",x"39b4",x"36eb",x"bbfd",x"212b",x"29e6",x"3942",x"3166"),
(x"2fc4",x"39d8",x"36ee",x"b52c",x"bb8d",x"ac0b",x"38b1",x"318d",x"2f3e",x"39d9",x"36ee",x"3123",x"bbe4",x"a874",x"38b1",x"31b1",x"2fc2",x"39d7",x"3713",x"b46c",x"bbaf",x"a5f6",x"38ba",x"318f"),
(x"2f0c",x"397d",x"3718",x"3a6d",x"3838",x"3468",x"38ba",x"3073",x"2f2a",x"3983",x"36eb",x"3a79",x"3840",x"3401",x"38af",x"3089",x"301e",x"397e",x"3718",x"b98b",x"396b",x"33db",x"38bf",x"30c2"),
(x"2e24",x"3969",x"36eb",x"b6d0",x"bb39",x"2ab1",x"393a",x"3210",x"2e32",x"396a",x"3714",x"af03",x"bbf3",x"23ef",x"3930",x"3204",x"3079",x"3969",x"36eb",x"3409",x"bbbc",x"27db",x"392b",x"32c5"),
(x"2eed",x"39c9",x"3716",x"3ba8",x"349f",x"2474",x"38ba",x"31dd",x"2ef0",x"39c9",x"36ee",x"3b71",x"35c6",x"2c00",x"38b0",x"31db",x"2f16",x"39c0",x"3716",x"3ba5",x"3473",x"2e24",x"38ba",x"31f3"),
(x"3007",x"3b85",x"3715",x"ad56",x"20d0",x"3bf8",x"3980",x"3980",x"2f10",x"3b90",x"370e",x"afd2",x"2717",x"3bef",x"396f",x"3984",x"2fbb",x"3ba1",x"3716",x"b0f9",x"a8b2",x"3be5",x"3979",x"398f"),
(x"3007",x"3b85",x"3715",x"3bc5",x"2b9a",x"3358",x"396e",x"3078",x"2fbb",x"3ba1",x"3716",x"3add",x"375a",x"334d",x"396e",x"3097",x"301b",x"3b86",x"36eb",x"3b99",x"3315",x"330d",x"3973",x"3076"),
(x"301b",x"3b03",x"3713",x"291b",x"2b55",x"3bfb",x"3988",x"3936",x"2fb0",x"3b06",x"3714",x"2c39",x"29a5",x"3bf9",x"397f",x"3937",x"3001",x"3b16",x"3712",x"2a69",x"287e",x"3bfc",x"3984",x"3940"),
(x"303e",x"3b06",x"3712",x"2a73",x"2a97",x"3bfa",x"398d",x"3938",x"3017",x"3b1a",x"3711",x"2994",x"2977",x"3bfc",x"3987",x"3943",x"304c",x"3b12",x"3711",x"2481",x"2546",x"3bff",x"398e",x"393e"),
(x"3017",x"3b1a",x"3711",x"2994",x"2977",x"3bfc",x"3987",x"3943",x"303e",x"3b06",x"3712",x"2a73",x"2a97",x"3bfa",x"398d",x"3938",x"3001",x"3b16",x"3712",x"2a69",x"287e",x"3bfc",x"3984",x"3940"),
(x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d",x"2ff2",x"3afd",x"3718",x"2e36",x"a153",x"3bf6",x"3984",x"3932",x"302f",x"3afb",x"3711",x"2fec",x"ac2c",x"3beb",x"398b",x"3931"),
(x"3040",x"3acf",x"370f",x"1df0",x"a631",x"3bff",x"398f",x"3918",x"301b",x"3acc",x"3713",x"2e9a",x"3366",x"3bbd",x"398a",x"3915",x"2ff4",x"3adb",x"370e",x"a6d5",x"25c2",x"3bfe",x"3985",x"391e"),
(x"2ff4",x"3adb",x"370e",x"a6d5",x"25c2",x"3bfe",x"3985",x"391e",x"3013",x"3ae4",x"3713",x"2538",x"ac79",x"3bfa",x"3988",x"3923",x"3040",x"3acf",x"370f",x"1df0",x"a631",x"3bff",x"398f",x"3918"),
(x"305c",x"3ad8",x"370f",x"2cd8",x"a71d",x"3bf9",x"3993",x"391e",x"3013",x"3ae4",x"3713",x"2538",x"ac79",x"3bfa",x"3988",x"3923",x"3058",x"3aeb",x"370f",x"2ec5",x"1a24",x"3bf4",x"3991",x"3928"),
(x"302f",x"3afb",x"3711",x"2fec",x"ac2c",x"3beb",x"398b",x"3931",x"3014",x"3ae7",x"3713",x"27e9",x"2849",x"3bfd",x"3988",x"3926",x"3000",x"3aec",x"3710",x"2c5b",x"b0a5",x"3be5",x"3985",x"3928"),
(x"2fd7",x"3a8d",x"3712",x"2f67",x"a981",x"3bf0",x"3983",x"38f2",x"2f48",x"3a8d",x"3715",x"26c2",x"ac65",x"3bfa",x"3979",x"38f2",x"2f7f",x"3a9c",x"3717",x"2ff2",x"aa7d",x"3bed",x"397d",x"38fa"),
(x"3044",x"3a9a",x"3714",x"9553",x"ab62",x"3bfc",x"398e",x"38f9",x"302b",x"3aae",x"3716",x"2cd8",x"a7e2",x"3bf9",x"398b",x"3905",x"3050",x"3aa2",x"3712",x"3163",x"a338",x"3be2",x"3990",x"38fe"),
(x"302b",x"3aae",x"3716",x"2cd8",x"a7e2",x"3bf9",x"398b",x"3905",x"3044",x"3a9a",x"3714",x"9553",x"ab62",x"3bfc",x"398e",x"38f9",x"300a",x"3aad",x"3716",x"a818",x"ad04",x"3bf8",x"3986",x"3904"),
(x"3000",x"3a94",x"3711",x"a40b",x"ad5c",x"3bf8",x"3985",x"38f6",x"2fd3",x"3aa6",x"3714",x"24fd",x"ada9",x"3bf7",x"3982",x"3900",x"300a",x"3aad",x"3716",x"a818",x"ad04",x"3bf8",x"3986",x"3904"),
(x"2fa9",x"3aa0",x"3714",x"3036",x"a73e",x"3bed",x"397f",x"38fc",x"3000",x"3a94",x"3711",x"a40b",x"ad5c",x"3bf8",x"3985",x"38f6",x"2fe3",x"3a91",x"3711",x"327d",x"175f",x"3bd5",x"3983",x"38f4"),
(x"302e",x"3a60",x"3711",x"3115",x"27d5",x"3be4",x"398c",x"38d9",x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"2fe6",x"3a82",x"3712",x"3146",x"2c91",x"3bde",x"3984",x"38ec"),
(x"2ef4",x"3a6b",x"3719",x"23bb",x"27c8",x"3bfe",x"3974",x"38de",x"2f3d",x"3a6b",x"3718",x"a138",x"ae95",x"3bf4",x"3979",x"38de",x"2ef3",x"3a69",x"3719",x"290e",x"af00",x"3bf2",x"3974",x"38dd"),
(x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"2f4b",x"3a60",x"3715",x"a8bf",x"afdb",x"3bef",x"397a",x"38d8",x"2f3d",x"3a6b",x"3718",x"a138",x"ae95",x"3bf4",x"3979",x"38de"),
(x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"2f3d",x"3a6b",x"3718",x"a138",x"ae95",x"3bf4",x"3979",x"38de",x"2f49",x"3a6d",x"3718",x"ab4f",x"2525",x"3bfc",x"3979",x"38df"),
(x"2f1d",x"3a89",x"3717",x"ad2d",x"2ecb",x"3bed",x"3976",x"38ef",x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2ede",x"3a7e",x"3718",x"acf2",x"18ea",x"3bf9",x"3972",x"38e9"),
(x"2ede",x"3a7e",x"3718",x"acf2",x"18ea",x"3bf9",x"3972",x"38e9",x"2ed4",x"3a86",x"3712",x"b59c",x"336a",x"3b42",x"3971",x"38ee",x"2f1d",x"3a89",x"3717",x"ad2d",x"2ecb",x"3bed",x"3976",x"38ef"),
(x"2fe6",x"3a82",x"3712",x"3146",x"2c91",x"3bde",x"3984",x"38ec",x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2f3a",x"3a8a",x"3716",x"3009",x"2da6",x"3be7",x"3978",x"38f0"),
(x"2f48",x"3a8d",x"3715",x"26c2",x"ac65",x"3bfa",x"3979",x"38f2",x"2fd7",x"3a8d",x"3712",x"2f67",x"a981",x"3bf0",x"3983",x"38f2",x"2f3a",x"3a8a",x"3716",x"3009",x"2da6",x"3be7",x"3978",x"38f0"),
(x"2f5a",x"3a9f",x"3717",x"17c8",x"9f93",x"3c00",x"397a",x"38fc",x"2f48",x"3a8d",x"3715",x"26c2",x"ac65",x"3bfa",x"3979",x"38f2",x"2f3c",x"3a92",x"3714",x"257a",x"ae8a",x"3bf4",x"3978",x"38f5"),
(x"2ece",x"3ab8",x"3714",x"adba",x"2266",x"3bf7",x"3971",x"390a",x"2f11",x"3aa9",x"3715",x"251e",x"2d06",x"3bf9",x"3975",x"3901",x"2e9f",x"3ab2",x"3714",x"975f",x"2c2c",x"3bfb",x"396e",x"3906"),
(x"2ec2",x"3ace",x"3715",x"b468",x"247a",x"3bb0",x"3971",x"3916",x"2ece",x"3ab8",x"3714",x"adba",x"2266",x"3bf7",x"3971",x"390a",x"2e7c",x"3acb",x"3712",x"b106",x"273e",x"3be5",x"396c",x"3915"),
(x"2ed8",x"3adf",x"3717",x"b273",x"2f43",x"3bc8",x"3972",x"3920",x"2ec2",x"3ace",x"3715",x"b468",x"247a",x"3bb0",x"3971",x"3916",x"2ea0",x"3ae3",x"3710",x"b550",x"2e33",x"3b81",x"396e",x"3922"),
(x"2f3c",x"3aed",x"3711",x"2e23",x"2a2e",x"3bf4",x"3978",x"3928",x"2ed8",x"3adf",x"3717",x"b273",x"2f43",x"3bc8",x"3972",x"3920",x"2ef8",x"3af2",x"3712",x"ab5f",x"2345",x"3bfc",x"3974",x"392b"),
(x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d",x"2fc1",x"3aef",x"3713",x"a5b5",x"b7de",x"3af6",x"3981",x"392a",x"2f7e",x"3aef",x"3712",x"add2",x"b04b",x"3be4",x"397d",x"3929"),
(x"2fc5",x"3b01",x"3716",x"2553",x"32c7",x"3bd1",x"3981",x"3934",x"2ff2",x"3afd",x"3718",x"2e36",x"a153",x"3bf6",x"3984",x"3932",x"2fad",x"3afe",x"3716",x"af4d",x"aa5f",x"3bf0",x"397f",x"3932"),
(x"300c",x"3aff",x"3716",x"2f15",x"329c",x"3bc6",x"3986",x"3933",x"2ff2",x"3afd",x"3718",x"2e36",x"a153",x"3bf6",x"3984",x"3932",x"2fc5",x"3b01",x"3716",x"2553",x"32c7",x"3bd1",x"3981",x"3934"),
(x"2f8e",x"3b1f",x"370f",x"2edc",x"2cd0",x"3bee",x"397d",x"3945",x"2fe3",x"3b15",x"3713",x"2da1",x"2f14",x"3beb",x"3982",x"3940",x"2f3b",x"3b15",x"3717",x"30e7",x"3057",x"3bd4",x"3977",x"393f"),
(x"2f5a",x"3b33",x"3716",x"2adf",x"a6b5",x"3bfc",x"3978",x"3951",x"2f8e",x"3b1f",x"370f",x"2edc",x"2cd0",x"3bee",x"397d",x"3945",x"2eeb",x"3b30",x"3713",x"29b8",x"a6e9",x"3bfd",x"3971",x"394e"),
(x"2f5a",x"3b33",x"3716",x"2adf",x"a6b5",x"3bfc",x"3978",x"3951",x"2eeb",x"3b30",x"3713",x"29b8",x"a6e9",x"3bfd",x"3971",x"394e",x"2ee1",x"3b4b",x"3717",x"2bf6",x"25ae",x"3bfb",x"396f",x"395d"),
(x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971",x"2ee1",x"3b4b",x"3717",x"2bf6",x"25ae",x"3bfb",x"396f",x"395d",x"2ebe",x"3b62",x"370f",x"b6c9",x"2fac",x"3b2e",x"396c",x"396a"),
(x"2ebe",x"3b62",x"370f",x"b6c9",x"2fac",x"3b2e",x"396c",x"396a",x"2ecd",x"3b69",x"370d",x"b809",x"2e09",x"3add",x"396c",x"396e",x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971"),
(x"2f10",x"3b90",x"370e",x"afd2",x"2717",x"3bef",x"396f",x"3984",x"3007",x"3b85",x"3715",x"ad56",x"20d0",x"3bf8",x"3980",x"3980",x"2efa",x"3b7a",x"3712",x"a9f0",x"2b1d",x"3bfa",x"396e",x"3978"),
(x"2ffb",x"3b6c",x"3715",x"3b82",x"b440",x"330f",x"396d",x"305d",x"300f",x"3b6a",x"36eb",x"3b89",x"b473",x"31fc",x"3972",x"3059",x"2f8b",x"3b48",x"370e",x"3b5f",x"b5f1",x"2f4d",x"396b",x"3036"),
(x"302f",x"3a2c",x"3710",x"bbfd",x"a997",x"a09b",x"3964",x"3071",x"302b",x"3a1c",x"3714",x"bbeb",x"308b",x"98b5",x"3964",x"3061",x"302e",x"3a20",x"36eb",x"bbf5",x"2e59",x"2467",x"395f",x"3064"),
(x"2ff3",x"3a58",x"3714",x"bb1c",x"b754",x"223f",x"3964",x"30a1",x"3024",x"3a3e",x"3713",x"bba5",x"b497",x"ac28",x"3964",x"3084",x"3029",x"3a3e",x"36eb",x"bba1",x"b4cc",x"1f45",x"395f",x"3084"),
(x"3021",x"3a14",x"3712",x"bb76",x"35c5",x"204d",x"3964",x"3057",x"300e",x"3a0d",x"3714",x"b95a",x"39f1",x"2032",x"3964",x"304f",x"301c",x"3a11",x"36eb",x"bab1",x"3862",x"21f0",x"395f",x"3054"),
(x"2fe4",x"3a08",x"3714",x"b5bf",x"3b76",x"27db",x"3964",x"3046",x"2fe9",x"3a09",x"36eb",x"b7e1",x"3af5",x"269a",x"395f",x"3046",x"300e",x"3a0d",x"3714",x"b95a",x"39f1",x"2032",x"3964",x"304f"),
(x"2f7e",x"3a04",x"3715",x"2836",x"3bfd",x"294f",x"3964",x"3038",x"2f83",x"3a06",x"36eb",x"b03c",x"3beb",x"299b",x"395f",x"3038",x"2fe4",x"3a08",x"3714",x"b5bf",x"3b76",x"27db",x"3964",x"3046"),
(x"2f19",x"3a07",x"3716",x"386f",x"3aa7",x"2604",x"3964",x"302a",x"2f1b",x"3a08",x"36eb",x"3868",x"3aab",x"296a",x"395f",x"302b",x"2f7e",x"3a04",x"3715",x"2836",x"3bfd",x"294f",x"3964",x"3038"),
(x"2f19",x"3a07",x"3716",x"386f",x"3aa7",x"2604",x"3964",x"302a",x"2ec8",x"3a14",x"3714",x"3b01",x"37b5",x"2839",x"3964",x"301a",x"2f1b",x"3a08",x"36eb",x"3868",x"3aab",x"296a",x"395f",x"302b"),
(x"2eb5",x"3a1f",x"3714",x"3be6",x"b10f",x"9bfc",x"3964",x"300d",x"2eb5",x"3a1e",x"36eb",x"3bf9",x"2d11",x"2511",x"395f",x"300f",x"2ec8",x"3a14",x"3714",x"3b01",x"37b5",x"2839",x"3964",x"301a"),
(x"2ed5",x"3a28",x"3715",x"3928",x"ba1d",x"1553",x"3964",x"3003",x"2ecf",x"3a28",x"36eb",x"390c",x"ba34",x"2532",x"395f",x"3005",x"2eb5",x"3a1f",x"3714",x"3be6",x"b10f",x"9bfc",x"3964",x"300d"),
(x"2ed5",x"3a28",x"3715",x"3928",x"ba1d",x"1553",x"3bac",x"3ad8",x"2f14",x"3a29",x"3714",x"afe2",x"bbee",x"28fd",x"3baa",x"3ad9",x"2ecf",x"3a28",x"36eb",x"390c",x"ba34",x"2532",x"3bad",x"3add"),
(x"2f14",x"3a29",x"3714",x"afe2",x"bbee",x"28fd",x"3baa",x"3ad9",x"2f4a",x"3a25",x"3711",x"b64f",x"bb52",x"2d1b",x"3ba8",x"3ada",x"2f19",x"3a28",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3baa",x"3add"),
(x"2f99",x"3a42",x"3713",x"3bc2",x"33a4",x"298a",x"3b9c",x"3ad9",x"2f9f",x"3a42",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b9b",x"3ade",x"2faf",x"3a3e",x"3711",x"3a7a",x"38b0",x"283c",x"3b9d",x"3ada"),
(x"2f4a",x"3a25",x"3711",x"b64f",x"bb52",x"2d1b",x"3ba8",x"3ada",x"2f9c",x"3a24",x"3710",x"3416",x"bbad",x"2f8d",x"3ba5",x"3ada",x"2f44",x"3a23",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3ba9",x"3ade"),
(x"301b",x"3acc",x"3713",x"b583",x"bb63",x"3153",x"3958",x"2f26",x"3013",x"3ac9",x"36eb",x"b5e4",x"bb4d",x"31a2",x"395a",x"2f00",x"2ff0",x"3ad5",x"370f",x"ba9c",x"b854",x"30fa",x"3955",x"2f17"),
(x"2ffb",x"3b6c",x"3715",x"3b82",x"b440",x"330f",x"396d",x"305d",x"3007",x"3b85",x"3715",x"3bc5",x"2b9a",x"3358",x"396e",x"3078",x"300f",x"3b6a",x"36eb",x"3b89",x"b473",x"31fc",x"3972",x"3059"),
(x"2faf",x"3a3e",x"3711",x"340c",x"26c2",x"3bbc",x"3981",x"38c5",x"2fd1",x"3a38",x"3710",x"2856",x"a9ab",x"3bfc",x"3983",x"38c2",x"2f3e",x"3a43",x"3718",x"2b65",x"b528",x"3b8f",x"3979",x"38c8"),
(x"2f14",x"3b70",x"3715",x"bbd7",x"b1f9",x"2c2a",x"3967",x"30d0",x"2f10",x"3b6d",x"3716",x"b8de",x"3a56",x"297d",x"3967",x"30d2",x"2f0d",x"3b6e",x"36eb",x"bbe3",x"2ce8",x"30c3",x"396b",x"30de"),
(x"2ef8",x"3af2",x"3712",x"b84e",x"3ab0",x"2ec7",x"3966",x"2ab9",x"2ea0",x"3ae3",x"3710",x"bb6a",x"35bb",x"2efe",x"3967",x"2b07",x"2ee2",x"3af4",x"36eb",x"b958",x"39de",x"2fe4",x"396b",x"2ab5"),
(x"2fc4",x"3a29",x"3711",x"3a7e",x"b887",x"3089",x"3ba3",x"3ada",x"2fd3",x"3a27",x"36eb",x"3aa4",x"b859",x"2fe5",x"3ba3",x"3ade",x"2f9c",x"3a24",x"3710",x"3416",x"bbad",x"2f8d",x"3ba5",x"3ada"),
(x"2f55",x"3a48",x"3718",x"bbe6",x"309e",x"2baa",x"3930",x"2400",x"2f4a",x"3a48",x"36eb",x"bbe6",x"308e",x"2c41",x"3935",x"238d",x"2f5a",x"3a5b",x"3715",x"bbfa",x"a70a",x"2c48",x"392e",x"22c2"),
(x"2fc4",x"3a29",x"3711",x"3a7e",x"b887",x"3089",x"3ba3",x"3ada",x"2fdc",x"3a30",x"3710",x"3bcc",x"b227",x"2f2f",x"3ba1",x"3ada",x"2fd3",x"3a27",x"36eb",x"3aa4",x"b859",x"2fe5",x"3ba3",x"3ade"),
(x"2ff0",x"3ad5",x"370f",x"ba9c",x"b854",x"30fa",x"3955",x"2f17",x"2fdc",x"3ad4",x"36eb",x"bb7d",x"b521",x"3095",x"3957",x"2ef3",x"2ff4",x"3adb",x"370e",x"bb25",x"370e",x"2d6a",x"3954",x"2f12"),
(x"3044",x"3a9a",x"3714",x"3972",x"b9bb",x"30de",x"3914",x"2857",x"3048",x"3a97",x"36eb",x"36fe",x"bb25",x"2ea4",x"3919",x"283d",x"3000",x"3a94",x"3711",x"34dc",x"bb97",x"2d61",x"3913",x"280e"),
(x"2faf",x"3a3e",x"3711",x"3a7a",x"38b0",x"283c",x"3b9d",x"3ada",x"2fb1",x"3a3e",x"36eb",x"39db",x"396c",x"2c1a",x"3b9d",x"3ade",x"2fd1",x"3a38",x"3710",x"3b2f",x"36d9",x"2e52",x"3b9f",x"3ada"),
(x"2fad",x"3afe",x"3716",x"b7e9",x"3af1",x"2aa7",x"3965",x"2a51",x"2ef8",x"3af2",x"3712",x"b84e",x"3ab0",x"2ec7",x"3966",x"2ab9",x"2fb4",x"3b00",x"36eb",x"b776",x"3b0b",x"2d41",x"396a",x"2a3e"),
(x"2f4b",x"3a60",x"3715",x"b95d",x"b9e3",x"2de3",x"392e",x"2274",x"2f5a",x"3a5b",x"3715",x"bbfa",x"a70a",x"2c48",x"392e",x"22c2",x"2f48",x"3a5e",x"36eb",x"b9df",x"b964",x"2d28",x"3933",x"222b"),
(x"3013",x"3ae4",x"3713",x"bb5b",x"3634",x"2c08",x"3951",x"2f12",x"2ff4",x"3adb",x"370e",x"bb25",x"370e",x"2d6a",x"3954",x"2f12",x"300f",x"3ae5",x"36eb",x"bad3",x"3822",x"2c4d",x"3953",x"2ee9"),
(x"2f5a",x"3b33",x"3716",x"3bff",x"20a8",x"2138",x"3969",x"3021",x"2f8b",x"3b48",x"370e",x"3b5f",x"b5f1",x"2f4d",x"396b",x"3036",x"2f5b",x"3b33",x"36eb",x"3bfe",x"1e8d",x"2828",x"396e",x"301b"),
(x"2fad",x"3afe",x"3716",x"b7e9",x"3af1",x"2aa7",x"3965",x"2a51",x"2fb4",x"3b00",x"36eb",x"b776",x"3b0b",x"2d41",x"396a",x"2a3e",x"2fc5",x"3b01",x"3716",x"bbde",x"31b5",x"2825",x"3965",x"2a3f"),
(x"2ef3",x"3a69",x"3719",x"b9a6",x"b994",x"2faf",x"392d",x"2190",x"2f4b",x"3a60",x"3715",x"b95d",x"b9e3",x"2de3",x"392e",x"2274",x"2ed5",x"3a69",x"36eb",x"b9ed",x"b94b",x"2f45",x"3932",x"2101"),
(x"2fe3",x"3a91",x"3711",x"3b12",x"b763",x"2ca3",x"392c",x"2a7d",x"3000",x"3a94",x"3711",x"34dc",x"bb97",x"2d61",x"392b",x"2a91",x"2ff6",x"3a93",x"36eb",x"37d8",x"baf6",x"2a35",x"3930",x"2a9b"),
(x"3014",x"3ae7",x"3713",x"bb09",x"b791",x"2ab8",x"3950",x"2f10",x"3013",x"3ae4",x"3713",x"bb5b",x"3634",x"2c08",x"3951",x"2f12",x"3010",x"3ae7",x"36eb",x"b9e9",x"b955",x"2e31",x"3952",x"2ee7"),
(x"2f5a",x"3b33",x"3716",x"3bff",x"20a8",x"2138",x"3969",x"3021",x"2f5b",x"3b33",x"36eb",x"3bfe",x"1e8d",x"2828",x"396e",x"301b",x"2f8e",x"3b1f",x"370f",x"3ad7",x"3821",x"29e6",x"3969",x"300a"),
(x"2fc5",x"3b01",x"3716",x"bbde",x"31b5",x"2825",x"3950",x"3126",x"2fc0",x"3b01",x"36eb",x"bb24",x"b71c",x"2cde",x"3954",x"3138",x"2fb0",x"3b06",x"3714",x"b9e8",x"b951",x"2f27",x"3952",x"3123"),
(x"2ef3",x"3a69",x"3719",x"b9a6",x"b994",x"2faf",x"392d",x"2190",x"2ed5",x"3a69",x"36eb",x"b9ed",x"b94b",x"2f45",x"3932",x"2101",x"2ef4",x"3a6b",x"3719",x"b250",x"3bca",x"2f22",x"392d",x"2173"),
(x"2fd7",x"3a8d",x"3712",x"3bf7",x"2843",x"2d8f",x"392c",x"2a6d",x"2fe5",x"3a8c",x"36eb",x"3bf8",x"a379",x"2d44",x"3930",x"2a7d",x"2fe6",x"3a82",x"3712",x"3b92",x"3509",x"2cb4",x"392d",x"2a40"),
(x"3000",x"3aec",x"3710",x"b833",x"bac7",x"2d1d",x"3915",x"2b3b",x"3014",x"3ae7",x"3713",x"bb09",x"b791",x"2ab8",x"3915",x"2b58",x"3010",x"3ae7",x"36eb",x"b9e9",x"b955",x"2e31",x"391a",x"2b4c"),
(x"2fe3",x"3b15",x"3713",x"37c2",x"3af3",x"2e28",x"3968",x"2ff8",x"2f8e",x"3b1f",x"370f",x"3ad7",x"3821",x"29e6",x"3969",x"300a",x"2fee",x"3b17",x"36eb",x"373f",x"3b1a",x"2d3c",x"396d",x"2fef"),
(x"2fb0",x"3b06",x"3714",x"b9e8",x"b951",x"2f27",x"3952",x"3123",x"2f9f",x"3b05",x"36eb",x"b97a",x"b9b6",x"309a",x"3955",x"3135",x"2f3b",x"3b15",x"3717",x"ba77",x"b889",x"310c",x"3956",x"3116"),
(x"2f3d",x"3a6b",x"3718",x"b0c6",x"3be6",x"2ad9",x"392b",x"20f4",x"2ef4",x"3a6b",x"3719",x"b250",x"3bca",x"2f22",x"392d",x"2173",x"2f48",x"3a6c",x"36eb",x"bb01",x"3745",x"3141",x"3930",x"2008"),
(x"2fe6",x"3a82",x"3712",x"3b92",x"3509",x"2cb4",x"392d",x"2a40",x"2fee",x"3a84",x"36eb",x"3b57",x"3625",x"2e99",x"3931",x"2a5c",x"302e",x"3a60",x"3711",x"3b70",x"3585",x"3014",x"392f",x"29ac"),
(x"2f7e",x"3aef",x"3712",x"32e8",x"bbcb",x"2c10",x"3914",x"2af5",x"2fc1",x"3aef",x"3713",x"b0a8",x"bbea",x"22dc",x"3914",x"2b18",x"2fb8",x"3aef",x"36eb",x"b046",x"bbe8",x"2cb7",x"3919",x"2b0c"),
(x"2fe3",x"3b15",x"3713",x"37c2",x"3af3",x"2e28",x"3968",x"2ff8",x"2fee",x"3b17",x"36eb",x"373f",x"3b1a",x"2d3c",x"396d",x"2fef",x"3001",x"3b16",x"3712",x"b721",x"3b24",x"2bf2",x"3968",x"2fef"),
(x"2f3b",x"3b15",x"3717",x"ba77",x"b889",x"310c",x"3956",x"3116",x"2f20",x"3b14",x"36eb",x"baff",x"b73c",x"3197",x"3959",x"3128",x"2eeb",x"3b30",x"3713",x"bbc6",x"b1be",x"30de",x"395c",x"3104"),
(x"302e",x"3a60",x"3711",x"3b70",x"3585",x"3014",x"392f",x"29ac",x"303d",x"3a5e",x"36eb",x"3b99",x"345f",x"30d6",x"3934",x"29b7",x"3046",x"3a41",x"3711",x"3be4",x"2d1d",x"308b",x"3931",x"292a"),
(x"2ed8",x"3adf",x"3717",x"3b6f",x"b5e5",x"261e",x"3913",x"2a83",x"2f3c",x"3aed",x"3711",x"3934",x"ba0d",x"2c18",x"3914",x"2ad1",x"2ede",x"3adf",x"36eb",x"3aaf",x"b860",x"2a70",x"3919",x"2a84"),
(x"3001",x"3b16",x"3712",x"b721",x"3b24",x"2bf2",x"3968",x"2fef",x"3004",x"3b18",x"36eb",x"b8ae",x"3a73",x"2d49",x"396c",x"2fe8",x"3017",x"3b1a",x"3711",x"b5dd",x"3b65",x"2eae",x"3968",x"2fe1"),
(x"2ee1",x"3b4b",x"3717",x"bbf0",x"af10",x"2aec",x"3960",x"30ef",x"2eeb",x"3b30",x"3713",x"bbc6",x"b1be",x"30de",x"395c",x"3104",x"2ed7",x"3b4b",x"36eb",x"bbea",x"ae09",x"2f12",x"3964",x"3101"),
(x"2f49",x"3a6d",x"3718",x"baf5",x"b7e1",x"2460",x"3965",x"2ca9",x"2f3d",x"3a6b",x"3718",x"b0c6",x"3be6",x"2ad9",x"3965",x"2cae",x"2f48",x"3a6c",x"36eb",x"bb01",x"3745",x"3141",x"396a",x"2cb1"),
(x"3046",x"3a1f",x"3714",x"3bec",x"ad02",x"2f52",x"3933",x"289e",x"3046",x"3a41",x"3711",x"3be4",x"2d1d",x"308b",x"3931",x"292a",x"304f",x"3a1e",x"36eb",x"3be8",x"ad66",x"3010",x"3938",x"28b0"),
(x"2ec2",x"3ace",x"3715",x"3bfe",x"2412",x"2867",x"3914",x"2a3d",x"2ed8",x"3adf",x"3717",x"3b6f",x"b5e5",x"261e",x"3913",x"2a83",x"2ec6",x"3acf",x"36eb",x"3bfa",x"ac62",x"2617",x"3919",x"2a40"),
(x"3017",x"3b1a",x"3711",x"b5dd",x"3b65",x"2eae",x"3968",x"2fe1",x"3014",x"3b1c",x"36eb",x"ae29",x"3be6",x"3005",x"396c",x"2fdc",x"3038",x"3b19",x"3712",x"35a5",x"3b63",x"30cc",x"3967",x"2fd0"),
(x"2ee1",x"3b4b",x"3717",x"bbf0",x"af10",x"2aec",x"3960",x"30ef",x"2ed7",x"3b4b",x"36eb",x"bbea",x"ae09",x"2f12",x"3964",x"3101",x"2ebe",x"3b62",x"370f",x"bbdd",x"b0de",x"2e6c",x"3965",x"30e2"),
(x"2f16",x"3a73",x"3715",x"b9d1",x"b974",x"2cc6",x"3966",x"2c96",x"2ef5",x"3a75",x"36eb",x"ba0e",x"b929",x"2e78",x"396b",x"2c95",x"2ede",x"3a7e",x"3718",x"bb13",x"b732",x"2fec",x"3966",x"2c7c"),
(x"3046",x"3a1f",x"3714",x"3bec",x"ad02",x"2f52",x"3933",x"289e",x"304f",x"3a1e",x"36eb",x"3be8",x"ad66",x"3010",x"3938",x"28b0",x"3036",x"3a0f",x"3712",x"3b45",x"b640",x"30a6",x"3934",x"285e"),
(x"2fdc",x"3a30",x"3710",x"3bcc",x"b227",x"2f2f",x"3ba1",x"3ada",x"2fd1",x"3a38",x"3710",x"3b2f",x"36d9",x"2e52",x"3b9f",x"3ada",x"2fec",x"3a30",x"36eb",x"3bf4",x"9ef6",x"2eb6",x"3ba1",x"3ade"),
(x"2ece",x"3ab8",x"3714",x"3b81",x"3558",x"2da6",x"3914",x"29e0",x"2ec2",x"3ace",x"3715",x"3bfe",x"2412",x"2867",x"3914",x"2a3d",x"2ed7",x"3aba",x"36eb",x"3bcf",x"32aa",x"2bc8",x"3919",x"29e8"),
(x"3038",x"3b19",x"3712",x"35a5",x"3b63",x"30cc",x"3967",x"2fd0",x"3043",x"3b1c",x"36eb",x"3913",x"3a0d",x"310f",x"396c",x"2fc3",x"304c",x"3b12",x"3711",x"3bb2",x"332f",x"30f4",x"3967",x"2fbd"),
(x"2ebe",x"3b62",x"370f",x"bbdd",x"b0de",x"2e6c",x"3965",x"30e2",x"2eaa",x"3b61",x"36eb",x"bbe4",x"aadf",x"30ee",x"3968",x"30f1",x"2ecd",x"3b69",x"370d",x"bb0d",x"370c",x"3169",x"3966",x"30de"),
(x"2ede",x"3a7e",x"3718",x"bb13",x"b732",x"2fec",x"3966",x"2c7c",x"2ec6",x"3a7d",x"36eb",x"bbbf",x"b333",x"2ed2",x"396b",x"2c80",x"2ed4",x"3a86",x"3712",x"bbf0",x"2c20",x"2e95",x"3967",x"2c6b"),
(x"3036",x"3a0f",x"3712",x"3b45",x"b640",x"30a6",x"3934",x"285e",x"303e",x"3a0c",x"36eb",x"3ab2",x"b834",x"30cf",x"3939",x"2865",x"3003",x"3a00",x"3715",x"393c",x"b9e9",x"311d",x"3934",x"280a"),
(x"2f11",x"3aa9",x"3715",x"3a65",x"38c1",x"2d9e",x"3914",x"2997",x"2ece",x"3ab8",x"3714",x"3b81",x"3558",x"2da6",x"3914",x"29e0",x"2f1f",x"3aaa",x"36eb",x"3ac2",x"3833",x"2e85",x"3919",x"299b"),
(x"304c",x"3b12",x"3711",x"3bb2",x"332f",x"30f4",x"3967",x"2fbd",x"3057",x"3b12",x"36eb",x"3be5",x"adbc",x"3036",x"396b",x"2fae",x"303e",x"3b06",x"3712",x"3ae4",x"b7c4",x"30c9",x"3965",x"2fa8"),
(x"2ee7",x"3b6c",x"3713",x"b451",x"3bac",x"2d81",x"3966",x"30d8",x"2ecd",x"3b69",x"370d",x"bb0d",x"370c",x"3169",x"3966",x"30de",x"2ee1",x"3b6e",x"36eb",x"b571",x"3b6d",x"30cc",x"396a",x"30e3"),
(x"2ed4",x"3a86",x"3712",x"bbf0",x"2c20",x"2e95",x"3967",x"2c6b",x"2ecb",x"3a89",x"36eb",x"bbbf",x"3370",x"2dad",x"396c",x"2c68",x"2ee4",x"3a89",x"3712",x"b297",x"3bcc",x"2d84",x"3967",x"2c63"),
(x"3003",x"3a00",x"3715",x"393c",x"b9e9",x"311d",x"3934",x"280a",x"3007",x"39fc",x"36eb",x"37cb",x"bae6",x"3068",x"393a",x"280f",x"2f91",x"39fb",x"3715",x"1ef6",x"bbee",x"302a",x"3935",x"2791"),
(x"2f5a",x"3a9f",x"3717",x"3939",x"3a0b",x"29e0",x"3914",x"2960",x"2f11",x"3aa9",x"3715",x"3a65",x"38c1",x"2d9e",x"3914",x"2997",x"2f61",x"3aa0",x"36eb",x"39cd",x"3979",x"2caa",x"3919",x"2965"),
(x"303e",x"3b06",x"3712",x"3ae4",x"b7c4",x"30c9",x"3965",x"2fa8",x"3044",x"3b03",x"36eb",x"3902",x"ba23",x"306a",x"3969",x"2f90",x"301b",x"3b03",x"3713",x"3607",x"bb5e",x"2e4f",x"3964",x"2f98"),
(x"2f10",x"3b6d",x"3716",x"b8de",x"3a56",x"297d",x"3967",x"30d2",x"2ee7",x"3b6c",x"3713",x"b451",x"3bac",x"2d81",x"3966",x"30d8",x"2f0d",x"3b6e",x"36eb",x"bbe3",x"2ce8",x"30c3",x"396b",x"30de"),
(x"2f1d",x"3a89",x"3717",x"aa07",x"3bfc",x"284d",x"3966",x"2c54",x"2ee4",x"3a89",x"3712",x"b297",x"3bcc",x"2d84",x"3967",x"2c63",x"2f24",x"3a8a",x"36eb",x"ac58",x"3bf7",x"2bc1",x"396b",x"2c4e"),
(x"2f0e",x"3a00",x"3713",x"b82e",x"baba",x"306c",x"3935",x"2702",x"2f91",x"39fb",x"3715",x"1ef6",x"bbee",x"302a",x"3935",x"2791",x"2f13",x"39fc",x"36eb",x"b66a",x"bb44",x"2f81",x"393a",x"270e"),
(x"2f7f",x"3a9c",x"3717",x"ac93",x"3bf9",x"2918",x"3914",x"2949",x"2f5a",x"3a9f",x"3717",x"3939",x"3a0b",x"29e0",x"3914",x"2960",x"2f7e",x"3a9d",x"36eb",x"b5a6",x"3b74",x"2d53",x"3919",x"2952"),
(x"300c",x"3aff",x"3716",x"3ac7",x"383c",x"283f",x"3963",x"2f91",x"301b",x"3b03",x"3713",x"3607",x"bb5e",x"2e4f",x"3964",x"2f98",x"300f",x"3aff",x"36eb",x"394d",x"39f2",x"2dc5",x"3967",x"2f78"),
(x"2f8b",x"3b48",x"370e",x"3004",x"a717",x"3bef",x"397b",x"395d",x"2f5a",x"3b33",x"3716",x"2adf",x"a6b5",x"3bfc",x"3978",x"3951",x"2ee1",x"3b4b",x"3717",x"2bf6",x"25ae",x"3bfb",x"396f",x"395d"),
(x"2f1d",x"3a89",x"3717",x"aa07",x"3bfc",x"284d",x"3966",x"2c54",x"2f24",x"3a8a",x"36eb",x"ac58",x"3bf7",x"2bc1",x"396b",x"2c4e",x"2f3a",x"3a8a",x"3716",x"b8f4",x"3a42",x"2c09",x"3966",x"2c4c"),
(x"2e95",x"3a0c",x"3715",x"bae0",x"b7cf",x"30d4",x"3934",x"265f",x"2f0e",x"3a00",x"3713",x"b82e",x"baba",x"306c",x"3935",x"2702",x"2e80",x"3a0a",x"36eb",x"b9f2",x"b938",x"30b5",x"393a",x"2650"),
(x"2fa9",x"3aa0",x"3714",x"b9a7",x"399f",x"2d1e",x"3914",x"2930",x"2f7f",x"3a9c",x"3717",x"ac93",x"3bf9",x"2918",x"3914",x"2949",x"2f7e",x"3a9d",x"36eb",x"b5a6",x"3b74",x"2d53",x"3919",x"2952"),
(x"300c",x"3aff",x"3716",x"3ac7",x"383c",x"283f",x"3963",x"2f91",x"300f",x"3aff",x"36eb",x"394d",x"39f2",x"2dc5",x"3967",x"2f78",x"302f",x"3afb",x"3711",x"38c8",x"3a4e",x"30a8",x"3962",x"2f7c"),
(x"2f3a",x"3a8a",x"3716",x"b8f4",x"3a42",x"2c09",x"3966",x"2c4c",x"2f37",x"3a8c",x"36eb",x"bb71",x"b58a",x"2fc3",x"396b",x"2c47",x"2f48",x"3a8d",x"3715",x"bac1",x"b812",x"3146",x"3966",x"2c44"),
(x"2e5f",x"3a1e",x"3715",x"bbec",x"abe2",x"2fce",x"3934",x"25be",x"2e95",x"3a0c",x"3715",x"bae0",x"b7cf",x"30d4",x"3934",x"265f",x"2e4e",x"3a1d",x"36eb",x"bbc4",x"b27a",x"3012",x"3939",x"25a9"),
(x"2fd3",x"3aa6",x"3714",x"b97e",x"39c5",x"2dbf",x"3915",x"290e",x"2fd6",x"3aa9",x"36eb",x"b976",x"39cc",x"2dcc",x"391a",x"290f",x"300a",x"3aad",x"3716",x"b7d6",x"3af0",x"2d8e",x"3915",x"28e1"),
(x"302f",x"3afb",x"3711",x"38c8",x"3a4e",x"30a8",x"3962",x"2f7c",x"303f",x"3afc",x"36eb",x"39ec",x"392b",x"31e5",x"3966",x"2f62",x"3058",x"3aeb",x"370f",x"3b4b",x"35cc",x"3223",x"395f",x"2f5b"),
(x"2efa",x"3b7a",x"3712",x"bbcf",x"b081",x"3141",x"3969",x"30c7",x"2edb",x"3b7b",x"36eb",x"bbdb",x"1c67",x"320a",x"396d",x"30d2",x"2f10",x"3b90",x"370e",x"bb7b",x"34a9",x"3270",x"396c",x"30b5"),
(x"2f3c",x"3a92",x"3714",x"3879",x"347b",x"3a3d",x"3966",x"2c3b",x"2f48",x"3a8d",x"3715",x"bac1",x"b812",x"3146",x"3966",x"2c44",x"2f06",x"3a9a",x"3718",x"bac6",x"b7dc",x"3286",x"3966",x"2c25"),
(x"2e70",x"3a2f",x"3717",x"bb55",x"35fd",x"307e",x"3933",x"2533",x"2e5f",x"3a1e",x"3715",x"bbec",x"abe2",x"2fce",x"3934",x"25be",x"2e58",x"3a30",x"36eb",x"bb6e",x"3575",x"309e",x"3938",x"250b"),
(x"2ff3",x"3a58",x"3714",x"305e",x"2194",x"3bec",x"3985",x"38d4",x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"302e",x"3a60",x"3711",x"3115",x"27d5",x"3be4",x"398c",x"38d9"),
(x"300a",x"3aad",x"3716",x"b7d6",x"3af0",x"2d8e",x"3915",x"28e1",x"3008",x"3aae",x"36eb",x"b53f",x"3b87",x"2d28",x"391a",x"28e9",x"302b",x"3aae",x"3716",x"2345",x"3bf7",x"2dcc",x"3915",x"28be"),
(x"3058",x"3aeb",x"370f",x"3b4b",x"35cc",x"3223",x"395f",x"2f5b",x"3065",x"3aeb",x"36eb",x"3bbc",x"3212",x"3175",x"3963",x"2f41",x"305c",x"3ad8",x"370f",x"3bd3",x"af46",x"3182",x"395c",x"2f3f"),
(x"2f06",x"3a9a",x"3718",x"bac6",x"b7dc",x"3286",x"3966",x"2c25",x"2ed7",x"3a9c",x"36eb",x"badb",x"b7e7",x"30ac",x"396c",x"2c1e",x"2e9f",x"3ab2",x"3714",x"bb6b",x"b587",x"3096",x"3967",x"2bd9"),
(x"2e70",x"3a2f",x"3717",x"bb55",x"35fd",x"307e",x"3933",x"2533",x"2e58",x"3a30",x"36eb",x"bb6e",x"3575",x"309e",x"3938",x"250b",x"2ec0",x"3a3d",x"3711",x"b8a4",x"3a69",x"309a",x"3932",x"24a5"),
(x"302b",x"3aae",x"3716",x"2345",x"3bf7",x"2dcc",x"3915",x"28be",x"302e",x"3ab0",x"36eb",x"33e5",x"3bb4",x"2ec2",x"391a",x"28c0",x"3045",x"3aab",x"3714",x"3976",x"39c0",x"3024",x"3915",x"289f"),
(x"305c",x"3ad8",x"370f",x"3bd3",x"af46",x"3182",x"395c",x"2f3f",x"3068",x"3ad7",x"36eb",x"3b61",x"b5a0",x"3119",x"395f",x"2f23",x"3040",x"3acf",x"370f",x"3891",x"ba72",x"30f5",x"395a",x"2f2e"),
(x"2f10",x"3b90",x"370e",x"bb7b",x"34a9",x"3270",x"396c",x"30b5",x"2ef9",x"3b92",x"36eb",x"bade",x"37ab",x"31d3",x"3970",x"30bd",x"2f7a",x"3ba1",x"3712",x"b8b5",x"3a3e",x"32bc",x"396e",x"30a0"),
(x"2e9f",x"3ab2",x"3714",x"bb6b",x"b587",x"3096",x"3967",x"2bd9",x"2e89",x"3ab2",x"36eb",x"bbba",x"b376",x"2f14",x"396c",x"2bd6",x"2e7c",x"3acb",x"3712",x"bbf0",x"aa00",x"2f46",x"3967",x"2b6e"),
(x"2f3e",x"3a43",x"3718",x"b8ae",x"3a78",x"2b7c",x"3930",x"242e",x"2ec0",x"3a3d",x"3711",x"b8a4",x"3a69",x"309a",x"3932",x"24a5",x"2f34",x"3a43",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3935",x"23da"),
(x"3045",x"3aab",x"3714",x"3976",x"39c0",x"3024",x"3915",x"289f",x"3050",x"3aac",x"36eb",x"3acb",x"3812",x"3064",x"391a",x"2898",x"3050",x"3aa2",x"3712",x"3be0",x"2e5e",x"30a3",x"3915",x"287a"),
(x"301b",x"3acc",x"3713",x"b583",x"bb63",x"3153",x"3958",x"2f26",x"3040",x"3acf",x"370f",x"3891",x"ba72",x"30f5",x"395a",x"2f2e",x"3013",x"3ac9",x"36eb",x"b5e4",x"bb4d",x"31a2",x"395a",x"2f00"),
(x"2fbb",x"3ba1",x"3716",x"3add",x"375a",x"334d",x"396e",x"3097",x"2f7a",x"3ba1",x"3712",x"b8b5",x"3a3e",x"32bc",x"396e",x"30a0",x"2fd0",x"3ba6",x"36eb",x"3996",x"395f",x"33ec",x"3973",x"309a"),
(x"2e7c",x"3acb",x"3712",x"bbf0",x"aa00",x"2f46",x"3967",x"2b6e",x"2e6b",x"3acc",x"36eb",x"bbef",x"2d0b",x"2e69",x"396c",x"2b67",x"2ea0",x"3ae3",x"3710",x"bb6a",x"35bb",x"2efe",x"3967",x"2b07"),
(x"2f55",x"3a48",x"3718",x"bbe6",x"309e",x"2baa",x"3930",x"2400",x"2f3e",x"3a43",x"3718",x"b8ae",x"3a78",x"2b7c",x"3930",x"242e",x"2f4a",x"3a48",x"36eb",x"bbe6",x"308e",x"2c41",x"3935",x"238d"),
(x"3050",x"3aa2",x"3712",x"3be0",x"2e5e",x"30a3",x"3915",x"287a",x"305c",x"3aa1",x"36eb",x"3bcf",x"b173",x"3043",x"391a",x"286a",x"3044",x"3a9a",x"3714",x"3972",x"b9bb",x"30de",x"3914",x"2857"),
(x"3046",x"3a41",x"3711",x"2cd1",x"2504",x"3bf9",x"398f",x"38c7",x"3046",x"3a1f",x"3714",x"aeb0",x"28fa",x"3bf3",x"3990",x"38b4",x"302f",x"3a2c",x"3710",x"a828",x"260a",x"3bfe",x"398d",x"38bb"),
(x"3036",x"3a0f",x"3712",x"2587",x"208e",x"3bff",x"398e",x"38ab",x"300e",x"3a0d",x"3714",x"28bf",x"2c22",x"3bfa",x"3989",x"38aa",x"3021",x"3a14",x"3712",x"a953",x"27ae",x"3bfd",x"398b",x"38ae"),
(x"3036",x"3a0f",x"3712",x"2587",x"208e",x"3bff",x"398e",x"38ab",x"3003",x"3a00",x"3715",x"20ea",x"2afd",x"3bfc",x"3988",x"38a2",x"300e",x"3a0d",x"3714",x"28bf",x"2c22",x"3bfa",x"3989",x"38aa"),
(x"3003",x"3a00",x"3715",x"20ea",x"2afd",x"3bfc",x"3988",x"38a2",x"2f91",x"39fb",x"3715",x"a7e2",x"29b2",x"3bfc",x"3980",x"389f",x"2fe4",x"3a08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3986",x"38a7"),
(x"2f91",x"39fb",x"3715",x"a7e2",x"29b2",x"3bfc",x"3980",x"389f",x"2f0e",x"3a00",x"3713",x"ab1d",x"aee4",x"3bf0",x"3978",x"38a1",x"2f7e",x"3a04",x"3715",x"a70a",x"a779",x"3bfe",x"397f",x"38a4"),
(x"2f0e",x"3a00",x"3713",x"ab1d",x"aee4",x"3bf0",x"3978",x"38a1",x"2e95",x"3a0c",x"3715",x"2266",x"9d87",x"3bff",x"3970",x"38a8",x"2f19",x"3a07",x"3716",x"a4bc",x"aceb",x"3bf9",x"3978",x"38a5"),
(x"2e95",x"3a0c",x"3715",x"2266",x"9d87",x"3bff",x"3970",x"38a8",x"2e5f",x"3a1e",x"3715",x"2891",x"a7ce",x"3bfd",x"396c",x"38b2",x"2ec8",x"3a14",x"3714",x"28e0",x"299e",x"3bfc",x"3973",x"38ac"),
(x"2eb5",x"3a1f",x"3714",x"2538",x"a9ab",x"3bfd",x"3971",x"38b2",x"2e5f",x"3a1e",x"3715",x"2891",x"a7ce",x"3bfd",x"396c",x"38b2",x"2ed5",x"3a28",x"3715",x"2c67",x"28a5",x"3bf9",x"3973",x"38b8"),
(x"2e70",x"3a2f",x"3717",x"2d06",x"2793",x"3bf8",x"396c",x"38bb",x"2ec0",x"3a3d",x"3711",x"28d9",x"a52b",x"3bfe",x"3971",x"38c3",x"2ed5",x"3a28",x"3715",x"2c67",x"28a5",x"3bf9",x"3973",x"38b8"),
(x"2f14",x"3a29",x"3714",x"2a45",x"2b10",x"3bfa",x"3977",x"38b8",x"2fc4",x"3a29",x"3711",x"2bef",x"a8a8",x"3bfa",x"3982",x"38b9",x"2f4a",x"3a25",x"3711",x"2a66",x"b319",x"3bca",x"397b",x"38b6"),
(x"2f55",x"3a48",x"3718",x"3420",x"1418",x"3bba",x"397a",x"38cb",x"2f99",x"3a42",x"3713",x"341f",x"ac3a",x"3bb6",x"397f",x"38c7",x"2f3e",x"3a43",x"3718",x"2b65",x"b528",x"3b8f",x"3979",x"38c8"),
(x"2f5a",x"3a5b",x"3715",x"27ae",x"a4f0",x"3bfe",x"397b",x"38d6",x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"2f94",x"3a4b",x"3714",x"2de0",x"a4c2",x"3bf6",x"397f",x"38cc"),
(x"2fd1",x"3a38",x"3710",x"2856",x"a9ab",x"3bfc",x"3983",x"38c2",x"2fc4",x"3a29",x"3711",x"2bef",x"a8a8",x"3bfa",x"3982",x"38b9",x"2f14",x"3a29",x"3714",x"2a45",x"2b10",x"3bfa",x"3977",x"38b8"),
(x"3056",x"3980",x"3718",x"26a1",x"97c8",x"3bff",x"3977",x"31ab",x"301e",x"397e",x"3718",x"224c",x"a379",x"3bff",x"3973",x"31a9",x"3033",x"39b8",x"3715",x"21a1",x"23fc",x"3bff",x"3974",x"31f5"),
(x"2f5a",x"3a5b",x"3715",x"27ae",x"a4f0",x"3bfe",x"397b",x"38d6",x"2f4b",x"3a60",x"3715",x"a8bf",x"afdb",x"3bef",x"397a",x"38d8",x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da"),
(x"2f94",x"3a4b",x"3714",x"3bf3",x"ae23",x"2b27",x"3b9a",x"3ad9",x"2fb5",x"3a63",x"3718",x"39e5",x"b968",x"0000",x"3b93",x"3ad8",x"2fb5",x"3a63",x"36eb",x"3469",x"bb91",x"316a",x"3b93",x"3add"),
(x"2f13",x"3798",x"3715",x"2d56",x"a0d0",x"3bf8",x"394e",x"397d",x"3008",x"3783",x"370e",x"2fd2",x"a717",x"3bef",x"393d",x"3981",x"2f67",x"3761",x"3716",x"30f9",x"28b2",x"3be5",x"3947",x"398c"),
(x"2f13",x"3798",x"3715",x"bbc5",x"ab9a",x"3358",x"3993",x"306e",x"2f67",x"3761",x"3716",x"badd",x"b75a",x"334d",x"3994",x"308d",x"2eeb",x"3797",x"36eb",x"bb99",x"b315",x"330d",x"3998",x"306b"),
(x"2eea",x"384e",x"3713",x"a91b",x"ab55",x"3bfb",x"3956",x"3932",x"2f72",x"384b",x"3714",x"ac39",x"a9a5",x"3bf9",x"394d",x"3934",x"2f20",x"383b",x"3712",x"aa69",x"a87e",x"3bfc",x"3952",x"393d"),
(x"2ea4",x"384b",x"3712",x"aa73",x"aa97",x"3bfa",x"395b",x"3934",x"2ef3",x"3837",x"3711",x"a994",x"a977",x"3bfc",x"3955",x"393f",x"2e89",x"383f",x"3711",x"a481",x"a546",x"3bff",x"395c",x"393b"),
(x"2ef3",x"3837",x"3711",x"a994",x"a977",x"3bfc",x"3955",x"393f",x"2ea4",x"384b",x"3712",x"aa73",x"aa97",x"3bfa",x"395b",x"3934",x"2f20",x"383b",x"3712",x"aa69",x"a87e",x"3bfc",x"3952",x"393d"),
(x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929",x"2f2f",x"3854",x"3718",x"ae36",x"2153",x"3bf6",x"3952",x"392e",x"2ec3",x"3856",x"3711",x"afec",x"2c2c",x"3beb",x"3959",x"392e"),
(x"2ea1",x"3883",x"370f",x"9df0",x"2631",x"3bff",x"395d",x"3914",x"2eec",x"3885",x"3713",x"ae9c",x"b367",x"3bbd",x"3958",x"3912",x"2f2d",x"3876",x"370e",x"26d5",x"a5c2",x"3bfe",x"3953",x"391a"),
(x"2f2d",x"3876",x"370e",x"26d5",x"a5c2",x"3bfe",x"3953",x"391a",x"2efb",x"386d",x"3713",x"a538",x"2c79",x"3bfa",x"3956",x"3920",x"2ea1",x"3883",x"370f",x"9df0",x"2631",x"3bff",x"395d",x"3914"),
(x"2e69",x"3879",x"370f",x"acd8",x"271d",x"3bf9",x"3960",x"391a",x"2efb",x"386d",x"3713",x"a538",x"2c79",x"3bfa",x"3956",x"3920",x"2e71",x"3866",x"370f",x"aec5",x"9a24",x"3bf4",x"395f",x"3925"),
(x"2ec3",x"3856",x"3711",x"afec",x"2c2c",x"3beb",x"3959",x"392e",x"2efa",x"386a",x"3713",x"a7ef",x"a849",x"3bfd",x"3956",x"3922",x"2f21",x"3865",x"3710",x"ac5b",x"30a5",x"3be5",x"3953",x"3925"),
(x"2f4a",x"38c4",x"3712",x"af67",x"2981",x"3bf0",x"3950",x"38ef",x"2fda",x"38c4",x"3715",x"a6c2",x"2c63",x"3bfa",x"3947",x"38ee",x"2fa2",x"38b5",x"3717",x"aff2",x"2a7a",x"3bed",x"394b",x"38f7"),
(x"2e99",x"38b7",x"3714",x"1553",x"2b62",x"3bfc",x"395c",x"38f6",x"2ecb",x"38a3",x"3716",x"acd8",x"27e2",x"3bf9",x"3959",x"3901",x"2e81",x"38af",x"3712",x"b162",x"2345",x"3be2",x"395e",x"38fb"),
(x"2ecb",x"38a3",x"3716",x"acd8",x"27e2",x"3bf9",x"3959",x"3901",x"2e99",x"38b7",x"3714",x"1553",x"2b62",x"3bfc",x"395c",x"38f6",x"2f0c",x"38a4",x"3716",x"2818",x"2d04",x"3bf8",x"3954",x"3900"),
(x"2f21",x"38bd",x"3711",x"240b",x"2d5c",x"3bf8",x"3953",x"38f2",x"2f4f",x"38ab",x"3714",x"a4fd",x"2da9",x"3bf7",x"3950",x"38fd",x"2f0c",x"38a4",x"3716",x"2818",x"2d04",x"3bf8",x"3954",x"3900"),
(x"2f79",x"38b1",x"3714",x"b036",x"273e",x"3bed",x"394d",x"38f9",x"2f21",x"38bd",x"3711",x"240b",x"2d5c",x"3bf8",x"3953",x"38f2",x"2f3f",x"38c0",x"3711",x"b27d",x"975f",x"3bd5",x"3951",x"38f1"),
(x"2ec5",x"38f1",x"3711",x"b115",x"a7d5",x"3be4",x"395a",x"38d5",x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2f3b",x"38cf",x"3712",x"b146",x"ac91",x"3bde",x"3952",x"38e8"),
(x"3017",x"38e6",x"3719",x"a3bb",x"a7b4",x"3bfe",x"3942",x"38db",x"2fe4",x"38e6",x"3718",x"2138",x"2e95",x"3bf4",x"3947",x"38db",x"3017",x"38e8",x"3719",x"a90e",x"2f00",x"3bf2",x"3942",x"38da"),
(x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2fd6",x"38f1",x"3715",x"28bf",x"2fda",x"3bef",x"3948",x"38d5",x"2fe4",x"38e6",x"3718",x"2138",x"2e95",x"3bf4",x"3947",x"38db"),
(x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2fe4",x"38e6",x"3718",x"2138",x"2e95",x"3bf4",x"3947",x"38db",x"2fd8",x"38e4",x"3718",x"2b4f",x"a525",x"3bfc",x"3947",x"38dc"),
(x"3002",x"38c8",x"3717",x"2d2d",x"aecd",x"3bed",x"3944",x"38ec",x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"3022",x"38d3",x"3718",x"2cf2",x"991e",x"3bf9",x"3940",x"38e5"),
(x"3022",x"38d3",x"3718",x"2cf2",x"991e",x"3bf9",x"3940",x"38e5",x"3027",x"38cb",x"3712",x"359c",x"b36a",x"3b42",x"393f",x"38ea",x"3002",x"38c8",x"3717",x"2d2d",x"aecd",x"3bed",x"3944",x"38ec"),
(x"2f3b",x"38cf",x"3712",x"b146",x"ac91",x"3bde",x"3952",x"38e8",x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"2fe7",x"38c7",x"3716",x"b009",x"ada6",x"3be7",x"3946",x"38ec"),
(x"2fda",x"38c4",x"3715",x"a6c2",x"2c63",x"3bfa",x"3947",x"38ee",x"2f4a",x"38c4",x"3712",x"af67",x"2981",x"3bf0",x"3950",x"38ef",x"2fe7",x"38c7",x"3716",x"b009",x"ada6",x"3be7",x"3946",x"38ec"),
(x"2fc7",x"38b2",x"3717",x"97c8",x"1f79",x"3c00",x"3948",x"38f8",x"2fda",x"38c4",x"3715",x"a6c2",x"2c63",x"3bfa",x"3947",x"38ee",x"2fe5",x"38bf",x"3714",x"a581",x"2e8a",x"3bf4",x"3946",x"38f1"),
(x"302a",x"3899",x"3714",x"2dba",x"a266",x"3bf7",x"393f",x"3906",x"3008",x"38a8",x"3715",x"a51e",x"ad06",x"3bf9",x"3943",x"38fe",x"3041",x"389f",x"3714",x"175f",x"ac2c",x"3bfb",x"393c",x"3903"),
(x"302f",x"3883",x"3715",x"3468",x"a47a",x"3bb0",x"393e",x"3913",x"302a",x"3899",x"3714",x"2dba",x"a266",x"3bf7",x"393f",x"3906",x"3052",x"3886",x"3712",x"3106",x"a738",x"3be5",x"393a",x"3911"),
(x"3025",x"3872",x"3717",x"3273",x"af43",x"3bc8",x"3940",x"391c",x"302f",x"3883",x"3715",x"3468",x"a47a",x"3bb0",x"393e",x"3913",x"3041",x"386e",x"3710",x"3550",x"ae33",x"3b81",x"393c",x"391f"),
(x"2fe6",x"3864",x"3711",x"ae24",x"aa2e",x"3bf4",x"3946",x"3924",x"3025",x"3872",x"3717",x"3273",x"af43",x"3bc8",x"3940",x"391c",x"3015",x"385f",x"3712",x"2b5f",x"a345",x"3bfc",x"3942",x"3927"),
(x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929",x"2f61",x"3862",x"3713",x"25b5",x"37de",x"3af6",x"394f",x"3926",x"2fa3",x"3862",x"3712",x"2dd2",x"304b",x"3be4",x"394b",x"3926"),
(x"2f5c",x"3850",x"3716",x"a559",x"b2c7",x"3bd1",x"394f",x"3931",x"2f2f",x"3854",x"3718",x"ae36",x"2153",x"3bf6",x"3952",x"392e",x"2f75",x"3853",x"3716",x"2f4d",x"2a5f",x"3bf0",x"394d",x"392f"),
(x"2f0a",x"3852",x"3716",x"af15",x"b29c",x"3bc7",x"3954",x"3930",x"2f2f",x"3854",x"3718",x"ae36",x"2153",x"3bf6",x"3952",x"392e",x"2f5c",x"3850",x"3716",x"a559",x"b2c7",x"3bd1",x"394f",x"3931"),
(x"2f93",x"3832",x"370f",x"aedc",x"acd0",x"3bee",x"394b",x"3942",x"2f3e",x"383c",x"3713",x"ada3",x"af14",x"3beb",x"3950",x"393c",x"2fe6",x"383c",x"3717",x"b0e7",x"b057",x"3bd4",x"3945",x"393c"),
(x"2fc8",x"381e",x"3716",x"aadf",x"26b5",x"3bfc",x"3946",x"394d",x"2f93",x"3832",x"370f",x"aedc",x"acd0",x"3bee",x"394b",x"3942",x"301b",x"3821",x"3713",x"a9b8",x"26e9",x"3bfd",x"393f",x"394b"),
(x"2fc8",x"381e",x"3716",x"aadf",x"26b5",x"3bfc",x"3946",x"394d",x"301b",x"3821",x"3713",x"a9b8",x"26e9",x"3bfd",x"393f",x"394b",x"3020",x"3806",x"3717",x"abf6",x"a5ae",x"3bfb",x"393d",x"395a"),
(x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d",x"3020",x"3806",x"3717",x"abf6",x"a5ae",x"3bfb",x"393d",x"395a",x"3031",x"37df",x"370f",x"36c9",x"afac",x"3b2e",x"3939",x"3966"),
(x"3031",x"37df",x"370f",x"36c9",x"afac",x"3b2e",x"3939",x"3966",x"302a",x"37d1",x"370d",x"3809",x"ae09",x"3add",x"393a",x"396b",x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d"),
(x"3008",x"3783",x"370e",x"2fd2",x"a717",x"3bef",x"393d",x"3981",x"2f13",x"3798",x"3715",x"2d56",x"a0d0",x"3bf8",x"394e",x"397d",x"3013",x"37ae",x"3712",x"29f0",x"ab1d",x"3bfa",x"393c",x"3975"),
(x"2f27",x"37cb",x"3715",x"bb82",x"3440",x"330f",x"3992",x"3053",x"2f02",x"37ce",x"36eb",x"bb89",x"3473",x"31fc",x"3997",x"304e",x"2f97",x"3809",x"370e",x"bb5f",x"35f1",x"2f4f",x"3991",x"302c"),
(x"2ec4",x"3925",x"3710",x"3bfd",x"2997",x"a09b",x"394a",x"29a0",x"2eca",x"3935",x"3714",x"3beb",x"b08a",x"98ea",x"394a",x"29e1",x"2ec5",x"3931",x"36eb",x"3bf5",x"ae59",x"2467",x"394f",x"29ce"),
(x"2f2f",x"38f9",x"3714",x"3b1c",x"3754",x"223f",x"3949",x"28de",x"2ed8",x"3913",x"3713",x"3ba5",x"3497",x"ac28",x"3949",x"2954",x"2ece",x"3913",x"36eb",x"3ba1",x"34cc",x"1f45",x"394e",x"2951"),
(x"2edf",x"393d",x"3712",x"3b76",x"b5c5",x"204d",x"394a",x"2a06",x"2f06",x"3944",x"3714",x"395a",x"b9f1",x"2032",x"394a",x"2a28",x"2ee8",x"3940",x"36eb",x"3ab1",x"b862",x"21f0",x"394f",x"2a10"),
(x"2f3d",x"3949",x"3714",x"35bf",x"bb76",x"27db",x"394a",x"2a4c",x"2f38",x"3948",x"36eb",x"37e1",x"baf5",x"269a",x"394f",x"2a46",x"2f06",x"3944",x"3714",x"395a",x"b9f1",x"2032",x"394a",x"2a28"),
(x"2fa3",x"394d",x"3715",x"a836",x"bbfd",x"294f",x"394a",x"2a84",x"2f9e",x"394c",x"36eb",x"303c",x"bbeb",x"299b",x"394f",x"2a7d",x"2f3d",x"3949",x"3714",x"35bf",x"bb76",x"27db",x"394a",x"2a4c"),
(x"3004",x"394a",x"3716",x"b86f",x"baa7",x"2604",x"394a",x"2aba",x"3003",x"3949",x"36eb",x"b868",x"baab",x"296a",x"394f",x"2ab4",x"2fa3",x"394d",x"3715",x"a836",x"bbfd",x"294f",x"394a",x"2a84"),
(x"3004",x"394a",x"3716",x"b86f",x"baa7",x"2604",x"394a",x"2aba",x"302c",x"393d",x"3714",x"bb01",x"b7b5",x"2839",x"394a",x"2afc",x"3003",x"3949",x"36eb",x"b868",x"baab",x"296a",x"394f",x"2ab4"),
(x"3036",x"3932",x"3714",x"bbe6",x"310f",x"9bfc",x"394b",x"2b2d",x"3036",x"3933",x"36eb",x"bbf9",x"ad11",x"2511",x"3950",x"2b22",x"302c",x"393d",x"3714",x"bb01",x"b7b5",x"2839",x"394a",x"2afc"),
(x"3026",x"3929",x"3715",x"b928",x"3a1d",x"1553",x"394b",x"2b57",x"3029",x"3929",x"36eb",x"b90c",x"3a34",x"2532",x"3950",x"2b4b",x"3036",x"3932",x"3714",x"bbe6",x"310f",x"9bfc",x"394b",x"2b2d"),
(x"3026",x"3929",x"3715",x"b928",x"3a1d",x"1553",x"394b",x"2b57",x"3006",x"3928",x"3714",x"2fe4",x"3bee",x"28fd",x"394b",x"2b79",x"3029",x"3929",x"36eb",x"b90c",x"3a34",x"2532",x"3950",x"2b4b"),
(x"3006",x"3928",x"3714",x"2fe4",x"3bee",x"28fd",x"394b",x"2b79",x"2fd7",x"392c",x"3711",x"364f",x"3b52",x"2d1b",x"394c",x"2b98",x"3004",x"3929",x"36eb",x"35dd",x"3b6d",x"2be9",x"3950",x"2b72"),
(x"2f89",x"3910",x"3713",x"bbc2",x"b3a4",x"298a",x"394a",x"2c28",x"2f82",x"390f",x"36eb",x"bbf6",x"aa70",x"2d61",x"394f",x"2c30",x"2f73",x"3913",x"3711",x"ba7a",x"b8af",x"283c",x"394b",x"2c1f"),
(x"2fd7",x"392c",x"3711",x"364f",x"3b52",x"2d1b",x"394c",x"2b98",x"2f85",x"392d",x"3710",x"b416",x"3bad",x"2f8b",x"394c",x"2bc3",x"2fdd",x"392e",x"36eb",x"32b2",x"3bc8",x"2e54",x"3950",x"2b90"),
(x"2eec",x"3885",x"3713",x"3583",x"3b63",x"3153",x"3972",x"2c1a",x"2efa",x"3888",x"36eb",x"35e4",x"3b4d",x"31a2",x"3977",x"2c09",x"2f31",x"387c",x"370f",x"3a9c",x"3854",x"30fa",x"3972",x"2c00"),
(x"2f27",x"37cb",x"3715",x"bb82",x"3440",x"330f",x"3992",x"3053",x"2f13",x"3798",x"3715",x"bbc5",x"ab9a",x"3358",x"3993",x"306e",x"2f02",x"37ce",x"36eb",x"bb89",x"3473",x"31fc",x"3997",x"304e"),
(x"2f73",x"3913",x"3711",x"b40c",x"a6bb",x"3bbc",x"394f",x"38c1",x"2f51",x"3919",x"3710",x"a856",x"29ab",x"3bfc",x"3951",x"38bf",x"2fe3",x"390e",x"3718",x"ab65",x"3528",x"3b8f",x"3947",x"38c4"),
(x"3006",x"37c2",x"3715",x"3bd7",x"31f9",x"2c2a",x"398d",x"30c6",x"3008",x"37c9",x"3716",x"38dd",x"ba57",x"297d",x"398d",x"30c9",x"300a",x"37c7",x"36eb",x"3be3",x"ace8",x"30c3",x"3991",x"30d4"),
(x"3015",x"385f",x"3712",x"384e",x"bab0",x"2ec8",x"3920",x"29dd",x"3041",x"386e",x"3710",x"3b6b",x"b5ba",x"2efe",x"3920",x"2a2b",x"301f",x"385d",x"36eb",x"3958",x"b9de",x"2fe4",x"3925",x"29dd"),
(x"2f5e",x"3928",x"3711",x"ba7e",x"3887",x"3089",x"394c",x"2be1",x"2f4e",x"392a",x"36eb",x"baa4",x"3859",x"2fe4",x"3950",x"2be3",x"2f85",x"392d",x"3710",x"b416",x"3bad",x"2f8b",x"394c",x"2bc3"),
(x"2fcc",x"3909",x"3718",x"3be6",x"b09f",x"2baa",x"3998",x"2fd9",x"2fd8",x"3909",x"36eb",x"3be6",x"b08e",x"2c41",x"399b",x"2fcd",x"2fc7",x"38f6",x"3715",x"3bfa",x"2710",x"2c48",x"3996",x"2fc6"),
(x"2f5e",x"3928",x"3711",x"ba7e",x"3887",x"3089",x"394c",x"2be1",x"2f45",x"3921",x"3710",x"bbcc",x"3227",x"2f2f",x"394c",x"2bff",x"2f4e",x"392a",x"36eb",x"baa4",x"3859",x"2fe4",x"3950",x"2be3"),
(x"2f31",x"387c",x"370f",x"3a9c",x"3854",x"30fa",x"3972",x"2c00",x"2f46",x"387d",x"36eb",x"3b7d",x"3521",x"3096",x"3975",x"2bdb",x"2f2d",x"3876",x"370e",x"3b25",x"b70d",x"2d6a",x"3971",x"2bec"),
(x"2e99",x"38b7",x"3714",x"b972",x"39bb",x"30de",x"399d",x"308e",x"2e90",x"38ba",x"36eb",x"b6fe",x"3b25",x"2ea4",x"39a1",x"308f",x"2f21",x"38bd",x"3711",x"b4dc",x"3b97",x"2d60",x"399e",x"3084"),
(x"2f73",x"3913",x"3711",x"ba7a",x"b8af",x"283c",x"394b",x"2c1f",x"2f71",x"3913",x"36eb",x"b9db",x"b96c",x"2c1a",x"394f",x"2c28",x"2f51",x"3919",x"3710",x"bb2f",x"b6d9",x"2e52",x"394b",x"2c11"),
(x"2f75",x"3853",x"3716",x"37e9",x"baf1",x"2aa7",x"391f",x"2974",x"3015",x"385f",x"3712",x"384e",x"bab0",x"2ec8",x"3920",x"29dd",x"2f6d",x"3851",x"36eb",x"3776",x"bb0b",x"2d41",x"3924",x"2965"),
(x"2fd6",x"38f1",x"3715",x"395d",x"39e3",x"2de3",x"3996",x"2fc1",x"2fc7",x"38f6",x"3715",x"3bfa",x"2710",x"2c48",x"3996",x"2fc6",x"2fd9",x"38f3",x"36eb",x"39df",x"3964",x"2d28",x"3999",x"2fb8"),
(x"2efb",x"386d",x"3713",x"3b5b",x"b634",x"2c08",x"396f",x"2bcc",x"2f2d",x"3876",x"370e",x"3b25",x"b70d",x"2d6a",x"3971",x"2bec",x"2f02",x"386c",x"36eb",x"3ad3",x"b822",x"2c4d",x"3973",x"2b9a"),
(x"2fc8",x"381e",x"3716",x"bbff",x"a0b5",x"2138",x"398e",x"3017",x"2f97",x"3809",x"370e",x"bb5f",x"35f1",x"2f4f",x"3991",x"302c",x"2fc6",x"381e",x"36eb",x"bbfe",x"9ea7",x"2828",x"3993",x"3011"),
(x"2f75",x"3853",x"3716",x"37e9",x"baf1",x"2aa7",x"391f",x"2974",x"2f6d",x"3851",x"36eb",x"3776",x"bb0b",x"2d41",x"3924",x"2965",x"2f5c",x"3850",x"3716",x"3bde",x"b1b5",x"2825",x"391f",x"2962"),
(x"3017",x"38e8",x"3719",x"39a6",x"3994",x"2fb1",x"3995",x"2fb4",x"2fd6",x"38f1",x"3715",x"395d",x"39e3",x"2de3",x"3996",x"2fc1",x"3026",x"38e8",x"36eb",x"39ed",x"394b",x"2f45",x"3998",x"2fa6"),
(x"2f3f",x"38c0",x"3711",x"bb12",x"3763",x"2ca3",x"399e",x"3082",x"2f21",x"38bd",x"3711",x"b4dc",x"3b97",x"2d60",x"399e",x"3084",x"2f2b",x"38be",x"36eb",x"b7d8",x"3af6",x"2a35",x"39a1",x"3084"),
(x"2efa",x"386a",x"3713",x"3b09",x"3791",x"2ab5",x"3994",x"30ed",x"2efb",x"386d",x"3713",x"3b5b",x"b634",x"2c08",x"3994",x"30ef",x"2f01",x"386a",x"36eb",x"39e9",x"3955",x"2e31",x"3997",x"30f0"),
(x"2fc8",x"381e",x"3716",x"bbff",x"a0b5",x"2138",x"398e",x"3017",x"2fc6",x"381e",x"36eb",x"bbfe",x"9ea7",x"2828",x"3993",x"3011",x"2f93",x"3832",x"370f",x"bad7",x"b821",x"29e6",x"398e",x"3000"),
(x"2f5c",x"3850",x"3716",x"3bde",x"b1b5",x"2825",x"391f",x"2962",x"2f62",x"3850",x"36eb",x"3b24",x"371c",x"2cde",x"3924",x"295c",x"2f72",x"384b",x"3714",x"39e8",x"3951",x"2f27",x"391f",x"2948"),
(x"3017",x"38e8",x"3719",x"39a6",x"3994",x"2fb1",x"3995",x"2fb4",x"3026",x"38e8",x"36eb",x"39ed",x"394b",x"2f45",x"3998",x"2fa6",x"3017",x"38e6",x"3719",x"3250",x"bbca",x"2f22",x"3995",x"2fb2"),
(x"2f4a",x"38c4",x"3712",x"bbf7",x"a83f",x"2d8f",x"399e",x"3080",x"2f3c",x"38c5",x"36eb",x"bbf8",x"2379",x"2d44",x"39a1",x"3080",x"2f3b",x"38cf",x"3712",x"bb92",x"b509",x"2cb4",x"399e",x"307a"),
(x"2f21",x"3865",x"3710",x"3833",x"3ac7",x"2d1d",x"3994",x"30ea",x"2efa",x"386a",x"3713",x"3b09",x"3791",x"2ab5",x"3994",x"30ed",x"2f01",x"386a",x"36eb",x"39e9",x"3955",x"2e31",x"3997",x"30f0"),
(x"2f3e",x"383c",x"3713",x"b7c2",x"baf3",x"2e28",x"398d",x"2fe4",x"2f93",x"3832",x"370f",x"bad7",x"b821",x"29e6",x"398e",x"3000",x"2f33",x"383a",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3991",x"2fdb"),
(x"2f72",x"384b",x"3714",x"39e8",x"3951",x"2f27",x"391f",x"2948",x"2f83",x"384c",x"36eb",x"397a",x"39b6",x"3099",x"3924",x"2945",x"2fe6",x"383c",x"3717",x"3a77",x"3889",x"310c",x"391f",x"28f0"),
(x"2fe4",x"38e6",x"3718",x"30c5",x"bbe6",x"2ad9",x"3994",x"2fab",x"3017",x"38e6",x"3719",x"3250",x"bbca",x"2f22",x"3995",x"2fb2",x"2fda",x"38e5",x"36eb",x"3b01",x"b745",x"3141",x"3996",x"2f98"),
(x"2f3b",x"38cf",x"3712",x"bb92",x"b509",x"2cb4",x"399e",x"307a",x"2f33",x"38cd",x"36eb",x"bb57",x"b625",x"2e97",x"39a1",x"307b",x"2ec5",x"38f1",x"3711",x"bb70",x"b585",x"3014",x"399f",x"3065"),
(x"2fa3",x"3862",x"3712",x"b2e8",x"3bcb",x"2c10",x"3995",x"30e1",x"2f61",x"3862",x"3713",x"30a8",x"3bea",x"22dc",x"3994",x"30e5",x"2f69",x"3862",x"36eb",x"3046",x"3be8",x"2cb7",x"3997",x"30e7"),
(x"2f3e",x"383c",x"3713",x"b7c2",x"baf3",x"2e28",x"396f",x"2d11",x"2f33",x"383a",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3973",x"2d26",x"2f20",x"383b",x"3712",x"3722",x"bb24",x"2bf2",x"3970",x"2d0b"),
(x"2fe6",x"383c",x"3717",x"3a77",x"3889",x"310c",x"391f",x"28f0",x"3000",x"383d",x"36eb",x"3aff",x"373c",x"3197",x"3925",x"28ea",x"301b",x"3821",x"3713",x"3bc6",x"31be",x"30de",x"391f",x"2878"),
(x"2ec5",x"38f1",x"3711",x"bb70",x"b585",x"3014",x"399f",x"3065",x"2ea7",x"38f3",x"36eb",x"bb99",x"b45f",x"30d6",x"39a2",x"3065",x"2e95",x"3910",x"3711",x"bbe4",x"ad1d",x"308b",x"399f",x"3054"),
(x"3025",x"3872",x"3717",x"bb6f",x"35e4",x"261e",x"3996",x"30d2",x"2fe6",x"3864",x"3711",x"b934",x"3a0d",x"2c16",x"3995",x"30dc",x"3021",x"3872",x"36eb",x"baaf",x"3860",x"2a70",x"3999",x"30d6"),
(x"2f20",x"383b",x"3712",x"3722",x"bb24",x"2bf2",x"3970",x"2d0b",x"2f19",x"3839",x"36eb",x"38ae",x"ba73",x"2d49",x"3974",x"2d1f",x"2ef3",x"3837",x"3711",x"35dd",x"bb65",x"2eae",x"3971",x"2d00"),
(x"3020",x"3806",x"3717",x"3bf0",x"2f10",x"2aec",x"391e",x"2808",x"301b",x"3821",x"3713",x"3bc6",x"31be",x"30de",x"391f",x"2878",x"3025",x"3806",x"36eb",x"3bea",x"2e0a",x"2f10",x"3923",x"27f7"),
(x"2fd8",x"38e4",x"3718",x"3af6",x"37e0",x"2460",x"3956",x"30de",x"2fe4",x"38e6",x"3718",x"30c5",x"bbe6",x"2ad9",x"3956",x"30e0",x"2fda",x"38e5",x"36eb",x"3b01",x"b745",x"3141",x"395b",x"30e0"),
(x"2e95",x"3932",x"3714",x"bbec",x"2d02",x"2f52",x"399f",x"3041",x"2e95",x"3910",x"3711",x"bbe4",x"ad1d",x"308b",x"399f",x"3054",x"2e82",x"3933",x"36eb",x"bbe8",x"2d66",x"3010",x"39a3",x"3041"),
(x"302f",x"3883",x"3715",x"bbfe",x"a412",x"2867",x"3997",x"30ca",x"3025",x"3872",x"3717",x"bb6f",x"35e4",x"261e",x"3996",x"30d2",x"302e",x"3882",x"36eb",x"bbfa",x"2c62",x"2617",x"399a",x"30ce"),
(x"2ef3",x"3837",x"3711",x"35dd",x"bb65",x"2eae",x"3971",x"2d00",x"2efa",x"3835",x"36eb",x"2e28",x"bbe6",x"3005",x"3975",x"2d16",x"2eb1",x"3838",x"3712",x"b5a6",x"bb63",x"30cc",x"3972",x"2cf1"),
(x"3020",x"3806",x"3717",x"3bf0",x"2f10",x"2aec",x"391e",x"2808",x"3025",x"3806",x"36eb",x"3bea",x"2e0a",x"2f10",x"3923",x"27f7",x"3031",x"37df",x"370f",x"3bdd",x"30de",x"2e6c",x"391e",x"2750"),
(x"3006",x"38de",x"3715",x"39d1",x"3974",x"2cc6",x"3956",x"30d4",x"3016",x"38dc",x"36eb",x"3a0e",x"3929",x"2e76",x"395c",x"30d2",x"3022",x"38d3",x"3718",x"3b13",x"3732",x"2fec",x"3956",x"30c7"),
(x"2e95",x"3932",x"3714",x"bbec",x"2d02",x"2f52",x"399f",x"3041",x"2e82",x"3933",x"36eb",x"bbe8",x"2d66",x"3010",x"39a3",x"3041",x"2eb5",x"3942",x"3712",x"bb45",x"3640",x"30a6",x"399f",x"3038"),
(x"2f45",x"3921",x"3710",x"bbcc",x"3227",x"2f2f",x"394c",x"2bff",x"2f51",x"3919",x"3710",x"bb2f",x"b6d9",x"2e52",x"394b",x"2c11",x"2f36",x"3921",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3950",x"2c05"),
(x"302a",x"3899",x"3714",x"bb81",x"b558",x"2da6",x"3998",x"30be",x"302f",x"3883",x"3715",x"bbfe",x"a412",x"2867",x"3997",x"30ca",x"3025",x"3897",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"399b",x"30c3"),
(x"2eb1",x"3838",x"3712",x"b5a6",x"bb63",x"30cc",x"3972",x"2cf1",x"2e9b",x"3835",x"36eb",x"b913",x"ba0d",x"310f",x"3976",x"2d00",x"2e89",x"383f",x"3711",x"bbb2",x"b32f",x"30f4",x"3972",x"2cdf"),
(x"3031",x"37df",x"370f",x"3bdd",x"30de",x"2e6c",x"391e",x"2750",x"303b",x"37e1",x"36eb",x"3be4",x"2adf",x"30ee",x"3923",x"273f",x"302a",x"37d1",x"370d",x"3b0d",x"b70c",x"3169",x"391e",x"2711"),
(x"3022",x"38d3",x"3718",x"3b13",x"3732",x"2fec",x"3956",x"30c7",x"302e",x"38d4",x"36eb",x"3bbf",x"3333",x"2ed0",x"395c",x"30c7",x"3027",x"38cb",x"3712",x"3bf0",x"ac20",x"2e95",x"3957",x"30be"),
(x"2eb5",x"3942",x"3712",x"bb45",x"3640",x"30a6",x"399f",x"3038",x"2ea5",x"3945",x"36eb",x"bab2",x"3834",x"30cf",x"39a3",x"3037",x"2f1a",x"3951",x"3715",x"b93c",x"39e9",x"311d",x"399f",x"302d"),
(x"3008",x"38a8",x"3715",x"ba65",x"b8c1",x"2d9e",x"3999",x"30b5",x"302a",x"3899",x"3714",x"bb81",x"b558",x"2da6",x"3998",x"30be",x"3001",x"38a7",x"36eb",x"bac2",x"b833",x"2e85",x"399c",x"30ba"),
(x"2e89",x"383f",x"3711",x"bbb2",x"b32f",x"30f4",x"3972",x"2cdf",x"2e73",x"383f",x"36eb",x"bbe5",x"2dbc",x"3036",x"3977",x"2ceb",x"2ea4",x"384b",x"3712",x"bae4",x"37c3",x"30c9",x"3973",x"2cc7"),
(x"301d",x"37cb",x"3713",x"3451",x"bbac",x"2d81",x"391d",x"26f7",x"302a",x"37d1",x"370d",x"3b0d",x"b70c",x"3169",x"391e",x"2711",x"3020",x"37c6",x"36eb",x"3571",x"bb6d",x"30cc",x"3922",x"26b4"),
(x"3027",x"38cb",x"3712",x"3bf0",x"ac20",x"2e95",x"3957",x"30be",x"302b",x"38c8",x"36eb",x"3bbf",x"b371",x"2dad",x"395c",x"30bb",x"301e",x"38c8",x"3712",x"3297",x"bbcc",x"2d84",x"3957",x"30ba"),
(x"2f1a",x"3951",x"3715",x"b93c",x"39e9",x"311d",x"399f",x"302d",x"2f13",x"3955",x"36eb",x"b7cb",x"3ae6",x"3068",x"39a2",x"302c",x"2f91",x"3956",x"3715",x"9ef6",x"3bee",x"302a",x"399f",x"3025"),
(x"2fc7",x"38b2",x"3717",x"b939",x"ba0b",x"29e0",x"399a",x"30ae",x"3008",x"38a8",x"3715",x"ba65",x"b8c1",x"2d9e",x"3999",x"30b5",x"2fc1",x"38b1",x"36eb",x"b9cd",x"b979",x"2caa",x"399d",x"30b3"),
(x"2ea4",x"384b",x"3712",x"bae4",x"37c3",x"30c9",x"3973",x"2cc7",x"2e9a",x"384e",x"36eb",x"b902",x"3a23",x"306a",x"3978",x"2ccb",x"2eea",x"384e",x"3713",x"b607",x"3b5e",x"2e4d",x"3973",x"2cb3"),
(x"3008",x"37c9",x"3716",x"38dd",x"ba57",x"297d",x"391d",x"26d4",x"301d",x"37cb",x"3713",x"3451",x"bbac",x"2d81",x"391d",x"26f7",x"300a",x"37c7",x"36eb",x"3be3",x"ace8",x"30c3",x"3922",x"268a"),
(x"3002",x"38c8",x"3717",x"2a07",x"bbfc",x"284d",x"3956",x"30b3",x"301e",x"38c8",x"3712",x"3297",x"bbcc",x"2d84",x"3957",x"30ba",x"2ffe",x"38c7",x"36eb",x"2c58",x"bbf7",x"2bc5",x"395b",x"30ae"),
(x"300a",x"3951",x"3713",x"382e",x"3aba",x"306c",x"399e",x"301c",x"2f91",x"3956",x"3715",x"9ef6",x"3bee",x"302a",x"399f",x"3025",x"3007",x"3955",x"36eb",x"366a",x"3b44",x"2f81",x"39a2",x"301a"),
(x"2fa2",x"38b5",x"3717",x"2c95",x"bbf9",x"2918",x"399a",x"30ac",x"2fc7",x"38b2",x"3717",x"b939",x"ba0b",x"29e0",x"399a",x"30ae",x"2fa3",x"38b4",x"36eb",x"35a6",x"bb74",x"2d53",x"399d",x"30b1"),
(x"2f0a",x"3852",x"3716",x"bac7",x"b83c",x"283f",x"3973",x"2ca8",x"2eea",x"384e",x"3713",x"b607",x"3b5e",x"2e4d",x"3973",x"2cb3",x"2f03",x"3852",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3978",x"2cad"),
(x"2f97",x"3809",x"370e",x"b004",x"271d",x"3bef",x"3949",x"3959",x"2fc8",x"381e",x"3716",x"aadf",x"26b5",x"3bfc",x"3946",x"394d",x"3020",x"3806",x"3717",x"abf6",x"a5ae",x"3bfb",x"393d",x"395a"),
(x"3002",x"38c8",x"3717",x"2a07",x"bbfc",x"284d",x"3956",x"30b3",x"2ffe",x"38c7",x"36eb",x"2c58",x"bbf7",x"2bc5",x"395b",x"30ae",x"2fe7",x"38c7",x"3716",x"38f4",x"ba42",x"2c09",x"3956",x"30af"),
(x"3046",x"3945",x"3715",x"3ae0",x"37cf",x"30d4",x"399d",x"3011",x"300a",x"3951",x"3713",x"382e",x"3aba",x"306c",x"399e",x"301c",x"3051",x"3947",x"36eb",x"39f2",x"3938",x"30b5",x"39a1",x"300e"),
(x"2f79",x"38b1",x"3714",x"39a7",x"b99f",x"2d1e",x"399b",x"30a9",x"2fa2",x"38b5",x"3717",x"2c95",x"bbf9",x"2918",x"399a",x"30ac",x"2fa3",x"38b4",x"36eb",x"35a6",x"bb74",x"2d53",x"399d",x"30b1"),
(x"2f0a",x"3852",x"3716",x"bac7",x"b83c",x"283f",x"3973",x"2ca8",x"2f03",x"3852",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3978",x"2cad",x"2ec3",x"3856",x"3711",x"b8c8",x"ba4e",x"30a8",x"3974",x"2c94"),
(x"2fe7",x"38c7",x"3716",x"38f4",x"ba42",x"2c09",x"3956",x"30af",x"2fea",x"38c5",x"36eb",x"3a76",x"b8ad",x"2cce",x"395b",x"30ab",x"2fda",x"38c4",x"3715",x"3b3f",x"b6b6",x"2b9d",x"3956",x"30ab"),
(x"3061",x"3933",x"3715",x"3bec",x"2be2",x"2fce",x"399c",x"3007",x"3046",x"3945",x"3715",x"3ae0",x"37cf",x"30d4",x"399d",x"3011",x"306a",x"3934",x"36eb",x"3bc4",x"327a",x"3012",x"39a0",x"3004"),
(x"2f4f",x"38ab",x"3714",x"397e",x"b9c5",x"2dbf",x"399b",x"30a5",x"2f4c",x"38a8",x"36eb",x"3976",x"b9cc",x"2dcc",x"399e",x"30a9",x"2f0c",x"38a4",x"3716",x"37d6",x"baf0",x"2d8e",x"399c",x"309f"),
(x"2ec3",x"3856",x"3711",x"b8c8",x"ba4e",x"30a8",x"3974",x"2c94",x"2ea2",x"3855",x"36eb",x"b9ec",x"b92b",x"31e4",x"3979",x"2c94",x"2e71",x"3866",x"370f",x"bb4b",x"b5cc",x"3223",x"3974",x"2c6c"),
(x"3013",x"37ae",x"3712",x"3bcf",x"3081",x"3141",x"398f",x"30be",x"3023",x"37ad",x"36eb",x"3bdb",x"9c67",x"320a",x"3993",x"30c8",x"3008",x"3783",x"370e",x"3b7b",x"b4a9",x"3270",x"3992",x"30ab"),
(x"2fe5",x"38bf",x"3714",x"b879",x"b47b",x"3a3d",x"391d",x"2b97",x"2fda",x"38c4",x"3715",x"3a5f",x"3873",x"3387",x"391d",x"2bab",x"300d",x"38b7",x"3718",x"3ac6",x"37dc",x"3285",x"391d",x"2b6d"),
(x"3058",x"3922",x"3717",x"3b55",x"b5fd",x"307e",x"399b",x"2ffe",x"3061",x"3933",x"3715",x"3bec",x"2be2",x"2fce",x"399c",x"3007",x"3065",x"3921",x"36eb",x"3b6e",x"b575",x"309e",x"399e",x"2ff4"),
(x"2f2f",x"38f9",x"3714",x"b05e",x"a194",x"3bec",x"3953",x"38d0",x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2ec5",x"38f1",x"3711",x"b115",x"a7d5",x"3be4",x"395a",x"38d5"),
(x"2f0c",x"38a4",x"3716",x"37d6",x"baf0",x"2d8e",x"399c",x"309f",x"2f11",x"38a3",x"36eb",x"353f",x"bb87",x"2d28",x"399f",x"30a4",x"2ecb",x"38a3",x"3716",x"a345",x"bbf7",x"2dcc",x"399c",x"309b"),
(x"2e71",x"3866",x"370f",x"bb4b",x"b5cc",x"3223",x"3974",x"2c6c",x"2e56",x"3866",x"36eb",x"bbbc",x"b212",x"3175",x"3979",x"2c6b",x"2e69",x"3879",x"370f",x"bbd3",x"2f46",x"3182",x"3974",x"2c45"),
(x"300d",x"38b7",x"3718",x"3ac6",x"37dc",x"3286",x"391d",x"2b6d",x"3025",x"38b5",x"36eb",x"3afe",x"375c",x"30f4",x"3923",x"2b64",x"3041",x"389f",x"3714",x"3b6b",x"3587",x"3095",x"391f",x"2afc"),
(x"3058",x"3922",x"3717",x"3b55",x"b5fd",x"307e",x"399b",x"2ffe",x"3065",x"3921",x"36eb",x"3b6e",x"b575",x"309e",x"399e",x"2ff4",x"3030",x"3914",x"3711",x"38a4",x"ba69",x"309a",x"399a",x"2fec"),
(x"2ecb",x"38a3",x"3716",x"a345",x"bbf7",x"2dcc",x"399c",x"309b",x"2ec4",x"38a1",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"39a0",x"309f",x"2e97",x"38a6",x"3714",x"b976",x"b9c0",x"3024",x"399d",x"3098"),
(x"2e69",x"3879",x"370f",x"bbd3",x"2f46",x"3182",x"3974",x"2c45",x"2e52",x"387a",x"36eb",x"bb61",x"35a0",x"3119",x"3978",x"2c41",x"2ea1",x"3883",x"370f",x"b891",x"3a72",x"30f5",x"3974",x"2c2c"),
(x"3008",x"3783",x"370e",x"3b7b",x"b4a9",x"3270",x"3992",x"30ab",x"3014",x"377e",x"36eb",x"3ade",x"b7ab",x"31d3",x"3996",x"30b2",x"2fa8",x"3761",x"3712",x"38b5",x"ba3e",x"32bc",x"3994",x"3095"),
(x"3041",x"389f",x"3714",x"3b6b",x"3587",x"3095",x"391f",x"2afc",x"304c",x"389f",x"36eb",x"3bba",x"3376",x"2f14",x"3924",x"2afe",x"3052",x"3886",x"3712",x"3bf0",x"2a00",x"2f46",x"3920",x"2a91"),
(x"2fe3",x"390e",x"3718",x"38ae",x"ba78",x"2b7c",x"3998",x"2fdf",x"3030",x"3914",x"3711",x"38a4",x"ba69",x"309a",x"399a",x"2fec",x"2fed",x"390e",x"36eb",x"360d",x"bb5a",x"2ef3",x"399b",x"2fd2"),
(x"2e97",x"38a6",x"3714",x"b976",x"b9c0",x"3024",x"399d",x"3098",x"2e81",x"38a5",x"36eb",x"bacb",x"b812",x"3064",x"39a0",x"309b",x"2e81",x"38af",x"3712",x"bbe0",x"ae5e",x"30a3",x"399d",x"3093"),
(x"2eec",x"3885",x"3713",x"3583",x"3b63",x"3153",x"3972",x"2c1a",x"2ea1",x"3883",x"370f",x"b891",x"3a72",x"30f5",x"3974",x"2c2c",x"2efa",x"3888",x"36eb",x"35e4",x"3b4d",x"31a2",x"3977",x"2c09"),
(x"2f67",x"3761",x"3716",x"badd",x"b75a",x"334d",x"3994",x"308d",x"2fa8",x"3761",x"3712",x"38b5",x"ba3e",x"32bc",x"3994",x"3095",x"2f52",x"3756",x"36eb",x"b996",x"b95e",x"33ec",x"3999",x"308f"),
(x"3052",x"3886",x"3712",x"3bf0",x"2a00",x"2f46",x"3920",x"2a91",x"305b",x"3885",x"36eb",x"3bef",x"ad09",x"2e69",x"3924",x"2a8f",x"3041",x"386e",x"3710",x"3b6b",x"b5ba",x"2efe",x"3920",x"2a2b"),
(x"2fcc",x"3909",x"3718",x"3be6",x"b09f",x"2baa",x"3998",x"2fd9",x"2fe3",x"390e",x"3718",x"38ae",x"ba78",x"2b7c",x"3998",x"2fdf",x"2fd8",x"3909",x"36eb",x"3be6",x"b08e",x"2c41",x"399b",x"2fcd"),
(x"2e81",x"38af",x"3712",x"bbe0",x"ae5e",x"30a3",x"399d",x"3093",x"2e6a",x"38b0",x"36eb",x"bbcf",x"3174",x"3043",x"39a1",x"3095",x"2e99",x"38b7",x"3714",x"b972",x"39bb",x"30de",x"399d",x"308e"),
(x"2e95",x"3910",x"3711",x"acd1",x"a504",x"3bf9",x"395d",x"38c4",x"2e95",x"3932",x"3714",x"2eb0",x"a8fa",x"3bf3",x"395e",x"38b1",x"2ec4",x"3925",x"3710",x"2828",x"a60a",x"3bfe",x"395a",x"38b8"),
(x"2eb5",x"3942",x"3712",x"a587",x"a08e",x"3bff",x"395c",x"38a8",x"2f06",x"3944",x"3714",x"a8bf",x"ac22",x"3bfa",x"3957",x"38a7",x"2edf",x"393d",x"3712",x"2953",x"a7ae",x"3bfd",x"3959",x"38aa"),
(x"2eb5",x"3942",x"3712",x"a587",x"a08e",x"3bff",x"395c",x"38a8",x"2f1a",x"3951",x"3715",x"a0ea",x"aafd",x"3bfc",x"3956",x"389f",x"2f06",x"3944",x"3714",x"a8bf",x"ac22",x"3bfa",x"3957",x"38a7"),
(x"2f1a",x"3951",x"3715",x"a0ea",x"aafd",x"3bfc",x"3956",x"389f",x"2f91",x"3956",x"3715",x"27e2",x"a9b5",x"3bfc",x"394e",x"389b",x"2f3d",x"3949",x"3714",x"231d",x"ab5f",x"3bfc",x"3953",x"38a3"),
(x"2f91",x"3956",x"3715",x"27e2",x"a9b5",x"3bfc",x"394e",x"389b",x"300a",x"3951",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3946",x"389e",x"2fa3",x"394d",x"3715",x"270a",x"2779",x"3bfe",x"394d",x"38a1"),
(x"300a",x"3951",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3946",x"389e",x"3046",x"3945",x"3715",x"a266",x"1d87",x"3bff",x"393e",x"38a4",x"3004",x"394a",x"3716",x"24bc",x"2ceb",x"3bf9",x"3946",x"38a2"),
(x"3046",x"3945",x"3715",x"a266",x"1d87",x"3bff",x"393e",x"38a4",x"3061",x"3933",x"3715",x"a891",x"27ce",x"3bfd",x"3939",x"38ae",x"302c",x"393d",x"3714",x"a8e0",x"a99e",x"3bfc",x"3941",x"38a9"),
(x"3036",x"3932",x"3714",x"a538",x"29ab",x"3bfd",x"393f",x"38af",x"3061",x"3933",x"3715",x"a891",x"27ce",x"3bfd",x"3939",x"38ae",x"3026",x"3929",x"3715",x"ac67",x"a8a5",x"3bf9",x"3941",x"38b4"),
(x"3058",x"3922",x"3717",x"ad04",x"a793",x"3bf8",x"393a",x"38b8",x"3030",x"3914",x"3711",x"a8d9",x"252b",x"3bfe",x"393f",x"38c0",x"3026",x"3929",x"3715",x"ac67",x"a8a5",x"3bf9",x"3941",x"38b4"),
(x"3006",x"3928",x"3714",x"aa45",x"ab10",x"3bfa",x"3945",x"38b5",x"2f5e",x"3928",x"3711",x"abef",x"28a8",x"3bfa",x"3950",x"38b6",x"2fd7",x"392c",x"3711",x"aa66",x"3318",x"3bca",x"3949",x"38b3"),
(x"2fcc",x"3909",x"3718",x"b420",x"9418",x"3bba",x"3948",x"38c7",x"2f89",x"3910",x"3713",x"b41f",x"2c3a",x"3bb6",x"394d",x"38c4",x"2fe3",x"390e",x"3718",x"ab65",x"3528",x"3b8f",x"3947",x"38c4"),
(x"2fc7",x"38f6",x"3715",x"a7ae",x"24ea",x"3bfe",x"3949",x"38d2",x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2f8e",x"3906",x"3714",x"ade0",x"24c2",x"3bf6",x"394d",x"38c9"),
(x"2f51",x"3919",x"3710",x"a856",x"29ab",x"3bfc",x"3951",x"38bf",x"2f5e",x"3928",x"3711",x"abef",x"28a8",x"3bfa",x"3950",x"38b6",x"3006",x"3928",x"3714",x"aa45",x"ab10",x"3bfa",x"3945",x"38b5"),
(x"2fc7",x"38f6",x"3715",x"a7ae",x"24ea",x"3bfe",x"3949",x"38d2",x"2fd6",x"38f1",x"3715",x"28bf",x"2fda",x"3bef",x"3948",x"38d5",x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7"),
(x"2f8e",x"3906",x"3714",x"bbf3",x"2e23",x"2b27",x"394a",x"2c3b",x"2f6c",x"38ee",x"3718",x"b9e5",x"3968",x"0000",x"3948",x"2c6e",x"2f6c",x"38ee",x"36eb",x"b46a",x"3b91",x"316a",x"394e",x"2c76"),
(x"2f37",x"3a8c",x"36eb",x"bb71",x"b58a",x"2fc3",x"396b",x"2c47",x"2ed7",x"3a9c",x"36eb",x"badb",x"b7e7",x"30ac",x"396c",x"2c1e",x"2f48",x"3a8d",x"3715",x"bac1",x"b812",x"3146",x"3966",x"2c44"),
(x"304f",x"39c2",x"36eb",x"3ba3",x"b452",x"2fdf",x"393f",x"3031",x"302e",x"39b8",x"36eb",x"3bf4",x"2d6d",x"ac2c",x"393c",x"3017",x"3033",x"39b8",x"3715",x"3bf4",x"2da3",x"2b3e",x"3933",x"302a"),
(x"3048",x"39d2",x"3715",x"3bda",x"2e4f",x"312f",x"3937",x"305f",x"3054",x"39d2",x"36eb",x"3b7a",x"3531",x"30a8",x"3942",x"3052",x"304f",x"39c2",x"36eb",x"3ba3",x"b452",x"2fdf",x"393f",x"3031"),
(x"3027",x"39e1",x"3714",x"3a0a",x"3915",x"3126",x"393a",x"3083",x"302b",x"39e5",x"36eb",x"38c7",x"3a49",x"310b",x"3944",x"307f",x"3054",x"39d2",x"36eb",x"3b7a",x"3531",x"30a8",x"3942",x"3052"),
(x"2fca",x"39e9",x"3714",x"3235",x"3bc0",x"30e0",x"393b",x"30aa",x"2fcc",x"39ec",x"36eb",x"23ae",x"3bec",x"306c",x"3945",x"30a6",x"302b",x"39e5",x"36eb",x"38c7",x"3a49",x"310b",x"3944",x"307f"),
(x"2ef2",x"39e6",x"3714",x"b35f",x"3baf",x"30fd",x"393c",x"30e4",x"2ed8",x"39e9",x"36eb",x"b6e0",x"3b1c",x"3118",x"3946",x"30e8",x"2fcc",x"39ec",x"36eb",x"23ae",x"3bec",x"306c",x"3945",x"30a6"),
(x"2e86",x"39db",x"3715",x"ba37",x"38de",x"311d",x"393b",x"310a",x"2e6e",x"39db",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3945",x"3110",x"2ed8",x"39e9",x"36eb",x"b6e0",x"3b1c",x"3118",x"3946",x"30e8"),
(x"2e63",x"39cc",x"3715",x"bbf2",x"2495",x"2f43",x"393a",x"312b",x"2e54",x"39cc",x"36eb",x"bbf7",x"2138",x"2dce",x"3944",x"3132",x"2e6e",x"39db",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3945",x"3110"),
(x"2e6b",x"39be",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3943",x"3150",x"2e54",x"39cc",x"36eb",x"bbf7",x"2138",x"2dce",x"3944",x"3132",x"2e63",x"39cc",x"3715",x"bbf2",x"2495",x"2f43",x"393a",x"312b"),
(x"2e93",x"39b4",x"36eb",x"bbfd",x"212b",x"29e6",x"3942",x"3166",x"2e6b",x"39be",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3943",x"3150",x"2e80",x"39be",x"3715",x"bb87",x"b537",x"2d81",x"3938",x"3149"),
(x"2e6c",x"3981",x"36eb",x"bb9b",x"34d2",x"2ca7",x"393d",x"31d3",x"2e77",x"3981",x"3717",x"bbe8",x"30a2",x"2973",x"3932",x"31ca",x"2e3f",x"397d",x"3714",x"bb74",x"35a7",x"2d5e",x"3933",x"31dc"),
(x"2f22",x"39b7",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38af",x"3208",x"2f13",x"39b7",x"3718",x"3bf1",x"95bc",x"2fb6",x"38bb",x"3207",x"2f16",x"39c0",x"3716",x"3ba5",x"3473",x"2e24",x"38ba",x"31f3"),
(x"2f2a",x"3983",x"36eb",x"3a79",x"3840",x"3401",x"38b0",x"3278",x"2f0c",x"397d",x"3718",x"3a6d",x"3838",x"3468",x"38bb",x"3284",x"2f13",x"39b7",x"3718",x"3bf1",x"95bc",x"2fb6",x"38bb",x"3207"),
(x"306e",x"397f",x"3715",x"3bb4",x"33e8",x"2ed7",x"3926",x"2f62",x"3077",x"3981",x"36eb",x"3bc6",x"328d",x"2f71",x"3930",x"2f41",x"3079",x"3969",x"36eb",x"3409",x"bbbc",x"27db",x"392b",x"2ee7"),
(x"2e24",x"3969",x"36eb",x"b6d0",x"bb39",x"2ab1",x"393a",x"3210",x"2e34",x"397f",x"36eb",x"bb76",x"3593",x"2dee",x"393d",x"31e3",x"2e3f",x"397d",x"3714",x"bb74",x"35a7",x"2d5e",x"3933",x"31dc"),
(x"2fc8",x"39b8",x"36eb",x"bbd3",x"b208",x"2da6",x"38b1",x"313c",x"2fc7",x"39c0",x"36ee",x"bb70",x"358e",x"2fc0",x"38b1",x"314f",x"2fd7",x"39bf",x"3715",x"bb88",x"3531",x"2dc2",x"38bb",x"314f"),
(x"2ffa",x"39c8",x"36ee",x"bb20",x"3725",x"2d51",x"38b2",x"3164",x"3005",x"39ca",x"3717",x"bbd6",x"323b",x"2a8a",x"38bc",x"3169",x"2fd7",x"39bf",x"3715",x"bb88",x"3531",x"2dc2",x"38bb",x"314f"),
(x"2fff",x"39d0",x"36ee",x"bb1d",x"b747",x"2911",x"38b1",x"3176",x"2fff",x"39d2",x"3716",x"baa5",x"b86c",x"2baa",x"38bb",x"317d",x"3005",x"39ca",x"3717",x"bbd6",x"323b",x"2a8a",x"38bc",x"3169"),
(x"2ef6",x"39d0",x"36ee",x"3a41",x"b8fc",x"243f",x"38b0",x"31cc",x"2ef1",x"39d0",x"3714",x"3b3d",x"b6cc",x"26f6",x"38ba",x"31ce",x"2f3a",x"39d8",x"3715",x"3670",x"bb52",x"9df0",x"38ba",x"31b4"),
(x"2fd9",x"39b7",x"3716",x"bbce",x"b2bb",x"2b41",x"38bc",x"313e",x"301e",x"397e",x"3718",x"b98b",x"396b",x"33db",x"38bf",x"30c2",x"3016",x"3985",x"36eb",x"bbe6",x"2cac",x"3077",x"38b3",x"30cc"),
(x"3033",x"39b8",x"3715",x"21a1",x"23fc",x"3bff",x"3974",x"31f5",x"2fd9",x"39b7",x"3716",x"282f",x"2804",x"3bfd",x"396f",x"31f4",x"2fd7",x"39bf",x"3715",x"a8d3",x"a80e",x"3bfd",x"396f",x"31ff"),
(x"303e",x"39c2",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3975",x"3203",x"2fd7",x"39bf",x"3715",x"a8d3",x"a80e",x"3bfd",x"396f",x"31ff",x"3005",x"39ca",x"3717",x"a511",x"281b",x"3bfe",x"3971",x"320c"),
(x"3048",x"39d2",x"3715",x"1e59",x"2bec",x"3bfc",x"3976",x"3218",x"3005",x"39ca",x"3717",x"a511",x"281b",x"3bfe",x"3971",x"320c",x"2fff",x"39d2",x"3716",x"a52b",x"2c98",x"3bfa",x"3971",x"3218"),
(x"3027",x"39e1",x"3714",x"a63f",x"27c1",x"3bfe",x"3973",x"322b",x"2fff",x"39d2",x"3716",x"a52b",x"2c98",x"3bfa",x"3971",x"3218",x"2fc2",x"39d7",x"3713",x"991e",x"9cd0",x"3c00",x"396f",x"321e"),
(x"2fca",x"39e9",x"3714",x"217a",x"a0ea",x"3bff",x"396f",x"3236",x"2fc2",x"39d7",x"3713",x"991e",x"9cd0",x"3c00",x"396f",x"321e",x"2f3a",x"39d8",x"3715",x"1c81",x"1953",x"3c00",x"396a",x"3220"),
(x"2ef2",x"39e6",x"3714",x"9dbc",x"247a",x"3bff",x"3967",x"3232",x"2f3a",x"39d8",x"3715",x"1c81",x"1953",x"3c00",x"396a",x"3220",x"2ef1",x"39d0",x"3714",x"1da1",x"252b",x"3bff",x"3967",x"3215"),
(x"2ef1",x"39d0",x"3714",x"1da1",x"252b",x"3bff",x"3967",x"3215",x"2eed",x"39c9",x"3716",x"a338",x"267a",x"3bff",x"3967",x"320c",x"2e63",x"39cc",x"3715",x"1818",x"26bb",x"3bff",x"3962",x"320f"),
(x"2eed",x"39c9",x"3716",x"a338",x"267a",x"3bff",x"3967",x"320c",x"2f16",x"39c0",x"3716",x"a4b5",x"2b17",x"3bfc",x"3969",x"3200",x"2e80",x"39be",x"3715",x"a64c",x"29dc",x"3bfd",x"3963",x"31fd"),
(x"2e80",x"39be",x"3715",x"a64c",x"29dc",x"3bfd",x"3963",x"31fd",x"2f16",x"39c0",x"3716",x"a4b5",x"2b17",x"3bfc",x"3969",x"3200",x"2f13",x"39b7",x"3718",x"a793",x"2439",x"3bfe",x"3968",x"31f3"),
(x"2e77",x"3981",x"3717",x"a984",x"a0c2",x"3bfd",x"3963",x"31ac",x"2e96",x"39b5",x"3717",x"a7d5",x"236c",x"3bfe",x"3964",x"31f0",x"2f13",x"39b7",x"3718",x"a793",x"2439",x"3bfe",x"3968",x"31f3"),
(x"2ef0",x"39c9",x"36ee",x"3b71",x"35c6",x"2c00",x"38b0",x"31db",x"2eed",x"39c9",x"3716",x"3ba8",x"349f",x"2474",x"38ba",x"31dd",x"2ef1",x"39d0",x"3714",x"3b3d",x"b6cc",x"26f6",x"38ba",x"31ce"),
(x"3033",x"39b8",x"3715",x"3bf4",x"2da3",x"2b3e",x"3933",x"302a",x"302e",x"39b8",x"36eb",x"3bf4",x"2d6d",x"ac2c",x"393c",x"3017",x"3065",x"3981",x"36eb",x"3baa",x"3479",x"2b93",x"3930",x"2f54"),
(x"306e",x"397f",x"3715",x"3bb4",x"33e8",x"2ed7",x"3926",x"2f62",x"3056",x"3980",x"3718",x"3ba4",x"33dc",x"313d",x"3926",x"2f7d",x"3065",x"3981",x"36eb",x"3baa",x"3479",x"2b93",x"3930",x"2f54"),
(x"2f0c",x"397d",x"3718",x"a3ae",x"ac2d",x"3bfb",x"3968",x"31a7",x"301e",x"397e",x"3718",x"224c",x"a379",x"3bff",x"3973",x"31a9",x"3072",x"3969",x"3715",x"2081",x"ad9e",x"3bf8",x"3979",x"318d"),
(x"2fff",x"39d0",x"36ee",x"bb1d",x"b747",x"2911",x"38b1",x"3176",x"2fc4",x"39d8",x"36ee",x"b52c",x"bb8d",x"ac0b",x"38b1",x"318d",x"2fc2",x"39d7",x"3713",x"b46c",x"bbaf",x"a5f6",x"38ba",x"318f"),
(x"2e77",x"3981",x"3717",x"bbe8",x"30a2",x"2973",x"3932",x"31ca",x"2e6c",x"3981",x"36eb",x"bb9b",x"34d2",x"2ca7",x"393d",x"31d3",x"2e93",x"39b4",x"36eb",x"bbfd",x"212b",x"29e6",x"3942",x"3166"),
(x"2f3e",x"39d9",x"36ee",x"3123",x"bbe4",x"a874",x"38b1",x"31b1",x"2f3a",x"39d8",x"3715",x"3670",x"bb52",x"9df0",x"38ba",x"31b4",x"2fc2",x"39d7",x"3713",x"b46c",x"bbaf",x"a5f6",x"38ba",x"318f"),
(x"2f2a",x"3983",x"36eb",x"3a79",x"3840",x"3401",x"38af",x"3089",x"3016",x"3985",x"36eb",x"bbe6",x"2cac",x"3077",x"38b3",x"30cc",x"301e",x"397e",x"3718",x"b98b",x"396b",x"33db",x"38bf",x"30c2"),
(x"2e32",x"396a",x"3714",x"af03",x"bbf3",x"23ef",x"3930",x"3204",x"3072",x"3969",x"3715",x"33c8",x"bbc2",x"235f",x"3921",x"32b2",x"3079",x"3969",x"36eb",x"3409",x"bbbc",x"27db",x"392b",x"32c5"),
(x"2ef0",x"39c9",x"36ee",x"3b71",x"35c6",x"2c00",x"38b0",x"31db",x"2f2c",x"39c2",x"36eb",x"3b82",x"350f",x"3071",x"38af",x"31f1",x"2f16",x"39c0",x"3716",x"3ba5",x"3473",x"2e24",x"38ba",x"31f3"),
(x"2f10",x"3b90",x"370e",x"afd2",x"2717",x"3bef",x"396f",x"3984",x"2f7a",x"3ba1",x"3712",x"b42b",x"2e69",x"3bae",x"3975",x"398f",x"2fbb",x"3ba1",x"3716",x"b0f9",x"a8b2",x"3be5",x"3979",x"398f"),
(x"2fbb",x"3ba1",x"3716",x"3add",x"375a",x"334d",x"396e",x"3097",x"2fd0",x"3ba6",x"36eb",x"3996",x"395f",x"33ec",x"3973",x"309a",x"301b",x"3b86",x"36eb",x"3b99",x"3315",x"330d",x"3973",x"3076"),
(x"2fb0",x"3b06",x"3714",x"2c39",x"29a5",x"3bf9",x"397f",x"3937",x"2fe3",x"3b15",x"3713",x"2da1",x"2f14",x"3beb",x"3982",x"3940",x"3001",x"3b16",x"3712",x"2a69",x"287e",x"3bfc",x"3984",x"3940"),
(x"3017",x"3b1a",x"3711",x"2994",x"2977",x"3bfc",x"3987",x"3943",x"3038",x"3b19",x"3712",x"aa38",x"ad35",x"3bf6",x"398c",x"3942",x"304c",x"3b12",x"3711",x"2481",x"2546",x"3bff",x"398e",x"393e"),
(x"303e",x"3b06",x"3712",x"2a73",x"2a97",x"3bfa",x"398d",x"3938",x"301b",x"3b03",x"3713",x"291b",x"2b55",x"3bfb",x"3988",x"3936",x"3001",x"3b16",x"3712",x"2a69",x"287e",x"3bfc",x"3984",x"3940"),
(x"2ff2",x"3afd",x"3718",x"2e36",x"a153",x"3bf6",x"3984",x"3932",x"300c",x"3aff",x"3716",x"2f15",x"329c",x"3bc6",x"3986",x"3933",x"302f",x"3afb",x"3711",x"2fec",x"ac2c",x"3beb",x"398b",x"3931"),
(x"301b",x"3acc",x"3713",x"2e9a",x"3366",x"3bbd",x"398a",x"3915",x"2ff0",x"3ad5",x"370f",x"ab8d",x"30ae",x"3be6",x"3985",x"391b",x"2ff4",x"3adb",x"370e",x"a6d5",x"25c2",x"3bfe",x"3985",x"391e"),
(x"3013",x"3ae4",x"3713",x"2538",x"ac79",x"3bfa",x"3988",x"3923",x"305c",x"3ad8",x"370f",x"2cd8",x"a71d",x"3bf9",x"3993",x"391e",x"3040",x"3acf",x"370f",x"1df0",x"a631",x"3bff",x"398f",x"3918"),
(x"3013",x"3ae4",x"3713",x"2538",x"ac79",x"3bfa",x"3988",x"3923",x"3014",x"3ae7",x"3713",x"27e9",x"2849",x"3bfd",x"3988",x"3926",x"3058",x"3aeb",x"370f",x"2ec5",x"1a24",x"3bf4",x"3991",x"3928"),
(x"302f",x"3afb",x"3711",x"2fec",x"ac2c",x"3beb",x"398b",x"3931",x"3058",x"3aeb",x"370f",x"2ec5",x"1a24",x"3bf4",x"3991",x"3928",x"3014",x"3ae7",x"3713",x"27e9",x"2849",x"3bfd",x"3988",x"3926"),
(x"3000",x"3aec",x"3710",x"2c5b",x"b0a5",x"3be5",x"3985",x"3928",x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d",x"302f",x"3afb",x"3711",x"2fec",x"ac2c",x"3beb",x"398b",x"3931"),
(x"3000",x"3aec",x"3710",x"2c5b",x"b0a5",x"3be5",x"3985",x"3928",x"2fc1",x"3aef",x"3713",x"a5b5",x"b7de",x"3af6",x"3981",x"392a",x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d"),
(x"2f48",x"3a8d",x"3715",x"26c2",x"ac65",x"3bfa",x"3979",x"38f2",x"2f5a",x"3a9f",x"3717",x"17c8",x"9f93",x"3c00",x"397a",x"38fc",x"2f7f",x"3a9c",x"3717",x"2ff2",x"aa7d",x"3bed",x"397d",x"38fa"),
(x"302b",x"3aae",x"3716",x"2cd8",x"a7e2",x"3bf9",x"398b",x"3905",x"3045",x"3aab",x"3714",x"2860",x"af8d",x"3bf0",x"398e",x"3903",x"3050",x"3aa2",x"3712",x"3163",x"a338",x"3be2",x"3990",x"38fe"),
(x"3044",x"3a9a",x"3714",x"9553",x"ab62",x"3bfc",x"398e",x"38f9",x"3000",x"3a94",x"3711",x"a40b",x"ad5c",x"3bf8",x"3985",x"38f6",x"300a",x"3aad",x"3716",x"a818",x"ad04",x"3bf8",x"3986",x"3904"),
(x"2fa9",x"3aa0",x"3714",x"3036",x"a73e",x"3bed",x"397f",x"38fc",x"2fd3",x"3aa6",x"3714",x"24fd",x"ada9",x"3bf7",x"3982",x"3900",x"3000",x"3a94",x"3711",x"a40b",x"ad5c",x"3bf8",x"3985",x"38f6"),
(x"2fe3",x"3a91",x"3711",x"327d",x"175f",x"3bd5",x"3983",x"38f4",x"2f7f",x"3a9c",x"3717",x"2ff2",x"aa7d",x"3bed",x"397d",x"38fa",x"2fa9",x"3aa0",x"3714",x"3036",x"a73e",x"3bed",x"397f",x"38fc"),
(x"2fe3",x"3a91",x"3711",x"327d",x"175f",x"3bd5",x"3983",x"38f4",x"2fd7",x"3a8d",x"3712",x"2f67",x"a981",x"3bf0",x"3983",x"38f2",x"2f7f",x"3a9c",x"3717",x"2ff2",x"aa7d",x"3bed",x"397d",x"38fa"),
(x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da",x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2fe6",x"3a82",x"3712",x"3146",x"2c91",x"3bde",x"3984",x"38ec"),
(x"2f3d",x"3a6b",x"3718",x"a138",x"ae95",x"3bf4",x"3979",x"38de",x"2f4b",x"3a60",x"3715",x"a8bf",x"afdb",x"3bef",x"397a",x"38d8",x"2ef3",x"3a69",x"3719",x"290e",x"af00",x"3bf2",x"3974",x"38dd"),
(x"2f49",x"3a6d",x"3718",x"ab4f",x"2525",x"3bfc",x"3979",x"38df",x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2fb5",x"3a63",x"3718",x"2e3b",x"1fae",x"3bf6",x"3981",x"38da"),
(x"2f49",x"3a6d",x"3718",x"ab4f",x"2525",x"3bfc",x"3979",x"38df",x"2f16",x"3a73",x"3715",x"ad65",x"ac5b",x"3bf3",x"3976",x"38e3",x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8"),
(x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2f16",x"3a73",x"3715",x"ad65",x"ac5b",x"3bf3",x"3976",x"38e3",x"2ede",x"3a7e",x"3718",x"acf2",x"18ea",x"3bf9",x"3972",x"38e9"),
(x"2ed4",x"3a86",x"3712",x"b59c",x"336a",x"3b42",x"3971",x"38ee",x"2ee4",x"3a89",x"3712",x"b541",x"30ba",x"3b76",x"3972",x"38f0",x"2f1d",x"3a89",x"3717",x"ad2d",x"2ecb",x"3bed",x"3976",x"38ef"),
(x"2f73",x"3a7c",x"3718",x"2bb4",x"28d3",x"3bfa",x"397c",x"38e8",x"2f1d",x"3a89",x"3717",x"ad2d",x"2ecb",x"3bed",x"3976",x"38ef",x"2f3a",x"3a8a",x"3716",x"3009",x"2da6",x"3be7",x"3978",x"38f0"),
(x"2fd7",x"3a8d",x"3712",x"2f67",x"a981",x"3bf0",x"3983",x"38f2",x"2fe6",x"3a82",x"3712",x"3146",x"2c91",x"3bde",x"3984",x"38ec",x"2f3a",x"3a8a",x"3716",x"3009",x"2da6",x"3be7",x"3978",x"38f0"),
(x"2f5a",x"3a9f",x"3717",x"17c8",x"9f93",x"3c00",x"397a",x"38fc",x"2f06",x"3a9a",x"3718",x"2c00",x"290e",x"3bfa",x"3975",x"38f9",x"2f11",x"3aa9",x"3715",x"251e",x"2d06",x"3bf9",x"3975",x"3901"),
(x"2f5a",x"3a9f",x"3717",x"17c8",x"9f93",x"3c00",x"397a",x"38fc",x"2f3c",x"3a92",x"3714",x"257a",x"ae8a",x"3bf4",x"3978",x"38f5",x"2f06",x"3a9a",x"3718",x"2c00",x"290e",x"3bfa",x"3975",x"38f9"),
(x"2f11",x"3aa9",x"3715",x"251e",x"2d06",x"3bf9",x"3975",x"3901",x"2f06",x"3a9a",x"3718",x"2c00",x"290e",x"3bfa",x"3975",x"38f9",x"2e9f",x"3ab2",x"3714",x"975f",x"2c2c",x"3bfb",x"396e",x"3906"),
(x"2ece",x"3ab8",x"3714",x"adba",x"2266",x"3bf7",x"3971",x"390a",x"2e9f",x"3ab2",x"3714",x"975f",x"2c2c",x"3bfb",x"396e",x"3906",x"2e7c",x"3acb",x"3712",x"b106",x"273e",x"3be5",x"396c",x"3915"),
(x"2ec2",x"3ace",x"3715",x"b468",x"247a",x"3bb0",x"3971",x"3916",x"2e7c",x"3acb",x"3712",x"b106",x"273e",x"3be5",x"396c",x"3915",x"2ea0",x"3ae3",x"3710",x"b550",x"2e33",x"3b81",x"396e",x"3922"),
(x"2ed8",x"3adf",x"3717",x"b273",x"2f43",x"3bc8",x"3972",x"3920",x"2ea0",x"3ae3",x"3710",x"b550",x"2e33",x"3b81",x"396e",x"3922",x"2ef8",x"3af2",x"3712",x"ab5f",x"2345",x"3bfc",x"3974",x"392b"),
(x"2f7e",x"3aef",x"3712",x"add2",x"b04b",x"3be4",x"397d",x"3929",x"2fad",x"3afe",x"3716",x"af4d",x"aa5f",x"3bf0",x"397f",x"3932",x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d"),
(x"2f7e",x"3aef",x"3712",x"add2",x"b04b",x"3be4",x"397d",x"3929",x"2ef8",x"3af2",x"3712",x"ab5f",x"2345",x"3bfc",x"3974",x"392b",x"2fad",x"3afe",x"3716",x"af4d",x"aa5f",x"3bf0",x"397f",x"3932"),
(x"2f7e",x"3aef",x"3712",x"add2",x"b04b",x"3be4",x"397d",x"3929",x"2f3c",x"3aed",x"3711",x"2e23",x"2a2e",x"3bf4",x"3978",x"3928",x"2ef8",x"3af2",x"3712",x"ab5f",x"2345",x"3bfc",x"3974",x"392b"),
(x"2ff2",x"3afd",x"3718",x"2e36",x"a153",x"3bf6",x"3984",x"3932",x"2fbb",x"3af4",x"3718",x"2c13",x"b1c5",x"3bda",x"3981",x"392d",x"2fad",x"3afe",x"3716",x"af4d",x"aa5f",x"3bf0",x"397f",x"3932"),
(x"300c",x"3aff",x"3716",x"2f15",x"329c",x"3bc6",x"3986",x"3933",x"2fb0",x"3b06",x"3714",x"2c39",x"29a5",x"3bf9",x"397f",x"3937",x"301b",x"3b03",x"3713",x"291b",x"2b55",x"3bfb",x"3988",x"3936"),
(x"300c",x"3aff",x"3716",x"2f15",x"329c",x"3bc6",x"3986",x"3933",x"2fc5",x"3b01",x"3716",x"2553",x"32c7",x"3bd1",x"3981",x"3934",x"2fb0",x"3b06",x"3714",x"2c39",x"29a5",x"3bf9",x"397f",x"3937"),
(x"2fe3",x"3b15",x"3713",x"2da1",x"2f14",x"3beb",x"3982",x"3940",x"2fb0",x"3b06",x"3714",x"2c39",x"29a5",x"3bf9",x"397f",x"3937",x"2f3b",x"3b15",x"3717",x"30e7",x"3057",x"3bd4",x"3977",x"393f"),
(x"2f8e",x"3b1f",x"370f",x"2edc",x"2cd0",x"3bee",x"397d",x"3945",x"2f3b",x"3b15",x"3717",x"30e7",x"3057",x"3bd4",x"3977",x"393f",x"2eeb",x"3b30",x"3713",x"29b8",x"a6e9",x"3bfd",x"3971",x"394e"),
(x"2ecd",x"3b69",x"370d",x"b809",x"2e09",x"3add",x"396c",x"396e",x"2ee7",x"3b6c",x"3713",x"af9d",x"b907",x"3a25",x"396e",x"3970",x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971"),
(x"3007",x"3b85",x"3715",x"ad56",x"20d0",x"3bf8",x"3980",x"3980",x"2ffb",x"3b6c",x"3715",x"99bc",x"a6cf",x"3bff",x"3980",x"3972",x"2efa",x"3b7a",x"3712",x"a9f0",x"2b1d",x"3bfa",x"396e",x"3978"),
(x"300f",x"3b6a",x"36eb",x"3b89",x"b473",x"31fc",x"3972",x"3059",x"2f92",x"3b47",x"36eb",x"3b4a",x"b677",x"2cf9",x"396f",x"3031",x"2f8b",x"3b48",x"370e",x"3b5f",x"b5f1",x"2f4d",x"396b",x"3036"),
(x"3029",x"3a3e",x"36eb",x"bba1",x"b4cc",x"1f45",x"395f",x"3084",x"3024",x"3a3e",x"3713",x"bba5",x"b497",x"ac28",x"3964",x"3084",x"302f",x"3a2c",x"3710",x"bbfd",x"a997",x"a09b",x"3964",x"3071"),
(x"302f",x"3a2c",x"3710",x"bbfd",x"a997",x"a09b",x"3964",x"3071",x"302e",x"3a20",x"36eb",x"bbf5",x"2e59",x"2467",x"395f",x"3064",x"3029",x"3a3e",x"36eb",x"bba1",x"b4cc",x"1f45",x"395f",x"3084"),
(x"2fb5",x"3a63",x"36eb",x"3469",x"bb91",x"316a",x"395f",x"30b0",x"2fb5",x"3a63",x"3718",x"39e5",x"b968",x"0000",x"3964",x"30b0",x"2ff3",x"3a58",x"3714",x"bb1c",x"b754",x"223f",x"3964",x"30a1"),
(x"2ff3",x"3a58",x"3714",x"bb1c",x"b754",x"223f",x"3964",x"30a1",x"3029",x"3a3e",x"36eb",x"bba1",x"b4cc",x"1f45",x"395f",x"3084",x"2fb5",x"3a63",x"36eb",x"3469",x"bb91",x"316a",x"395f",x"30b0"),
(x"302e",x"3a20",x"36eb",x"bbf5",x"2e59",x"2467",x"395f",x"3064",x"302b",x"3a1c",x"3714",x"bbeb",x"308b",x"98b5",x"3964",x"3061",x"3021",x"3a14",x"3712",x"bb76",x"35c5",x"204d",x"3964",x"3057"),
(x"3021",x"3a14",x"3712",x"bb76",x"35c5",x"204d",x"3964",x"3057",x"301c",x"3a11",x"36eb",x"bab1",x"3862",x"21f0",x"395f",x"3054",x"302e",x"3a20",x"36eb",x"bbf5",x"2e59",x"2467",x"395f",x"3064"),
(x"2fe9",x"3a09",x"36eb",x"b7e1",x"3af5",x"269a",x"395f",x"3046",x"301c",x"3a11",x"36eb",x"bab1",x"3862",x"21f0",x"395f",x"3054",x"300e",x"3a0d",x"3714",x"b95a",x"39f1",x"2032",x"3964",x"304f"),
(x"2f83",x"3a06",x"36eb",x"b03c",x"3beb",x"299b",x"395f",x"3038",x"2fe9",x"3a09",x"36eb",x"b7e1",x"3af5",x"269a",x"395f",x"3046",x"2fe4",x"3a08",x"3714",x"b5bf",x"3b76",x"27db",x"3964",x"3046"),
(x"2f1b",x"3a08",x"36eb",x"3868",x"3aab",x"296a",x"395f",x"302b",x"2f83",x"3a06",x"36eb",x"b03c",x"3beb",x"299b",x"395f",x"3038",x"2f7e",x"3a04",x"3715",x"2836",x"3bfd",x"294f",x"3964",x"3038"),
(x"2ec8",x"3a14",x"3714",x"3b01",x"37b5",x"2839",x"3964",x"301a",x"2ecf",x"3a14",x"36eb",x"3af3",x"37df",x"2b38",x"395f",x"301a",x"2f1b",x"3a08",x"36eb",x"3868",x"3aab",x"296a",x"395f",x"302b"),
(x"2eb5",x"3a1e",x"36eb",x"3bf9",x"2d11",x"2511",x"395f",x"300f",x"2ecf",x"3a14",x"36eb",x"3af3",x"37df",x"2b38",x"395f",x"301a",x"2ec8",x"3a14",x"3714",x"3b01",x"37b5",x"2839",x"3964",x"301a"),
(x"2ecf",x"3a28",x"36eb",x"390c",x"ba34",x"2532",x"395f",x"3005",x"2eb5",x"3a1e",x"36eb",x"3bf9",x"2d11",x"2511",x"395f",x"300f",x"2eb5",x"3a1f",x"3714",x"3be6",x"b10f",x"9bfc",x"3964",x"300d"),
(x"2f14",x"3a29",x"3714",x"afe2",x"bbee",x"28fd",x"3baa",x"3ad9",x"2f19",x"3a28",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3baa",x"3add",x"2ecf",x"3a28",x"36eb",x"390c",x"ba34",x"2532",x"3bad",x"3add"),
(x"2f4a",x"3a25",x"3711",x"b64f",x"bb52",x"2d1b",x"3ba8",x"3ada",x"2f44",x"3a23",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3ba9",x"3ade",x"2f19",x"3a28",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3baa",x"3add"),
(x"2f9f",x"3a42",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b9b",x"3ade",x"2fb1",x"3a3e",x"36eb",x"39db",x"396c",x"2c1a",x"3b9d",x"3ade",x"2faf",x"3a3e",x"3711",x"3a7a",x"38b0",x"283c",x"3b9d",x"3ada"),
(x"2f9c",x"3a24",x"3710",x"3416",x"bbad",x"2f8d",x"3ba5",x"3ada",x"2fa8",x"3a23",x"36eb",x"337e",x"bbba",x"2ef6",x"3ba5",x"3ade",x"2f44",x"3a23",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3ba9",x"3ade"),
(x"3013",x"3ac9",x"36eb",x"b5e4",x"bb4d",x"31a2",x"395a",x"2f00",x"2fdc",x"3ad4",x"36eb",x"bb7d",x"b521",x"3095",x"3957",x"2ef3",x"2ff0",x"3ad5",x"370f",x"ba9c",x"b854",x"30fa",x"3955",x"2f17"),
(x"3007",x"3b85",x"3715",x"3bc5",x"2b9a",x"3358",x"396e",x"3078",x"301b",x"3b86",x"36eb",x"3b99",x"3315",x"330d",x"3973",x"3076",x"300f",x"3b6a",x"36eb",x"3b89",x"b473",x"31fc",x"3972",x"3059"),
(x"2fd1",x"3a38",x"3710",x"2856",x"a9ab",x"3bfc",x"3983",x"38c2",x"2ec0",x"3a3d",x"3711",x"28d9",x"a52b",x"3bfe",x"3971",x"38c3",x"2f3e",x"3a43",x"3718",x"2b65",x"b528",x"3b8f",x"3979",x"38c8"),
(x"2f0d",x"3b6e",x"36eb",x"bbe3",x"2ce8",x"30c3",x"396b",x"30de",x"2efa",x"3b7a",x"3712",x"bbcf",x"b081",x"3141",x"3969",x"30c7",x"2f14",x"3b70",x"3715",x"bbd7",x"b1f9",x"2c2a",x"3967",x"30d0"),
(x"2f0d",x"3b6e",x"36eb",x"bbe3",x"2ce8",x"30c3",x"396b",x"30de",x"2edb",x"3b7b",x"36eb",x"bbdb",x"1c67",x"320a",x"396d",x"30d2",x"2efa",x"3b7a",x"3712",x"bbcf",x"b081",x"3141",x"3969",x"30c7"),
(x"2ea0",x"3ae3",x"3710",x"bb6a",x"35bb",x"2efe",x"3967",x"2b07",x"2e95",x"3ae4",x"36eb",x"bb75",x"35a2",x"2d46",x"396c",x"2b03",x"2ee2",x"3af4",x"36eb",x"b958",x"39de",x"2fe4",x"396b",x"2ab5"),
(x"2fd3",x"3a27",x"36eb",x"3aa4",x"b859",x"2fe5",x"3ba3",x"3ade",x"2fa8",x"3a23",x"36eb",x"337e",x"bbba",x"2ef6",x"3ba5",x"3ade",x"2f9c",x"3a24",x"3710",x"3416",x"bbad",x"2f8d",x"3ba5",x"3ada"),
(x"2f4a",x"3a48",x"36eb",x"bbe6",x"308e",x"2c41",x"3935",x"238d",x"2f4e",x"3a5b",x"36eb",x"bbfa",x"a0a8",x"2cbc",x"3933",x"2258",x"2f5a",x"3a5b",x"3715",x"bbfa",x"a70a",x"2c48",x"392e",x"22c2"),
(x"2fdc",x"3a30",x"3710",x"3bcc",x"b227",x"2f2f",x"3ba1",x"3ada",x"2fec",x"3a30",x"36eb",x"3bf4",x"9ef6",x"2eb6",x"3ba1",x"3ade",x"2fd3",x"3a27",x"36eb",x"3aa4",x"b859",x"2fe5",x"3ba3",x"3ade"),
(x"2fdc",x"3ad4",x"36eb",x"bb7d",x"b521",x"3095",x"3957",x"2ef3",x"2fe5",x"3ada",x"36eb",x"bb19",x"3744",x"2cf7",x"3956",x"2ef0",x"2ff4",x"3adb",x"370e",x"bb25",x"370e",x"2d6a",x"3954",x"2f12"),
(x"3048",x"3a97",x"36eb",x"36fe",x"bb25",x"2ea4",x"3919",x"283d",x"2ff6",x"3a93",x"36eb",x"37d8",x"baf6",x"2a35",x"3918",x"27dd",x"3000",x"3a94",x"3711",x"34dc",x"bb97",x"2d61",x"3913",x"280e"),
(x"2fb1",x"3a3e",x"36eb",x"39db",x"396c",x"2c1a",x"3b9d",x"3ade",x"2fe0",x"3a3a",x"36eb",x"3b02",x"3776",x"2fc8",x"3b9f",x"3ade",x"2fd1",x"3a38",x"3710",x"3b2f",x"36d9",x"2e52",x"3b9f",x"3ada"),
(x"2ef8",x"3af2",x"3712",x"b84e",x"3ab0",x"2ec7",x"3966",x"2ab9",x"2ee2",x"3af4",x"36eb",x"b958",x"39de",x"2fe4",x"396b",x"2ab5",x"2fb4",x"3b00",x"36eb",x"b776",x"3b0b",x"2d41",x"396a",x"2a3e"),
(x"2f5a",x"3a5b",x"3715",x"bbfa",x"a70a",x"2c48",x"392e",x"22c2",x"2f4e",x"3a5b",x"36eb",x"bbfa",x"a0a8",x"2cbc",x"3933",x"2258",x"2f48",x"3a5e",x"36eb",x"b9df",x"b964",x"2d28",x"3933",x"222b"),
(x"2ff4",x"3adb",x"370e",x"bb25",x"370e",x"2d6a",x"3954",x"2f12",x"2fe5",x"3ada",x"36eb",x"bb19",x"3744",x"2cf7",x"3956",x"2ef0",x"300f",x"3ae5",x"36eb",x"bad3",x"3822",x"2c4d",x"3953",x"2ee9"),
(x"2f8b",x"3b48",x"370e",x"3b5f",x"b5f1",x"2f4d",x"396b",x"3036",x"2f92",x"3b47",x"36eb",x"3b4a",x"b677",x"2cf9",x"396f",x"3031",x"2f5b",x"3b33",x"36eb",x"3bfe",x"1e8d",x"2828",x"396e",x"301b"),
(x"2fb4",x"3b00",x"36eb",x"b776",x"3b0b",x"2d41",x"396a",x"2a3e",x"2fc0",x"3b01",x"36eb",x"bb24",x"b71c",x"2cde",x"396a",x"2a35",x"2fc5",x"3b01",x"3716",x"bbde",x"31b5",x"2825",x"3965",x"2a3f"),
(x"2f4b",x"3a60",x"3715",x"b95d",x"b9e3",x"2de3",x"392e",x"2274",x"2f48",x"3a5e",x"36eb",x"b9df",x"b964",x"2d28",x"3933",x"222b",x"2ed5",x"3a69",x"36eb",x"b9ed",x"b94b",x"2f45",x"3932",x"2101"),
(x"2fe5",x"3a8c",x"36eb",x"3bf8",x"a379",x"2d44",x"3930",x"2a7d",x"2fd7",x"3a8d",x"3712",x"3bf7",x"2843",x"2d8f",x"392c",x"2a6d",x"2fe3",x"3a91",x"3711",x"3b12",x"b763",x"2ca3",x"392c",x"2a7d"),
(x"2fe3",x"3a91",x"3711",x"3b12",x"b763",x"2ca3",x"392c",x"2a7d",x"2ff6",x"3a93",x"36eb",x"37d8",x"baf6",x"2a35",x"3930",x"2a9b",x"2fe5",x"3a8c",x"36eb",x"3bf8",x"a379",x"2d44",x"3930",x"2a7d"),
(x"3013",x"3ae4",x"3713",x"bb5b",x"3634",x"2c08",x"3951",x"2f12",x"300f",x"3ae5",x"36eb",x"bad3",x"3822",x"2c4d",x"3953",x"2ee9",x"3010",x"3ae7",x"36eb",x"b9e9",x"b955",x"2e31",x"3952",x"2ee7"),
(x"2f5b",x"3b33",x"36eb",x"3bfe",x"1e8d",x"2828",x"396e",x"301b",x"2f92",x"3b20",x"36eb",x"3ab4",x"3859",x"2a59",x"396d",x"3006",x"2f8e",x"3b1f",x"370f",x"3ad7",x"3821",x"29e6",x"3969",x"300a"),
(x"2fc0",x"3b01",x"36eb",x"bb24",x"b71c",x"2cde",x"3954",x"3138",x"2f9f",x"3b05",x"36eb",x"b97a",x"b9b6",x"309a",x"3955",x"3135",x"2fb0",x"3b06",x"3714",x"b9e8",x"b951",x"2f27",x"3952",x"3123"),
(x"2ed5",x"3a69",x"36eb",x"b9ed",x"b94b",x"2f45",x"3932",x"2101",x"2edf",x"3a6d",x"36eb",x"b2cb",x"3bc1",x"2fc5",x"3932",x"20bd",x"2ef4",x"3a6b",x"3719",x"b250",x"3bca",x"2f22",x"392d",x"2173"),
(x"2fe5",x"3a8c",x"36eb",x"3bf8",x"a379",x"2d44",x"3930",x"2a7d",x"2fee",x"3a84",x"36eb",x"3b57",x"3625",x"2e99",x"3931",x"2a5c",x"2fe6",x"3a82",x"3712",x"3b92",x"3509",x"2cb4",x"392d",x"2a40"),
(x"2fb8",x"3aef",x"36eb",x"b046",x"bbe8",x"2cb7",x"3919",x"2b0c",x"2fc1",x"3aef",x"3713",x"b0a8",x"bbea",x"22dc",x"3914",x"2b18",x"3000",x"3aec",x"3710",x"b833",x"bac7",x"2d1d",x"3915",x"2b3b"),
(x"3000",x"3aec",x"3710",x"b833",x"bac7",x"2d1d",x"3915",x"2b3b",x"3010",x"3ae7",x"36eb",x"b9e9",x"b955",x"2e31",x"391a",x"2b4c",x"2fb8",x"3aef",x"36eb",x"b046",x"bbe8",x"2cb7",x"3919",x"2b0c"),
(x"2f8e",x"3b1f",x"370f",x"3ad7",x"3821",x"29e6",x"3969",x"300a",x"2f92",x"3b20",x"36eb",x"3ab4",x"3859",x"2a59",x"396d",x"3006",x"2fee",x"3b17",x"36eb",x"373f",x"3b1a",x"2d3c",x"396d",x"2fef"),
(x"2f9f",x"3b05",x"36eb",x"b97a",x"b9b6",x"309a",x"3955",x"3135",x"2f20",x"3b14",x"36eb",x"baff",x"b73c",x"3197",x"3959",x"3128",x"2f3b",x"3b15",x"3717",x"ba77",x"b889",x"310c",x"3956",x"3116"),
(x"2ef4",x"3a6b",x"3719",x"b250",x"3bca",x"2f22",x"392d",x"2173",x"2edf",x"3a6d",x"36eb",x"b2cb",x"3bc1",x"2fc5",x"3932",x"20bd",x"2f48",x"3a6c",x"36eb",x"bb01",x"3745",x"3141",x"3930",x"2008"),
(x"2fee",x"3a84",x"36eb",x"3b57",x"3625",x"2e99",x"3931",x"2a5c",x"303d",x"3a5e",x"36eb",x"3b99",x"345f",x"30d6",x"3934",x"29b7",x"302e",x"3a60",x"3711",x"3b70",x"3585",x"3014",x"392f",x"29ac"),
(x"2f42",x"3aeb",x"36eb",x"374a",x"bb15",x"2de4",x"3919",x"2acc",x"2f3c",x"3aed",x"3711",x"3934",x"ba0d",x"2c18",x"3914",x"2ad1",x"2f7e",x"3aef",x"3712",x"32e8",x"bbcb",x"2c10",x"3914",x"2af5"),
(x"2f7e",x"3aef",x"3712",x"32e8",x"bbcb",x"2c10",x"3914",x"2af5",x"2fb8",x"3aef",x"36eb",x"b046",x"bbe8",x"2cb7",x"3919",x"2b0c",x"2f42",x"3aeb",x"36eb",x"374a",x"bb15",x"2de4",x"3919",x"2acc"),
(x"2fee",x"3b17",x"36eb",x"373f",x"3b1a",x"2d3c",x"396d",x"2fef",x"3004",x"3b18",x"36eb",x"b8ae",x"3a73",x"2d49",x"396c",x"2fe8",x"3001",x"3b16",x"3712",x"b721",x"3b24",x"2bf2",x"3968",x"2fef"),
(x"2f20",x"3b14",x"36eb",x"baff",x"b73c",x"3197",x"3959",x"3128",x"2ecb",x"3b30",x"36eb",x"bbbf",x"b113",x"322d",x"395f",x"3114",x"2eeb",x"3b30",x"3713",x"bbc6",x"b1be",x"30de",x"395c",x"3104"),
(x"303d",x"3a5e",x"36eb",x"3b99",x"345f",x"30d6",x"3934",x"29b7",x"3051",x"3a41",x"36eb",x"3be6",x"2c77",x"308b",x"3936",x"293e",x"3046",x"3a41",x"3711",x"3be4",x"2d1d",x"308b",x"3931",x"292a"),
(x"2f3c",x"3aed",x"3711",x"3934",x"ba0d",x"2c18",x"3914",x"2ad1",x"2f42",x"3aeb",x"36eb",x"374a",x"bb15",x"2de4",x"3919",x"2acc",x"2ede",x"3adf",x"36eb",x"3aaf",x"b860",x"2a70",x"3919",x"2a84"),
(x"3004",x"3b18",x"36eb",x"b8ae",x"3a73",x"2d49",x"396c",x"2fe8",x"3014",x"3b1c",x"36eb",x"ae29",x"3be6",x"3005",x"396c",x"2fdc",x"3017",x"3b1a",x"3711",x"b5dd",x"3b65",x"2eae",x"3968",x"2fe1"),
(x"2eeb",x"3b30",x"3713",x"bbc6",x"b1be",x"30de",x"395c",x"3104",x"2ecb",x"3b30",x"36eb",x"bbbf",x"b113",x"322d",x"395f",x"3114",x"2ed7",x"3b4b",x"36eb",x"bbea",x"ae09",x"2f12",x"3964",x"3101"),
(x"2f48",x"3a6c",x"36eb",x"bb01",x"3745",x"3141",x"396a",x"2cb1",x"2f16",x"3a73",x"3715",x"b9d1",x"b974",x"2cc6",x"3966",x"2c96",x"2f49",x"3a6d",x"3718",x"baf5",x"b7e1",x"2460",x"3965",x"2ca9"),
(x"2f48",x"3a6c",x"36eb",x"bb01",x"3745",x"3141",x"396a",x"2cb1",x"2ef5",x"3a75",x"36eb",x"ba0e",x"b929",x"2e78",x"396b",x"2c95",x"2f16",x"3a73",x"3715",x"b9d1",x"b974",x"2cc6",x"3966",x"2c96"),
(x"3046",x"3a41",x"3711",x"3be4",x"2d1d",x"308b",x"3931",x"292a",x"3051",x"3a41",x"36eb",x"3be6",x"2c77",x"308b",x"3936",x"293e",x"304f",x"3a1e",x"36eb",x"3be8",x"ad66",x"3010",x"3938",x"28b0"),
(x"2ed8",x"3adf",x"3717",x"3b6f",x"b5e5",x"261e",x"3913",x"2a83",x"2ede",x"3adf",x"36eb",x"3aaf",x"b860",x"2a70",x"3919",x"2a84",x"2ec6",x"3acf",x"36eb",x"3bfa",x"ac62",x"2617",x"3919",x"2a40"),
(x"3014",x"3b1c",x"36eb",x"ae29",x"3be6",x"3005",x"396c",x"2fdc",x"3043",x"3b1c",x"36eb",x"3913",x"3a0d",x"310f",x"396c",x"2fc3",x"3038",x"3b19",x"3712",x"35a5",x"3b63",x"30cc",x"3967",x"2fd0"),
(x"2ed7",x"3b4b",x"36eb",x"bbea",x"ae09",x"2f12",x"3964",x"3101",x"2eaa",x"3b61",x"36eb",x"bbe4",x"aadf",x"30ee",x"3968",x"30f1",x"2ebe",x"3b62",x"370f",x"bbdd",x"b0de",x"2e6c",x"3965",x"30e2"),
(x"2ef5",x"3a75",x"36eb",x"ba0e",x"b929",x"2e78",x"396b",x"2c95",x"2ec6",x"3a7d",x"36eb",x"bbbf",x"b333",x"2ed2",x"396b",x"2c80",x"2ede",x"3a7e",x"3718",x"bb13",x"b732",x"2fec",x"3966",x"2c7c"),
(x"304f",x"3a1e",x"36eb",x"3be8",x"ad66",x"3010",x"3938",x"28b0",x"303e",x"3a0c",x"36eb",x"3ab2",x"b834",x"30cf",x"3939",x"2865",x"3036",x"3a0f",x"3712",x"3b45",x"b640",x"30a6",x"3934",x"285e"),
(x"2fd1",x"3a38",x"3710",x"3b2f",x"36d9",x"2e52",x"3b9f",x"3ada",x"2fe0",x"3a3a",x"36eb",x"3b02",x"3776",x"2fc8",x"3b9f",x"3ade",x"2fec",x"3a30",x"36eb",x"3bf4",x"9ef6",x"2eb6",x"3ba1",x"3ade"),
(x"2ec2",x"3ace",x"3715",x"3bfe",x"2412",x"2867",x"3914",x"2a3d",x"2ec6",x"3acf",x"36eb",x"3bfa",x"ac62",x"2617",x"3919",x"2a40",x"2ed7",x"3aba",x"36eb",x"3bcf",x"32aa",x"2bc8",x"3919",x"29e8"),
(x"3043",x"3b1c",x"36eb",x"3913",x"3a0d",x"310f",x"396c",x"2fc3",x"3057",x"3b12",x"36eb",x"3be5",x"adbc",x"3036",x"396b",x"2fae",x"304c",x"3b12",x"3711",x"3bb2",x"332f",x"30f4",x"3967",x"2fbd"),
(x"2eaa",x"3b61",x"36eb",x"bbe4",x"aadf",x"30ee",x"3968",x"30f1",x"2eb7",x"3b6c",x"36eb",x"baf6",x"3714",x"32f0",x"396a",x"30e8",x"2ecd",x"3b69",x"370d",x"bb0d",x"370c",x"3169",x"3966",x"30de"),
(x"2ec6",x"3a7d",x"36eb",x"bbbf",x"b333",x"2ed2",x"396b",x"2c80",x"2ecb",x"3a89",x"36eb",x"bbbf",x"3370",x"2dad",x"396c",x"2c68",x"2ed4",x"3a86",x"3712",x"bbf0",x"2c20",x"2e95",x"3967",x"2c6b"),
(x"303e",x"3a0c",x"36eb",x"3ab2",x"b834",x"30cf",x"3939",x"2865",x"3007",x"39fc",x"36eb",x"37cb",x"bae6",x"3068",x"393a",x"280f",x"3003",x"3a00",x"3715",x"393c",x"b9e9",x"311d",x"3934",x"280a"),
(x"2ece",x"3ab8",x"3714",x"3b81",x"3558",x"2da6",x"3914",x"29e0",x"2ed7",x"3aba",x"36eb",x"3bcf",x"32aa",x"2bc8",x"3919",x"29e8",x"2f1f",x"3aaa",x"36eb",x"3ac2",x"3833",x"2e85",x"3919",x"299b"),
(x"3057",x"3b12",x"36eb",x"3be5",x"adbc",x"3036",x"396b",x"2fae",x"3044",x"3b03",x"36eb",x"3902",x"ba23",x"306a",x"3969",x"2f90",x"303e",x"3b06",x"3712",x"3ae4",x"b7c4",x"30c9",x"3965",x"2fa8"),
(x"2ecd",x"3b69",x"370d",x"bb0d",x"370c",x"3169",x"3966",x"30de",x"2eb7",x"3b6c",x"36eb",x"baf6",x"3714",x"32f0",x"396a",x"30e8",x"2ee1",x"3b6e",x"36eb",x"b571",x"3b6d",x"30cc",x"396a",x"30e3"),
(x"2ecb",x"3a89",x"36eb",x"bbbf",x"3370",x"2dad",x"396c",x"2c68",x"2ed6",x"3a8b",x"36eb",x"aeda",x"3bea",x"2e47",x"396c",x"2c62",x"2ee4",x"3a89",x"3712",x"b297",x"3bcc",x"2d84",x"3967",x"2c63"),
(x"3007",x"39fc",x"36eb",x"37cb",x"bae6",x"3068",x"393a",x"280f",x"2f90",x"39f8",x"36eb",x"175f",x"bbf5",x"2e99",x"393a",x"2796",x"2f91",x"39fb",x"3715",x"1ef6",x"bbee",x"302a",x"3935",x"2791"),
(x"2f11",x"3aa9",x"3715",x"3a65",x"38c1",x"2d9e",x"3914",x"2997",x"2f1f",x"3aaa",x"36eb",x"3ac2",x"3833",x"2e85",x"3919",x"299b",x"2f61",x"3aa0",x"36eb",x"39cd",x"3979",x"2caa",x"3919",x"2965"),
(x"3044",x"3b03",x"36eb",x"3902",x"ba23",x"306a",x"3969",x"2f90",x"3017",x"3b01",x"36eb",x"33f1",x"bbbc",x"2b5c",x"3968",x"2f7d",x"301b",x"3b03",x"3713",x"3607",x"bb5e",x"2e4f",x"3964",x"2f98"),
(x"2ee7",x"3b6c",x"3713",x"b451",x"3bac",x"2d81",x"3966",x"30d8",x"2ee1",x"3b6e",x"36eb",x"b571",x"3b6d",x"30cc",x"396a",x"30e3",x"2f0d",x"3b6e",x"36eb",x"bbe3",x"2ce8",x"30c3",x"396b",x"30de"),
(x"2ee4",x"3a89",x"3712",x"b297",x"3bcc",x"2d84",x"3967",x"2c63",x"2ed6",x"3a8b",x"36eb",x"aeda",x"3bea",x"2e47",x"396c",x"2c62",x"2f24",x"3a8a",x"36eb",x"ac58",x"3bf7",x"2bc1",x"396b",x"2c4e"),
(x"2f91",x"39fb",x"3715",x"1ef6",x"bbee",x"302a",x"3935",x"2791",x"2f90",x"39f8",x"36eb",x"175f",x"bbf5",x"2e99",x"393a",x"2796",x"2f13",x"39fc",x"36eb",x"b66a",x"bb44",x"2f81",x"393a",x"270e"),
(x"2f5a",x"3a9f",x"3717",x"3939",x"3a0b",x"29e0",x"3914",x"2960",x"2f61",x"3aa0",x"36eb",x"39cd",x"3979",x"2caa",x"3919",x"2965",x"2f7e",x"3a9d",x"36eb",x"b5a6",x"3b74",x"2d53",x"3919",x"2952"),
(x"301b",x"3b03",x"3713",x"3607",x"bb5e",x"2e4f",x"3964",x"2f98",x"3017",x"3b01",x"36eb",x"33f1",x"bbbc",x"2b5c",x"3968",x"2f7d",x"300f",x"3aff",x"36eb",x"394d",x"39f2",x"2dc5",x"3967",x"2f78"),
(x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971",x"2ffb",x"3b6c",x"3715",x"99bc",x"a6cf",x"3bff",x"3980",x"3972",x"2f8b",x"3b48",x"370e",x"3004",x"a717",x"3bef",x"397b",x"395d"),
(x"2f14",x"3b70",x"3715",x"258e",x"307a",x"3beb",x"3971",x"3973",x"2efa",x"3b7a",x"3712",x"a9f0",x"2b1d",x"3bfa",x"396e",x"3978",x"2ffb",x"3b6c",x"3715",x"99bc",x"a6cf",x"3bff",x"3980",x"3972"),
(x"2ffb",x"3b6c",x"3715",x"99bc",x"a6cf",x"3bff",x"3980",x"3972",x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971",x"2f14",x"3b70",x"3715",x"258e",x"307a",x"3beb",x"3971",x"3973"),
(x"2f8b",x"3b48",x"370e",x"3004",x"a717",x"3bef",x"397b",x"395d",x"2ee1",x"3b4b",x"3717",x"2bf6",x"25ae",x"3bfb",x"396f",x"395d",x"2f10",x"3b6d",x"3716",x"20ea",x"a780",x"3bfe",x"3971",x"3971"),
(x"2f24",x"3a8a",x"36eb",x"ac58",x"3bf7",x"2bc1",x"396b",x"2c4e",x"2f37",x"3a8c",x"36eb",x"bb71",x"b58a",x"2fc3",x"396b",x"2c47",x"2f3a",x"3a8a",x"3716",x"b8f4",x"3a42",x"2c09",x"3966",x"2c4c"),
(x"2f0e",x"3a00",x"3713",x"b82e",x"baba",x"306c",x"3935",x"2702",x"2f13",x"39fc",x"36eb",x"b66a",x"bb44",x"2f81",x"393a",x"270e",x"2e80",x"3a0a",x"36eb",x"b9f2",x"b938",x"30b5",x"393a",x"2650"),
(x"2fd6",x"3aa9",x"36eb",x"b976",x"39cc",x"2dcc",x"391a",x"290f",x"2fd3",x"3aa6",x"3714",x"b97e",x"39c5",x"2dbf",x"3915",x"290e",x"2fa9",x"3aa0",x"3714",x"b9a7",x"399f",x"2d1e",x"3914",x"2930"),
(x"2fa9",x"3aa0",x"3714",x"b9a7",x"399f",x"2d1e",x"3914",x"2930",x"2f7e",x"3a9d",x"36eb",x"b5a6",x"3b74",x"2d53",x"3919",x"2952",x"2fd6",x"3aa9",x"36eb",x"b976",x"39cc",x"2dcc",x"391a",x"290f"),
(x"300f",x"3aff",x"36eb",x"394d",x"39f2",x"2dc5",x"3967",x"2f78",x"303f",x"3afc",x"36eb",x"39ec",x"392b",x"31e5",x"3966",x"2f62",x"302f",x"3afb",x"3711",x"38c8",x"3a4e",x"30a8",x"3962",x"2f7c"),
(x"2e95",x"3a0c",x"3715",x"bae0",x"b7cf",x"30d4",x"3934",x"265f",x"2e80",x"3a0a",x"36eb",x"b9f2",x"b938",x"30b5",x"393a",x"2650",x"2e4e",x"3a1d",x"36eb",x"bbc4",x"b27a",x"3012",x"3939",x"25a9"),
(x"2fd6",x"3aa9",x"36eb",x"b976",x"39cc",x"2dcc",x"391a",x"290f",x"3008",x"3aae",x"36eb",x"b53f",x"3b87",x"2d28",x"391a",x"28e9",x"300a",x"3aad",x"3716",x"b7d6",x"3af0",x"2d8e",x"3915",x"28e1"),
(x"303f",x"3afc",x"36eb",x"39ec",x"392b",x"31e5",x"3966",x"2f62",x"3065",x"3aeb",x"36eb",x"3bbc",x"3212",x"3175",x"3963",x"2f41",x"3058",x"3aeb",x"370f",x"3b4b",x"35cc",x"3223",x"395f",x"2f5b"),
(x"2edb",x"3b7b",x"36eb",x"bbdb",x"1c67",x"320a",x"396d",x"30d2",x"2ef9",x"3b92",x"36eb",x"bade",x"37ab",x"31d3",x"3970",x"30bd",x"2f10",x"3b90",x"370e",x"bb7b",x"34a9",x"3270",x"396c",x"30b5"),
(x"2f48",x"3a8d",x"3715",x"bac1",x"b812",x"3146",x"3966",x"2c44",x"2ed7",x"3a9c",x"36eb",x"badb",x"b7e7",x"30ac",x"396c",x"2c1e",x"2f06",x"3a9a",x"3718",x"bac6",x"b7dc",x"3286",x"3966",x"2c25"),
(x"2e5f",x"3a1e",x"3715",x"bbec",x"abe2",x"2fce",x"3934",x"25be",x"2e4e",x"3a1d",x"36eb",x"bbc4",x"b27a",x"3012",x"3939",x"25a9",x"2e58",x"3a30",x"36eb",x"bb6e",x"3575",x"309e",x"3938",x"250b"),
(x"2ff3",x"3a58",x"3714",x"305e",x"2194",x"3bec",x"3985",x"38d4",x"3046",x"3a41",x"3711",x"2cd1",x"2504",x"3bf9",x"398f",x"38c7",x"3024",x"3a3e",x"3713",x"30f4",x"1987",x"3be7",x"398b",x"38c5"),
(x"2ff3",x"3a58",x"3714",x"305e",x"2194",x"3bec",x"3985",x"38d4",x"302e",x"3a60",x"3711",x"3115",x"27d5",x"3be4",x"398c",x"38d9",x"3046",x"3a41",x"3711",x"2cd1",x"2504",x"3bf9",x"398f",x"38c7"),
(x"3008",x"3aae",x"36eb",x"b53f",x"3b87",x"2d28",x"391a",x"28e9",x"302e",x"3ab0",x"36eb",x"33e5",x"3bb4",x"2ec2",x"391a",x"28c0",x"302b",x"3aae",x"3716",x"2345",x"3bf7",x"2dcc",x"3915",x"28be"),
(x"3065",x"3aeb",x"36eb",x"3bbc",x"3212",x"3175",x"3963",x"2f41",x"3068",x"3ad7",x"36eb",x"3b61",x"b5a0",x"3119",x"395f",x"2f23",x"305c",x"3ad8",x"370f",x"3bd3",x"af46",x"3182",x"395c",x"2f3f"),
(x"2ed7",x"3a9c",x"36eb",x"badb",x"b7e7",x"30ac",x"396c",x"2c1e",x"2e89",x"3ab2",x"36eb",x"bbba",x"b376",x"2f14",x"396c",x"2bd6",x"2e9f",x"3ab2",x"3714",x"bb6b",x"b587",x"3096",x"3967",x"2bd9"),
(x"2e58",x"3a30",x"36eb",x"bb6e",x"3575",x"309e",x"3938",x"250b",x"2ead",x"3a40",x"36eb",x"b884",x"3a69",x"3249",x"3937",x"2473",x"2ec0",x"3a3d",x"3711",x"b8a4",x"3a69",x"309a",x"3932",x"24a5"),
(x"302e",x"3ab0",x"36eb",x"33e5",x"3bb4",x"2ec2",x"391a",x"28c0",x"3050",x"3aac",x"36eb",x"3acb",x"3812",x"3064",x"391a",x"2898",x"3045",x"3aab",x"3714",x"3976",x"39c0",x"3024",x"3915",x"289f"),
(x"3068",x"3ad7",x"36eb",x"3b61",x"b5a0",x"3119",x"395f",x"2f23",x"3042",x"3acb",x"36eb",x"386e",x"ba87",x"313e",x"395d",x"2f0e",x"3040",x"3acf",x"370f",x"3891",x"ba72",x"30f5",x"395a",x"2f2e"),
(x"2ef9",x"3b92",x"36eb",x"bade",x"37ab",x"31d3",x"3970",x"30bd",x"2f7f",x"3ba6",x"36eb",x"b8a6",x"3a54",x"3207",x"3973",x"30a4",x"2f7a",x"3ba1",x"3712",x"b8b5",x"3a3e",x"32bc",x"396e",x"30a0"),
(x"2e89",x"3ab2",x"36eb",x"bbba",x"b376",x"2f14",x"396c",x"2bd6",x"2e6b",x"3acc",x"36eb",x"bbef",x"2d0b",x"2e69",x"396c",x"2b67",x"2e7c",x"3acb",x"3712",x"bbf0",x"aa00",x"2f46",x"3967",x"2b6e"),
(x"2ec0",x"3a3d",x"3711",x"b8a4",x"3a69",x"309a",x"3932",x"24a5",x"2ead",x"3a40",x"36eb",x"b884",x"3a69",x"3249",x"3937",x"2473",x"2f34",x"3a43",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3935",x"23da"),
(x"3050",x"3aac",x"36eb",x"3acb",x"3812",x"3064",x"391a",x"2898",x"305c",x"3aa1",x"36eb",x"3bcf",x"b173",x"3043",x"391a",x"286a",x"3050",x"3aa2",x"3712",x"3be0",x"2e5e",x"30a3",x"3915",x"287a"),
(x"3040",x"3acf",x"370f",x"3891",x"ba72",x"30f5",x"395a",x"2f2e",x"3042",x"3acb",x"36eb",x"386e",x"ba87",x"313e",x"395d",x"2f0e",x"3013",x"3ac9",x"36eb",x"b5e4",x"bb4d",x"31a2",x"395a",x"2f00"),
(x"2f7a",x"3ba1",x"3712",x"b8b5",x"3a3e",x"32bc",x"396e",x"30a0",x"2f7f",x"3ba6",x"36eb",x"b8a6",x"3a54",x"3207",x"3973",x"30a4",x"2fd0",x"3ba6",x"36eb",x"3996",x"395f",x"33ec",x"3973",x"309a"),
(x"2e6b",x"3acc",x"36eb",x"bbef",x"2d0b",x"2e69",x"396c",x"2b67",x"2e95",x"3ae4",x"36eb",x"bb75",x"35a2",x"2d46",x"396c",x"2b03",x"2ea0",x"3ae3",x"3710",x"bb6a",x"35bb",x"2efe",x"3967",x"2b07"),
(x"2f3e",x"3a43",x"3718",x"b8ae",x"3a78",x"2b7c",x"3930",x"242e",x"2f34",x"3a43",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3935",x"23da",x"2f4a",x"3a48",x"36eb",x"bbe6",x"308e",x"2c41",x"3935",x"238d"),
(x"305c",x"3aa1",x"36eb",x"3bcf",x"b173",x"3043",x"391a",x"286a",x"3048",x"3a97",x"36eb",x"36fe",x"bb25",x"2ea4",x"3919",x"283d",x"3044",x"3a9a",x"3714",x"3972",x"b9bb",x"30de",x"3914",x"2857"),
(x"302f",x"3a2c",x"3710",x"a828",x"260a",x"3bfe",x"398d",x"38bb",x"3024",x"3a3e",x"3713",x"30f4",x"1987",x"3be7",x"398b",x"38c5",x"3046",x"3a41",x"3711",x"2cd1",x"2504",x"3bf9",x"398f",x"38c7"),
(x"3046",x"3a1f",x"3714",x"aeb0",x"28fa",x"3bf3",x"3990",x"38b4",x"302b",x"3a1c",x"3714",x"a946",x"1ffc",x"3bfe",x"398d",x"38b3",x"302f",x"3a2c",x"3710",x"a828",x"260a",x"3bfe",x"398d",x"38bb"),
(x"3036",x"3a0f",x"3712",x"2587",x"208e",x"3bff",x"398e",x"38ab",x"302b",x"3a1c",x"3714",x"a946",x"1ffc",x"3bfe",x"398d",x"38b3",x"3046",x"3a1f",x"3714",x"aeb0",x"28fa",x"3bf3",x"3990",x"38b4"),
(x"3036",x"3a0f",x"3712",x"2587",x"208e",x"3bff",x"398e",x"38ab",x"3021",x"3a14",x"3712",x"a953",x"27ae",x"3bfd",x"398b",x"38ae",x"302b",x"3a1c",x"3714",x"a946",x"1ffc",x"3bfe",x"398d",x"38b3"),
(x"3003",x"3a00",x"3715",x"20ea",x"2afd",x"3bfc",x"3988",x"38a2",x"2fe4",x"3a08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3986",x"38a7",x"300e",x"3a0d",x"3714",x"28bf",x"2c22",x"3bfa",x"3989",x"38aa"),
(x"2f91",x"39fb",x"3715",x"a7e2",x"29b2",x"3bfc",x"3980",x"389f",x"2f7e",x"3a04",x"3715",x"a70a",x"a779",x"3bfe",x"397f",x"38a4",x"2fe4",x"3a08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3986",x"38a7"),
(x"2f0e",x"3a00",x"3713",x"ab1d",x"aee4",x"3bf0",x"3978",x"38a1",x"2f19",x"3a07",x"3716",x"a4bc",x"aceb",x"3bf9",x"3978",x"38a5",x"2f7e",x"3a04",x"3715",x"a70a",x"a779",x"3bfe",x"397f",x"38a4"),
(x"2e95",x"3a0c",x"3715",x"2266",x"9d87",x"3bff",x"3970",x"38a8",x"2ec8",x"3a14",x"3714",x"28e0",x"299e",x"3bfc",x"3973",x"38ac",x"2f19",x"3a07",x"3716",x"a4bc",x"aceb",x"3bf9",x"3978",x"38a5"),
(x"2e5f",x"3a1e",x"3715",x"2891",x"a7ce",x"3bfd",x"396c",x"38b2",x"2eb5",x"3a1f",x"3714",x"2538",x"a9ab",x"3bfd",x"3971",x"38b2",x"2ec8",x"3a14",x"3714",x"28e0",x"299e",x"3bfc",x"3973",x"38ac"),
(x"2e5f",x"3a1e",x"3715",x"2891",x"a7ce",x"3bfd",x"396c",x"38b2",x"2e70",x"3a2f",x"3717",x"2d06",x"2793",x"3bf8",x"396c",x"38bb",x"2ed5",x"3a28",x"3715",x"2c67",x"28a5",x"3bf9",x"3973",x"38b8"),
(x"2ec0",x"3a3d",x"3711",x"28d9",x"a52b",x"3bfe",x"3971",x"38c3",x"2f14",x"3a29",x"3714",x"2a45",x"2b10",x"3bfa",x"3977",x"38b8",x"2ed5",x"3a28",x"3715",x"2c67",x"28a5",x"3bf9",x"3973",x"38b8"),
(x"2fc4",x"3a29",x"3711",x"2bef",x"a8a8",x"3bfa",x"3982",x"38b9",x"2f9c",x"3a24",x"3710",x"2352",x"ae80",x"3bf5",x"3980",x"38b6",x"2f4a",x"3a25",x"3711",x"2a66",x"b319",x"3bca",x"397b",x"38b6"),
(x"2f99",x"3a42",x"3713",x"341f",x"ac3a",x"3bb6",x"397f",x"38c7",x"2faf",x"3a3e",x"3711",x"340c",x"26c2",x"3bbc",x"3981",x"38c5",x"2f3e",x"3a43",x"3718",x"2b65",x"b528",x"3b8f",x"3979",x"38c8"),
(x"2f94",x"3a4b",x"3714",x"2de0",x"a4c2",x"3bf6",x"397f",x"38cc",x"2f55",x"3a48",x"3718",x"3420",x"1418",x"3bba",x"397a",x"38cb",x"2f5a",x"3a5b",x"3715",x"27ae",x"a4f0",x"3bfe",x"397b",x"38d6"),
(x"2f94",x"3a4b",x"3714",x"2de0",x"a4c2",x"3bf6",x"397f",x"38cc",x"2f99",x"3a42",x"3713",x"341f",x"ac3a",x"3bb6",x"397f",x"38c7",x"2f55",x"3a48",x"3718",x"3420",x"1418",x"3bba",x"397a",x"38cb"),
(x"2fc4",x"3a29",x"3711",x"2bef",x"a8a8",x"3bfa",x"3982",x"38b9",x"2fd1",x"3a38",x"3710",x"2856",x"a9ab",x"3bfc",x"3983",x"38c2",x"2fdc",x"3a30",x"3710",x"2a8d",x"2973",x"3bfb",x"3984",x"38bd"),
(x"2f14",x"3a29",x"3714",x"2a45",x"2b10",x"3bfa",x"3977",x"38b8",x"2ec0",x"3a3d",x"3711",x"28d9",x"a52b",x"3bfe",x"3971",x"38c3",x"2fd1",x"3a38",x"3710",x"2856",x"a9ab",x"3bfc",x"3983",x"38c2"),
(x"301e",x"397e",x"3718",x"224c",x"a379",x"3bff",x"3973",x"31a9",x"2fd9",x"39b7",x"3716",x"282f",x"2804",x"3bfd",x"396f",x"31f4",x"3033",x"39b8",x"3715",x"21a1",x"23fc",x"3bff",x"3974",x"31f5"),
(x"2f9f",x"3a42",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b9b",x"3ade",x"2f99",x"3a42",x"3713",x"3bc2",x"33a4",x"298a",x"3b9c",x"3ad9",x"2f94",x"3a4b",x"3714",x"3bf3",x"ae23",x"2b27",x"3b9a",x"3ad9"),
(x"2f94",x"3a4b",x"3714",x"3bf3",x"ae23",x"2b27",x"3b9a",x"3ad9",x"2fb5",x"3a63",x"36eb",x"3469",x"bb91",x"316a",x"3b93",x"3add",x"2f9f",x"3a42",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b9b",x"3ade"),
(x"3008",x"3783",x"370e",x"2fd2",x"a717",x"3bef",x"393d",x"3981",x"2fa8",x"3761",x"3712",x"342b",x"ae69",x"3bae",x"3943",x"398b",x"2f67",x"3761",x"3716",x"30f9",x"28b2",x"3be5",x"3947",x"398c"),
(x"2f67",x"3761",x"3716",x"badd",x"b75a",x"334d",x"3994",x"308d",x"2f52",x"3756",x"36eb",x"b996",x"b95e",x"33ec",x"3999",x"308f",x"2eeb",x"3797",x"36eb",x"bb99",x"b315",x"330d",x"3998",x"306b"),
(x"2f72",x"384b",x"3714",x"ac39",x"a9a5",x"3bf9",x"394d",x"3934",x"2f3e",x"383c",x"3713",x"ada3",x"af14",x"3beb",x"3950",x"393c",x"2f20",x"383b",x"3712",x"aa69",x"a87e",x"3bfc",x"3952",x"393d"),
(x"2ef3",x"3837",x"3711",x"a994",x"a977",x"3bfc",x"3955",x"393f",x"2eb1",x"3838",x"3712",x"2a38",x"2d35",x"3bf6",x"3959",x"393f",x"2e89",x"383f",x"3711",x"a481",x"a546",x"3bff",x"395c",x"393b"),
(x"2ea4",x"384b",x"3712",x"aa73",x"aa97",x"3bfa",x"395b",x"3934",x"2eea",x"384e",x"3713",x"a91b",x"ab55",x"3bfb",x"3956",x"3932",x"2f20",x"383b",x"3712",x"aa69",x"a87e",x"3bfc",x"3952",x"393d"),
(x"2f2f",x"3854",x"3718",x"ae36",x"2153",x"3bf6",x"3952",x"392e",x"2f0a",x"3852",x"3716",x"af15",x"b29c",x"3bc7",x"3954",x"3930",x"2ec3",x"3856",x"3711",x"afec",x"2c2c",x"3beb",x"3959",x"392e"),
(x"2eec",x"3885",x"3713",x"ae9c",x"b367",x"3bbd",x"3958",x"3912",x"2f31",x"387c",x"370f",x"2b8a",x"b0af",x"3be6",x"3953",x"3917",x"2f2d",x"3876",x"370e",x"26d5",x"a5c2",x"3bfe",x"3953",x"391a"),
(x"2efb",x"386d",x"3713",x"a538",x"2c79",x"3bfa",x"3956",x"3920",x"2e69",x"3879",x"370f",x"acd8",x"271d",x"3bf9",x"3960",x"391a",x"2ea1",x"3883",x"370f",x"9df0",x"2631",x"3bff",x"395d",x"3914"),
(x"2efb",x"386d",x"3713",x"a538",x"2c79",x"3bfa",x"3956",x"3920",x"2efa",x"386a",x"3713",x"a7ef",x"a849",x"3bfd",x"3956",x"3922",x"2e71",x"3866",x"370f",x"aec5",x"9a24",x"3bf4",x"395f",x"3925"),
(x"2ec3",x"3856",x"3711",x"afec",x"2c2c",x"3beb",x"3959",x"392e",x"2e71",x"3866",x"370f",x"aec5",x"9a24",x"3bf4",x"395f",x"3925",x"2efa",x"386a",x"3713",x"a7ef",x"a849",x"3bfd",x"3956",x"3922"),
(x"2f21",x"3865",x"3710",x"ac5b",x"30a5",x"3be5",x"3953",x"3925",x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929",x"2ec3",x"3856",x"3711",x"afec",x"2c2c",x"3beb",x"3959",x"392e"),
(x"2f21",x"3865",x"3710",x"ac5b",x"30a5",x"3be5",x"3953",x"3925",x"2f61",x"3862",x"3713",x"25b5",x"37de",x"3af6",x"394f",x"3926",x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929"),
(x"2fda",x"38c4",x"3715",x"a6c2",x"2c63",x"3bfa",x"3947",x"38ee",x"2fc7",x"38b2",x"3717",x"97c8",x"1f79",x"3c00",x"3948",x"38f8",x"2fa2",x"38b5",x"3717",x"aff2",x"2a7a",x"3bed",x"394b",x"38f7"),
(x"2ecb",x"38a3",x"3716",x"acd8",x"27e2",x"3bf9",x"3959",x"3901",x"2e97",x"38a6",x"3714",x"a860",x"2f8b",x"3bf0",x"395c",x"38ff",x"2e81",x"38af",x"3712",x"b162",x"2345",x"3be2",x"395e",x"38fb"),
(x"2e99",x"38b7",x"3714",x"1553",x"2b62",x"3bfc",x"395c",x"38f6",x"2f21",x"38bd",x"3711",x"240b",x"2d5c",x"3bf8",x"3953",x"38f2",x"2f0c",x"38a4",x"3716",x"2818",x"2d04",x"3bf8",x"3954",x"3900"),
(x"2f79",x"38b1",x"3714",x"b036",x"273e",x"3bed",x"394d",x"38f9",x"2f4f",x"38ab",x"3714",x"a4fd",x"2da9",x"3bf7",x"3950",x"38fd",x"2f21",x"38bd",x"3711",x"240b",x"2d5c",x"3bf8",x"3953",x"38f2"),
(x"2f3f",x"38c0",x"3711",x"b27d",x"975f",x"3bd5",x"3951",x"38f1",x"2fa2",x"38b5",x"3717",x"aff2",x"2a7a",x"3bed",x"394b",x"38f7",x"2f79",x"38b1",x"3714",x"b036",x"273e",x"3bed",x"394d",x"38f9"),
(x"2f3f",x"38c0",x"3711",x"b27d",x"975f",x"3bd5",x"3951",x"38f1",x"2f4a",x"38c4",x"3712",x"af67",x"2981",x"3bf0",x"3950",x"38ef",x"2fa2",x"38b5",x"3717",x"aff2",x"2a7a",x"3bed",x"394b",x"38f7"),
(x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7",x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"2f3b",x"38cf",x"3712",x"b146",x"ac91",x"3bde",x"3952",x"38e8"),
(x"2fe4",x"38e6",x"3718",x"2138",x"2e95",x"3bf4",x"3947",x"38db",x"2fd6",x"38f1",x"3715",x"28bf",x"2fda",x"3bef",x"3948",x"38d5",x"3017",x"38e8",x"3719",x"a90e",x"2f00",x"3bf2",x"3942",x"38da"),
(x"2fd8",x"38e4",x"3718",x"2b4f",x"a525",x"3bfc",x"3947",x"38dc",x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"2f6c",x"38ee",x"3718",x"ae3b",x"9fae",x"3bf6",x"394e",x"38d7"),
(x"2fd8",x"38e4",x"3718",x"2b4f",x"a525",x"3bfc",x"3947",x"38dc",x"3006",x"38de",x"3715",x"2d65",x"2c5a",x"3bf3",x"3944",x"38e0",x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5"),
(x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"3006",x"38de",x"3715",x"2d65",x"2c5a",x"3bf3",x"3944",x"38e0",x"3022",x"38d3",x"3718",x"2cf2",x"991e",x"3bf9",x"3940",x"38e5"),
(x"3027",x"38cb",x"3712",x"359c",x"b36a",x"3b42",x"393f",x"38ea",x"301e",x"38c8",x"3712",x"3541",x"b0b9",x"3b76",x"3940",x"38ec",x"3002",x"38c8",x"3717",x"2d2d",x"aecd",x"3bed",x"3944",x"38ec"),
(x"2faf",x"38d5",x"3718",x"abb4",x"a8d3",x"3bfa",x"394a",x"38e5",x"3002",x"38c8",x"3717",x"2d2d",x"aecd",x"3bed",x"3944",x"38ec",x"2fe7",x"38c7",x"3716",x"b009",x"ada6",x"3be7",x"3946",x"38ec"),
(x"2f4a",x"38c4",x"3712",x"af67",x"2981",x"3bf0",x"3950",x"38ef",x"2f3b",x"38cf",x"3712",x"b146",x"ac91",x"3bde",x"3952",x"38e8",x"2fe7",x"38c7",x"3716",x"b009",x"ada6",x"3be7",x"3946",x"38ec"),
(x"2fc7",x"38b2",x"3717",x"97c8",x"1f79",x"3c00",x"3948",x"38f8",x"300d",x"38b7",x"3718",x"ac00",x"a911",x"3bfa",x"3943",x"38f5",x"3008",x"38a8",x"3715",x"a51e",x"ad06",x"3bf9",x"3943",x"38fe"),
(x"2fc7",x"38b2",x"3717",x"97c8",x"1f79",x"3c00",x"3948",x"38f8",x"2fe5",x"38bf",x"3714",x"a581",x"2e8a",x"3bf4",x"3946",x"38f1",x"300d",x"38b7",x"3718",x"ac00",x"a911",x"3bfa",x"3943",x"38f5"),
(x"3008",x"38a8",x"3715",x"a51e",x"ad06",x"3bf9",x"3943",x"38fe",x"300d",x"38b7",x"3718",x"ac00",x"a911",x"3bfa",x"3943",x"38f5",x"3041",x"389f",x"3714",x"175f",x"ac2c",x"3bfb",x"393c",x"3903"),
(x"302a",x"3899",x"3714",x"2dba",x"a266",x"3bf7",x"393f",x"3906",x"3041",x"389f",x"3714",x"175f",x"ac2c",x"3bfb",x"393c",x"3903",x"3052",x"3886",x"3712",x"3106",x"a738",x"3be5",x"393a",x"3911"),
(x"302f",x"3883",x"3715",x"3468",x"a47a",x"3bb0",x"393e",x"3913",x"3052",x"3886",x"3712",x"3106",x"a738",x"3be5",x"393a",x"3911",x"3041",x"386e",x"3710",x"3550",x"ae33",x"3b81",x"393c",x"391f"),
(x"3025",x"3872",x"3717",x"3273",x"af43",x"3bc8",x"3940",x"391c",x"3041",x"386e",x"3710",x"3550",x"ae33",x"3b81",x"393c",x"391f",x"3015",x"385f",x"3712",x"2b5f",x"a345",x"3bfc",x"3942",x"3927"),
(x"2fa3",x"3862",x"3712",x"2dd2",x"304b",x"3be4",x"394b",x"3926",x"2f75",x"3853",x"3716",x"2f4d",x"2a5f",x"3bf0",x"394d",x"392f",x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929"),
(x"2fa3",x"3862",x"3712",x"2dd2",x"304b",x"3be4",x"394b",x"3926",x"3015",x"385f",x"3712",x"2b5f",x"a345",x"3bfc",x"3942",x"3927",x"2f75",x"3853",x"3716",x"2f4d",x"2a5f",x"3bf0",x"394d",x"392f"),
(x"2fa3",x"3862",x"3712",x"2dd2",x"304b",x"3be4",x"394b",x"3926",x"2fe6",x"3864",x"3711",x"ae24",x"aa2e",x"3bf4",x"3946",x"3924",x"3015",x"385f",x"3712",x"2b5f",x"a345",x"3bfc",x"3942",x"3927"),
(x"2f2f",x"3854",x"3718",x"ae36",x"2153",x"3bf6",x"3952",x"392e",x"2f67",x"385d",x"3718",x"ac13",x"31c5",x"3bda",x"394f",x"3929",x"2f75",x"3853",x"3716",x"2f4d",x"2a5f",x"3bf0",x"394d",x"392f"),
(x"2f0a",x"3852",x"3716",x"af15",x"b29c",x"3bc7",x"3954",x"3930",x"2f72",x"384b",x"3714",x"ac39",x"a9a5",x"3bf9",x"394d",x"3934",x"2eea",x"384e",x"3713",x"a91b",x"ab55",x"3bfb",x"3956",x"3932"),
(x"2f0a",x"3852",x"3716",x"af15",x"b29c",x"3bc7",x"3954",x"3930",x"2f5c",x"3850",x"3716",x"a559",x"b2c7",x"3bd1",x"394f",x"3931",x"2f72",x"384b",x"3714",x"ac39",x"a9a5",x"3bf9",x"394d",x"3934"),
(x"2f3e",x"383c",x"3713",x"ada3",x"af14",x"3beb",x"3950",x"393c",x"2f72",x"384b",x"3714",x"ac39",x"a9a5",x"3bf9",x"394d",x"3934",x"2fe6",x"383c",x"3717",x"b0e7",x"b057",x"3bd4",x"3945",x"393c"),
(x"2f93",x"3832",x"370f",x"aedc",x"acd0",x"3bee",x"394b",x"3942",x"2fe6",x"383c",x"3717",x"b0e7",x"b057",x"3bd4",x"3945",x"393c",x"301b",x"3821",x"3713",x"a9b8",x"26e9",x"3bfd",x"393f",x"394b"),
(x"302a",x"37d1",x"370d",x"3809",x"ae09",x"3add",x"393a",x"396b",x"301d",x"37cb",x"3713",x"2f9f",x"3907",x"3a25",x"393c",x"396d",x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d"),
(x"2f13",x"3798",x"3715",x"2d56",x"a0d0",x"3bf8",x"394e",x"397d",x"2f27",x"37cb",x"3715",x"19bc",x"26cf",x"3bff",x"394e",x"396e",x"3013",x"37ae",x"3712",x"29f0",x"ab1d",x"3bfa",x"393c",x"3975"),
(x"2f02",x"37ce",x"36eb",x"bb89",x"3473",x"31fc",x"3997",x"304e",x"2f8f",x"380a",x"36eb",x"bb4a",x"3677",x"2cfa",x"3995",x"3026",x"2f97",x"3809",x"370e",x"bb5f",x"35f1",x"2f4f",x"3991",x"302c"),
(x"2ece",x"3913",x"36eb",x"3ba1",x"34cc",x"1f45",x"394e",x"2951",x"2ed8",x"3913",x"3713",x"3ba5",x"3497",x"ac28",x"3949",x"2954",x"2ec4",x"3925",x"3710",x"3bfd",x"2997",x"a09b",x"394a",x"29a0"),
(x"2ec4",x"3925",x"3710",x"3bfd",x"2997",x"a09b",x"394a",x"29a0",x"2ec5",x"3931",x"36eb",x"3bf5",x"ae59",x"2467",x"394f",x"29ce",x"2ece",x"3913",x"36eb",x"3ba1",x"34cc",x"1f45",x"394e",x"2951"),
(x"2f6c",x"38ee",x"36eb",x"b46a",x"3b91",x"316a",x"394e",x"28a1",x"2f6c",x"38ee",x"3718",x"b9e5",x"3968",x"0000",x"3948",x"28a4",x"2f2f",x"38f9",x"3714",x"3b1c",x"3754",x"223f",x"3949",x"28de"),
(x"2f2f",x"38f9",x"3714",x"3b1c",x"3754",x"223f",x"3949",x"28de",x"2ece",x"3913",x"36eb",x"3ba1",x"34cc",x"1f45",x"394e",x"2951",x"2f6c",x"38ee",x"36eb",x"b46a",x"3b91",x"316a",x"394e",x"28a1"),
(x"2ec5",x"3931",x"36eb",x"3bf5",x"ae59",x"2467",x"394f",x"29ce",x"2eca",x"3935",x"3714",x"3beb",x"b08a",x"98ea",x"394a",x"29e1",x"2edf",x"393d",x"3712",x"3b76",x"b5c5",x"204d",x"394a",x"2a06"),
(x"2edf",x"393d",x"3712",x"3b76",x"b5c5",x"204d",x"394a",x"2a06",x"2ee8",x"3940",x"36eb",x"3ab1",x"b862",x"21f0",x"394f",x"2a10",x"2ec5",x"3931",x"36eb",x"3bf5",x"ae59",x"2467",x"394f",x"29ce"),
(x"2f38",x"3948",x"36eb",x"37e1",x"baf5",x"269a",x"394f",x"2a46",x"2ee8",x"3940",x"36eb",x"3ab1",x"b862",x"21f0",x"394f",x"2a10",x"2f06",x"3944",x"3714",x"395a",x"b9f1",x"2032",x"394a",x"2a28"),
(x"2f9e",x"394c",x"36eb",x"303c",x"bbeb",x"299b",x"394f",x"2a7d",x"2f38",x"3948",x"36eb",x"37e1",x"baf5",x"269a",x"394f",x"2a46",x"2f3d",x"3949",x"3714",x"35bf",x"bb76",x"27db",x"394a",x"2a4c"),
(x"3003",x"3949",x"36eb",x"b868",x"baab",x"296a",x"394f",x"2ab4",x"2f9e",x"394c",x"36eb",x"303c",x"bbeb",x"299b",x"394f",x"2a7d",x"2fa3",x"394d",x"3715",x"a836",x"bbfd",x"294f",x"394a",x"2a84"),
(x"302c",x"393d",x"3714",x"bb01",x"b7b5",x"2839",x"394a",x"2afc",x"3029",x"393d",x"36eb",x"baf3",x"b7df",x"2b38",x"394f",x"2af7",x"3003",x"3949",x"36eb",x"b868",x"baab",x"296a",x"394f",x"2ab4"),
(x"3036",x"3933",x"36eb",x"bbf9",x"ad11",x"2511",x"3950",x"2b22",x"3029",x"393d",x"36eb",x"baf3",x"b7df",x"2b38",x"394f",x"2af7",x"302c",x"393d",x"3714",x"bb01",x"b7b5",x"2839",x"394a",x"2afc"),
(x"3029",x"3929",x"36eb",x"b90c",x"3a34",x"2532",x"3950",x"2b4b",x"3036",x"3933",x"36eb",x"bbf9",x"ad11",x"2511",x"3950",x"2b22",x"3036",x"3932",x"3714",x"bbe6",x"310f",x"9bfc",x"394b",x"2b2d"),
(x"3006",x"3928",x"3714",x"2fe4",x"3bee",x"28fd",x"394b",x"2b79",x"3004",x"3929",x"36eb",x"35dd",x"3b6d",x"2be9",x"3950",x"2b72",x"3029",x"3929",x"36eb",x"b90c",x"3a34",x"2532",x"3950",x"2b4b"),
(x"2fd7",x"392c",x"3711",x"364f",x"3b52",x"2d1b",x"394c",x"2b98",x"2fdd",x"392e",x"36eb",x"32b2",x"3bc8",x"2e54",x"3950",x"2b90",x"3004",x"3929",x"36eb",x"35dd",x"3b6d",x"2be9",x"3950",x"2b72"),
(x"2f82",x"390f",x"36eb",x"bbf6",x"aa70",x"2d61",x"394f",x"2c30",x"2f71",x"3913",x"36eb",x"b9db",x"b96c",x"2c1a",x"394f",x"2c28",x"2f73",x"3913",x"3711",x"ba7a",x"b8af",x"283c",x"394b",x"2c1f"),
(x"2f85",x"392d",x"3710",x"b416",x"3bad",x"2f8b",x"394c",x"2bc3",x"2f79",x"392e",x"36eb",x"b37e",x"3bba",x"2ef6",x"3950",x"2bc4",x"2fdd",x"392e",x"36eb",x"32b2",x"3bc8",x"2e54",x"3950",x"2b90"),
(x"2efa",x"3888",x"36eb",x"35e4",x"3b4d",x"31a2",x"3977",x"2c09",x"2f46",x"387d",x"36eb",x"3b7d",x"3521",x"3096",x"3975",x"2bdb",x"2f31",x"387c",x"370f",x"3a9c",x"3854",x"30fa",x"3972",x"2c00"),
(x"2f13",x"3798",x"3715",x"bbc5",x"ab9a",x"3358",x"3993",x"306e",x"2eeb",x"3797",x"36eb",x"bb99",x"b315",x"330d",x"3998",x"306b",x"2f02",x"37ce",x"36eb",x"bb89",x"3473",x"31fc",x"3997",x"304e"),
(x"2f51",x"3919",x"3710",x"a856",x"29ab",x"3bfc",x"3951",x"38bf",x"3030",x"3914",x"3711",x"a8d9",x"252b",x"3bfe",x"393f",x"38c0",x"2fe3",x"390e",x"3718",x"ab65",x"3528",x"3b8f",x"3947",x"38c4"),
(x"300a",x"37c7",x"36eb",x"3be3",x"ace8",x"30c3",x"3991",x"30d4",x"3013",x"37ae",x"3712",x"3bcf",x"3081",x"3141",x"398f",x"30be",x"3006",x"37c2",x"3715",x"3bd7",x"31f9",x"2c2a",x"398d",x"30c6"),
(x"300a",x"37c7",x"36eb",x"3be3",x"ace8",x"30c3",x"3991",x"30d4",x"3023",x"37ad",x"36eb",x"3bdb",x"9c67",x"320a",x"3993",x"30c8",x"3013",x"37ae",x"3712",x"3bcf",x"3081",x"3141",x"398f",x"30be"),
(x"3041",x"386e",x"3710",x"3b6b",x"b5ba",x"2efe",x"3920",x"2a2b",x"3046",x"386d",x"36eb",x"3b75",x"b5a2",x"2d46",x"3925",x"2a2a",x"301f",x"385d",x"36eb",x"3958",x"b9de",x"2fe4",x"3925",x"29dd"),
(x"2f4e",x"392a",x"36eb",x"baa4",x"3859",x"2fe4",x"3950",x"2be3",x"2f79",x"392e",x"36eb",x"b37e",x"3bba",x"2ef6",x"3950",x"2bc4",x"2f85",x"392d",x"3710",x"b416",x"3bad",x"2f8b",x"394c",x"2bc3"),
(x"2fd8",x"3909",x"36eb",x"3be6",x"b08e",x"2c41",x"399b",x"2fcd",x"2fd4",x"38f6",x"36eb",x"3bfa",x"20b5",x"2cbc",x"399a",x"2fbb",x"2fc7",x"38f6",x"3715",x"3bfa",x"2710",x"2c48",x"3996",x"2fc6"),
(x"2f45",x"3921",x"3710",x"bbcc",x"3227",x"2f2f",x"394c",x"2bff",x"2f36",x"3921",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3950",x"2c05",x"2f4e",x"392a",x"36eb",x"baa4",x"3859",x"2fe4",x"3950",x"2be3"),
(x"2f46",x"387d",x"36eb",x"3b7d",x"3521",x"3096",x"3975",x"2bdb",x"2f3c",x"3877",x"36eb",x"3b19",x"b744",x"2cf7",x"3975",x"2bc7",x"2f2d",x"3876",x"370e",x"3b25",x"b70d",x"2d6a",x"3971",x"2bec"),
(x"2e90",x"38ba",x"36eb",x"b6fe",x"3b25",x"2ea4",x"39a1",x"308f",x"2f2b",x"38be",x"36eb",x"b7d8",x"3af6",x"2a35",x"39a1",x"3084",x"2f21",x"38bd",x"3711",x"b4dc",x"3b97",x"2d60",x"399e",x"3084"),
(x"2f71",x"3913",x"36eb",x"b9db",x"b96c",x"2c1a",x"394f",x"2c28",x"2f41",x"3917",x"36eb",x"bb02",x"b777",x"2fc8",x"3950",x"2c18",x"2f51",x"3919",x"3710",x"bb2f",x"b6d9",x"2e52",x"394b",x"2c11"),
(x"3015",x"385f",x"3712",x"384e",x"bab0",x"2ec8",x"3920",x"29dd",x"301f",x"385d",x"36eb",x"3958",x"b9de",x"2fe4",x"3925",x"29dd",x"2f6d",x"3851",x"36eb",x"3776",x"bb0b",x"2d41",x"3924",x"2965"),
(x"2fc7",x"38f6",x"3715",x"3bfa",x"2710",x"2c48",x"3996",x"2fc6",x"2fd4",x"38f6",x"36eb",x"3bfa",x"20b5",x"2cbc",x"399a",x"2fbb",x"2fd9",x"38f3",x"36eb",x"39df",x"3964",x"2d28",x"3999",x"2fb8"),
(x"2f2d",x"3876",x"370e",x"3b25",x"b70d",x"2d6a",x"3971",x"2bec",x"2f3c",x"3877",x"36eb",x"3b19",x"b744",x"2cf7",x"3975",x"2bc7",x"2f02",x"386c",x"36eb",x"3ad3",x"b822",x"2c4d",x"3973",x"2b9a"),
(x"2f97",x"3809",x"370e",x"bb5f",x"35f1",x"2f4f",x"3991",x"302c",x"2f8f",x"380a",x"36eb",x"bb4a",x"3677",x"2cfa",x"3995",x"3026",x"2fc6",x"381e",x"36eb",x"bbfe",x"9ea7",x"2828",x"3993",x"3011"),
(x"2f6d",x"3851",x"36eb",x"3776",x"bb0b",x"2d41",x"3924",x"2965",x"2f62",x"3850",x"36eb",x"3b24",x"371c",x"2cde",x"3924",x"295c",x"2f5c",x"3850",x"3716",x"3bde",x"b1b5",x"2825",x"391f",x"2962"),
(x"2fd6",x"38f1",x"3715",x"395d",x"39e3",x"2de3",x"3996",x"2fc1",x"2fd9",x"38f3",x"36eb",x"39df",x"3964",x"2d28",x"3999",x"2fb8",x"3026",x"38e8",x"36eb",x"39ed",x"394b",x"2f45",x"3998",x"2fa6"),
(x"2f3c",x"38c5",x"36eb",x"bbf8",x"2379",x"2d44",x"39a1",x"3080",x"2f4a",x"38c4",x"3712",x"bbf7",x"a83f",x"2d8f",x"399e",x"3080",x"2f3f",x"38c0",x"3711",x"bb12",x"3763",x"2ca3",x"399e",x"3082"),
(x"2f3f",x"38c0",x"3711",x"bb12",x"3763",x"2ca3",x"399e",x"3082",x"2f2b",x"38be",x"36eb",x"b7d8",x"3af6",x"2a35",x"39a1",x"3084",x"2f3c",x"38c5",x"36eb",x"bbf8",x"2379",x"2d44",x"39a1",x"3080"),
(x"2efb",x"386d",x"3713",x"3b5b",x"b634",x"2c08",x"3994",x"30ef",x"2f02",x"386c",x"36eb",x"3ad3",x"b822",x"2c4d",x"3997",x"30f1",x"2f01",x"386a",x"36eb",x"39e9",x"3955",x"2e31",x"3997",x"30f0"),
(x"2fc6",x"381e",x"36eb",x"bbfe",x"9ea7",x"2828",x"3993",x"3011",x"2f8f",x"3831",x"36eb",x"bab4",x"b859",x"2a59",x"3992",x"2ff8",x"2f93",x"3832",x"370f",x"bad7",x"b821",x"29e6",x"398e",x"3000"),
(x"2f62",x"3850",x"36eb",x"3b24",x"371c",x"2cde",x"3924",x"295c",x"2f83",x"384c",x"36eb",x"397a",x"39b6",x"3099",x"3924",x"2945",x"2f72",x"384b",x"3714",x"39e8",x"3951",x"2f27",x"391f",x"2948"),
(x"3026",x"38e8",x"36eb",x"39ed",x"394b",x"2f45",x"3998",x"2fa6",x"3021",x"38e4",x"36eb",x"32cb",x"bbc1",x"2fc5",x"3998",x"2fa2",x"3017",x"38e6",x"3719",x"3250",x"bbca",x"2f22",x"3995",x"2fb2"),
(x"2f3c",x"38c5",x"36eb",x"bbf8",x"2379",x"2d44",x"39a1",x"3080",x"2f33",x"38cd",x"36eb",x"bb57",x"b625",x"2e97",x"39a1",x"307b",x"2f3b",x"38cf",x"3712",x"bb92",x"b509",x"2cb4",x"399e",x"307a"),
(x"2f69",x"3862",x"36eb",x"3046",x"3be8",x"2cb7",x"3997",x"30e7",x"2f61",x"3862",x"3713",x"30a8",x"3bea",x"22dc",x"3994",x"30e5",x"2f21",x"3865",x"3710",x"3833",x"3ac7",x"2d1d",x"3994",x"30ea"),
(x"2f21",x"3865",x"3710",x"3833",x"3ac7",x"2d1d",x"3994",x"30ea",x"2f01",x"386a",x"36eb",x"39e9",x"3955",x"2e31",x"3997",x"30f0",x"2f69",x"3862",x"36eb",x"3046",x"3be8",x"2cb7",x"3997",x"30e7"),
(x"2f93",x"3832",x"370f",x"bad7",x"b821",x"29e6",x"398e",x"3000",x"2f8f",x"3831",x"36eb",x"bab4",x"b859",x"2a59",x"3992",x"2ff8",x"2f33",x"383a",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3991",x"2fdb"),
(x"2f83",x"384c",x"36eb",x"397a",x"39b6",x"3099",x"3924",x"2945",x"3000",x"383d",x"36eb",x"3aff",x"373c",x"3197",x"3925",x"28ea",x"2fe6",x"383c",x"3717",x"3a77",x"3889",x"310c",x"391f",x"28f0"),
(x"3017",x"38e6",x"3719",x"3250",x"bbca",x"2f22",x"3995",x"2fb2",x"3021",x"38e4",x"36eb",x"32cb",x"bbc1",x"2fc5",x"3998",x"2fa2",x"2fda",x"38e5",x"36eb",x"3b01",x"b745",x"3141",x"3996",x"2f98"),
(x"2f33",x"38cd",x"36eb",x"bb57",x"b625",x"2e97",x"39a1",x"307b",x"2ea7",x"38f3",x"36eb",x"bb99",x"b45f",x"30d6",x"39a2",x"3065",x"2ec5",x"38f1",x"3711",x"bb70",x"b585",x"3014",x"399f",x"3065"),
(x"2fdf",x"3866",x"36eb",x"b74a",x"3b15",x"2de4",x"3998",x"30df",x"2fe6",x"3864",x"3711",x"b934",x"3a0d",x"2c16",x"3995",x"30dc",x"2fa3",x"3862",x"3712",x"b2e8",x"3bcb",x"2c10",x"3995",x"30e1"),
(x"2fa3",x"3862",x"3712",x"b2e8",x"3bcb",x"2c10",x"3995",x"30e1",x"2f69",x"3862",x"36eb",x"3046",x"3be8",x"2cb7",x"3997",x"30e7",x"2fdf",x"3866",x"36eb",x"b74a",x"3b15",x"2de4",x"3998",x"30df"),
(x"2f33",x"383a",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3973",x"2d26",x"2f19",x"3839",x"36eb",x"38ae",x"ba73",x"2d49",x"3974",x"2d1f",x"2f20",x"383b",x"3712",x"3722",x"bb24",x"2bf2",x"3970",x"2d0b"),
(x"3000",x"383d",x"36eb",x"3aff",x"373c",x"3197",x"3925",x"28ea",x"302b",x"3821",x"36eb",x"3bbf",x"3113",x"322d",x"3924",x"286c",x"301b",x"3821",x"3713",x"3bc6",x"31be",x"30de",x"391f",x"2878"),
(x"2ea7",x"38f3",x"36eb",x"bb99",x"b45f",x"30d6",x"39a2",x"3065",x"2e7f",x"3910",x"36eb",x"bbe6",x"ac77",x"308b",x"39a2",x"3054",x"2e95",x"3910",x"3711",x"bbe4",x"ad1d",x"308b",x"399f",x"3054"),
(x"2fe6",x"3864",x"3711",x"b934",x"3a0d",x"2c16",x"3995",x"30dc",x"2fdf",x"3866",x"36eb",x"b74a",x"3b15",x"2de4",x"3998",x"30df",x"3021",x"3872",x"36eb",x"baaf",x"3860",x"2a70",x"3999",x"30d6"),
(x"2f19",x"3839",x"36eb",x"38ae",x"ba73",x"2d49",x"3974",x"2d1f",x"2efa",x"3835",x"36eb",x"2e28",x"bbe6",x"3005",x"3975",x"2d16",x"2ef3",x"3837",x"3711",x"35dd",x"bb65",x"2eae",x"3971",x"2d00"),
(x"301b",x"3821",x"3713",x"3bc6",x"31be",x"30de",x"391f",x"2878",x"302b",x"3821",x"36eb",x"3bbf",x"3113",x"322d",x"3924",x"286c",x"3025",x"3806",x"36eb",x"3bea",x"2e0a",x"2f10",x"3923",x"27f7"),
(x"2fda",x"38e5",x"36eb",x"3b01",x"b745",x"3141",x"395b",x"30e0",x"3006",x"38de",x"3715",x"39d1",x"3974",x"2cc6",x"3956",x"30d4",x"2fd8",x"38e4",x"3718",x"3af6",x"37e0",x"2460",x"3956",x"30de"),
(x"2fda",x"38e5",x"36eb",x"3b01",x"b745",x"3141",x"395b",x"30e0",x"3016",x"38dc",x"36eb",x"3a0e",x"3929",x"2e76",x"395c",x"30d2",x"3006",x"38de",x"3715",x"39d1",x"3974",x"2cc6",x"3956",x"30d4"),
(x"2e95",x"3910",x"3711",x"bbe4",x"ad1d",x"308b",x"399f",x"3054",x"2e7f",x"3910",x"36eb",x"bbe6",x"ac77",x"308b",x"39a2",x"3054",x"2e82",x"3933",x"36eb",x"bbe8",x"2d66",x"3010",x"39a3",x"3041"),
(x"3025",x"3872",x"3717",x"bb6f",x"35e4",x"261e",x"3996",x"30d2",x"3021",x"3872",x"36eb",x"baaf",x"3860",x"2a70",x"3999",x"30d6",x"302e",x"3882",x"36eb",x"bbfa",x"2c62",x"2617",x"399a",x"30ce"),
(x"2efa",x"3835",x"36eb",x"2e28",x"bbe6",x"3005",x"3975",x"2d16",x"2e9b",x"3835",x"36eb",x"b913",x"ba0d",x"310f",x"3976",x"2d00",x"2eb1",x"3838",x"3712",x"b5a6",x"bb63",x"30cc",x"3972",x"2cf1"),
(x"3025",x"3806",x"36eb",x"3bea",x"2e0a",x"2f10",x"3923",x"27f7",x"303b",x"37e1",x"36eb",x"3be4",x"2adf",x"30ee",x"3923",x"273f",x"3031",x"37df",x"370f",x"3bdd",x"30de",x"2e6c",x"391e",x"2750"),
(x"3016",x"38dc",x"36eb",x"3a0e",x"3929",x"2e76",x"395c",x"30d2",x"302e",x"38d4",x"36eb",x"3bbf",x"3333",x"2ed0",x"395c",x"30c7",x"3022",x"38d3",x"3718",x"3b13",x"3732",x"2fec",x"3956",x"30c7"),
(x"2e82",x"3933",x"36eb",x"bbe8",x"2d66",x"3010",x"39a3",x"3041",x"2ea5",x"3945",x"36eb",x"bab2",x"3834",x"30cf",x"39a3",x"3037",x"2eb5",x"3942",x"3712",x"bb45",x"3640",x"30a6",x"399f",x"3038"),
(x"2f51",x"3919",x"3710",x"bb2f",x"b6d9",x"2e52",x"394b",x"2c11",x"2f41",x"3917",x"36eb",x"bb02",x"b777",x"2fc8",x"3950",x"2c18",x"2f36",x"3921",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3950",x"2c05"),
(x"302f",x"3883",x"3715",x"bbfe",x"a412",x"2867",x"3997",x"30ca",x"302e",x"3882",x"36eb",x"bbfa",x"2c62",x"2617",x"399a",x"30ce",x"3025",x"3897",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"399b",x"30c3"),
(x"2e9b",x"3835",x"36eb",x"b913",x"ba0d",x"310f",x"3976",x"2d00",x"2e73",x"383f",x"36eb",x"bbe5",x"2dbc",x"3036",x"3977",x"2ceb",x"2e89",x"383f",x"3711",x"bbb2",x"b32f",x"30f4",x"3972",x"2cdf"),
(x"303b",x"37e1",x"36eb",x"3be4",x"2adf",x"30ee",x"3923",x"273f",x"3035",x"37ca",x"36eb",x"3af6",x"b714",x"32f0",x"3923",x"26e0",x"302a",x"37d1",x"370d",x"3b0d",x"b70c",x"3169",x"391e",x"2711"),
(x"302e",x"38d4",x"36eb",x"3bbf",x"3333",x"2ed0",x"395c",x"30c7",x"302b",x"38c8",x"36eb",x"3bbf",x"b371",x"2dad",x"395c",x"30bb",x"3027",x"38cb",x"3712",x"3bf0",x"ac20",x"2e95",x"3957",x"30be"),
(x"2ea5",x"3945",x"36eb",x"bab2",x"3834",x"30cf",x"39a3",x"3037",x"2f13",x"3955",x"36eb",x"b7cb",x"3ae6",x"3068",x"39a2",x"302c",x"2f1a",x"3951",x"3715",x"b93c",x"39e9",x"311d",x"399f",x"302d"),
(x"302a",x"3899",x"3714",x"bb81",x"b558",x"2da6",x"3998",x"30be",x"3025",x"3897",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"399b",x"30c3",x"3001",x"38a7",x"36eb",x"bac2",x"b833",x"2e85",x"399c",x"30ba"),
(x"2e73",x"383f",x"36eb",x"bbe5",x"2dbc",x"3036",x"3977",x"2ceb",x"2e9a",x"384e",x"36eb",x"b902",x"3a23",x"306a",x"3978",x"2ccb",x"2ea4",x"384b",x"3712",x"bae4",x"37c3",x"30c9",x"3973",x"2cc7"),
(x"302a",x"37d1",x"370d",x"3b0d",x"b70c",x"3169",x"391e",x"2711",x"3035",x"37ca",x"36eb",x"3af6",x"b714",x"32f0",x"3923",x"26e0",x"3020",x"37c6",x"36eb",x"3571",x"bb6d",x"30cc",x"3922",x"26b4"),
(x"302b",x"38c8",x"36eb",x"3bbf",x"b371",x"2dad",x"395c",x"30bb",x"3025",x"38c6",x"36eb",x"2eda",x"bbea",x"2e47",x"395c",x"30b8",x"301e",x"38c8",x"3712",x"3297",x"bbcc",x"2d84",x"3957",x"30ba"),
(x"2f13",x"3955",x"36eb",x"b7cb",x"3ae6",x"3068",x"39a2",x"302c",x"2f91",x"3959",x"36eb",x"95bc",x"3bf5",x"2e99",x"39a2",x"3023",x"2f91",x"3956",x"3715",x"9ef6",x"3bee",x"302a",x"399f",x"3025"),
(x"3008",x"38a8",x"3715",x"ba65",x"b8c1",x"2d9e",x"3999",x"30b5",x"3001",x"38a7",x"36eb",x"bac2",x"b833",x"2e85",x"399c",x"30ba",x"2fc1",x"38b1",x"36eb",x"b9cd",x"b979",x"2caa",x"399d",x"30b3"),
(x"2e9a",x"384e",x"36eb",x"b902",x"3a23",x"306a",x"3978",x"2ccb",x"2ef3",x"3850",x"36eb",x"b3f1",x"3bbc",x"2b58",x"3978",x"2cb3",x"2eea",x"384e",x"3713",x"b607",x"3b5e",x"2e4d",x"3973",x"2cb3"),
(x"301d",x"37cb",x"3713",x"3451",x"bbac",x"2d81",x"391d",x"26f7",x"3020",x"37c6",x"36eb",x"3571",x"bb6d",x"30cc",x"3922",x"26b4",x"300a",x"37c7",x"36eb",x"3be3",x"ace8",x"30c3",x"3922",x"268a"),
(x"301e",x"38c8",x"3712",x"3297",x"bbcc",x"2d84",x"3957",x"30ba",x"3025",x"38c6",x"36eb",x"2eda",x"bbea",x"2e47",x"395c",x"30b8",x"2ffe",x"38c7",x"36eb",x"2c58",x"bbf7",x"2bc5",x"395b",x"30ae"),
(x"2f91",x"3956",x"3715",x"9ef6",x"3bee",x"302a",x"399f",x"3025",x"2f91",x"3959",x"36eb",x"95bc",x"3bf5",x"2e99",x"39a2",x"3023",x"3007",x"3955",x"36eb",x"366a",x"3b44",x"2f81",x"39a2",x"301a"),
(x"2fc7",x"38b2",x"3717",x"b939",x"ba0b",x"29e0",x"399a",x"30ae",x"2fc1",x"38b1",x"36eb",x"b9cd",x"b979",x"2caa",x"399d",x"30b3",x"2fa3",x"38b4",x"36eb",x"35a6",x"bb74",x"2d53",x"399d",x"30b1"),
(x"2eea",x"384e",x"3713",x"b607",x"3b5e",x"2e4d",x"3973",x"2cb3",x"2ef3",x"3850",x"36eb",x"b3f1",x"3bbc",x"2b58",x"3978",x"2cb3",x"2f03",x"3852",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3978",x"2cad"),
(x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d",x"2f27",x"37cb",x"3715",x"19bc",x"26cf",x"3bff",x"394e",x"396e",x"2f97",x"3809",x"370e",x"b004",x"271d",x"3bef",x"3949",x"3959"),
(x"3006",x"37c2",x"3715",x"a58e",x"b07a",x"3beb",x"393f",x"396f",x"3013",x"37ae",x"3712",x"29f0",x"ab1d",x"3bfa",x"393c",x"3975",x"2f27",x"37cb",x"3715",x"19bc",x"26cf",x"3bff",x"394e",x"396e"),
(x"2f27",x"37cb",x"3715",x"19bc",x"26cf",x"3bff",x"394e",x"396e",x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d",x"3006",x"37c2",x"3715",x"a58e",x"b07a",x"3beb",x"393f",x"396f"),
(x"2f97",x"3809",x"370e",x"b004",x"271d",x"3bef",x"3949",x"3959",x"3020",x"3806",x"3717",x"abf6",x"a5ae",x"3bfb",x"393d",x"395a",x"3008",x"37c9",x"3716",x"a0ea",x"2786",x"3bfe",x"393f",x"396d"),
(x"2ffe",x"38c7",x"36eb",x"2c58",x"bbf7",x"2bc5",x"395b",x"30ae",x"2fea",x"38c5",x"36eb",x"3a76",x"b8ad",x"2cce",x"395b",x"30ab",x"2fe7",x"38c7",x"3716",x"38f4",x"ba42",x"2c09",x"3956",x"30af"),
(x"300a",x"3951",x"3713",x"382e",x"3aba",x"306c",x"399e",x"301c",x"3007",x"3955",x"36eb",x"366a",x"3b44",x"2f81",x"39a2",x"301a",x"3051",x"3947",x"36eb",x"39f2",x"3938",x"30b5",x"39a1",x"300e"),
(x"2f4c",x"38a8",x"36eb",x"3976",x"b9cc",x"2dcc",x"399e",x"30a9",x"2f4f",x"38ab",x"3714",x"397e",x"b9c5",x"2dbf",x"399b",x"30a5",x"2f79",x"38b1",x"3714",x"39a7",x"b99f",x"2d1e",x"399b",x"30a9"),
(x"2f79",x"38b1",x"3714",x"39a7",x"b99f",x"2d1e",x"399b",x"30a9",x"2fa3",x"38b4",x"36eb",x"35a6",x"bb74",x"2d53",x"399d",x"30b1",x"2f4c",x"38a8",x"36eb",x"3976",x"b9cc",x"2dcc",x"399e",x"30a9"),
(x"2f03",x"3852",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3978",x"2cad",x"2ea2",x"3855",x"36eb",x"b9ec",x"b92b",x"31e4",x"3979",x"2c94",x"2ec3",x"3856",x"3711",x"b8c8",x"ba4e",x"30a8",x"3974",x"2c94"),
(x"3046",x"3945",x"3715",x"3ae0",x"37cf",x"30d4",x"399d",x"3011",x"3051",x"3947",x"36eb",x"39f2",x"3938",x"30b5",x"39a1",x"300e",x"306a",x"3934",x"36eb",x"3bc4",x"327a",x"3012",x"39a0",x"3004"),
(x"2f4c",x"38a8",x"36eb",x"3976",x"b9cc",x"2dcc",x"399e",x"30a9",x"2f11",x"38a3",x"36eb",x"353f",x"bb87",x"2d28",x"399f",x"30a4",x"2f0c",x"38a4",x"3716",x"37d6",x"baf0",x"2d8e",x"399c",x"309f"),
(x"2ea2",x"3855",x"36eb",x"b9ec",x"b92b",x"31e4",x"3979",x"2c94",x"2e56",x"3866",x"36eb",x"bbbc",x"b212",x"3175",x"3979",x"2c6b",x"2e71",x"3866",x"370f",x"bb4b",x"b5cc",x"3223",x"3974",x"2c6c"),
(x"3023",x"37ad",x"36eb",x"3bdb",x"9c67",x"320a",x"3993",x"30c8",x"3014",x"377e",x"36eb",x"3ade",x"b7ab",x"31d3",x"3996",x"30b2",x"3008",x"3783",x"370e",x"3b7b",x"b4a9",x"3270",x"3992",x"30ab"),
(x"2fda",x"38c4",x"3715",x"3a5f",x"3873",x"3388",x"391d",x"2bab",x"3025",x"38b5",x"36eb",x"3afe",x"375c",x"30f4",x"3923",x"2b64",x"300d",x"38b7",x"3718",x"3ac6",x"37dc",x"3286",x"391d",x"2b6d"),
(x"3061",x"3933",x"3715",x"3bec",x"2be2",x"2fce",x"399c",x"3007",x"306a",x"3934",x"36eb",x"3bc4",x"327a",x"3012",x"39a0",x"3004",x"3065",x"3921",x"36eb",x"3b6e",x"b575",x"309e",x"399e",x"2ff4"),
(x"2f2f",x"38f9",x"3714",x"b05e",x"a194",x"3bec",x"3953",x"38d0",x"2e95",x"3910",x"3711",x"acd1",x"a504",x"3bf9",x"395d",x"38c4",x"2ed8",x"3913",x"3713",x"b0f4",x"99bc",x"3be7",x"3959",x"38c2"),
(x"2f2f",x"38f9",x"3714",x"b05e",x"a194",x"3bec",x"3953",x"38d0",x"2ec5",x"38f1",x"3711",x"b115",x"a7d5",x"3be4",x"395a",x"38d5",x"2e95",x"3910",x"3711",x"acd1",x"a504",x"3bf9",x"395d",x"38c4"),
(x"2f11",x"38a3",x"36eb",x"353f",x"bb87",x"2d28",x"399f",x"30a4",x"2ec4",x"38a1",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"39a0",x"309f",x"2ecb",x"38a3",x"3716",x"a345",x"bbf7",x"2dcc",x"399c",x"309b"),
(x"2e56",x"3866",x"36eb",x"bbbc",x"b212",x"3175",x"3979",x"2c6b",x"2e52",x"387a",x"36eb",x"bb61",x"35a0",x"3119",x"3978",x"2c41",x"2e69",x"3879",x"370f",x"bbd3",x"2f46",x"3182",x"3974",x"2c45"),
(x"3025",x"38b5",x"36eb",x"3afe",x"375c",x"30f4",x"3923",x"2b64",x"304c",x"389f",x"36eb",x"3bba",x"3376",x"2f14",x"3924",x"2afe",x"3041",x"389f",x"3714",x"3b6b",x"3587",x"3095",x"391f",x"2afc"),
(x"3065",x"3921",x"36eb",x"3b6e",x"b575",x"309e",x"399e",x"2ff4",x"303a",x"3911",x"36eb",x"3884",x"ba69",x"3249",x"399d",x"2fe2",x"3030",x"3914",x"3711",x"38a4",x"ba69",x"309a",x"399a",x"2fec"),
(x"2ec4",x"38a1",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"39a0",x"309f",x"2e81",x"38a5",x"36eb",x"bacb",x"b812",x"3064",x"39a0",x"309b",x"2e97",x"38a6",x"3714",x"b976",x"b9c0",x"3024",x"399d",x"3098"),
(x"2e52",x"387a",x"36eb",x"bb61",x"35a0",x"3119",x"3978",x"2c41",x"2e9d",x"3886",x"36eb",x"b86e",x"3a87",x"313e",x"3978",x"2c22",x"2ea1",x"3883",x"370f",x"b891",x"3a72",x"30f5",x"3974",x"2c2c"),
(x"3014",x"377e",x"36eb",x"3ade",x"b7ab",x"31d3",x"3996",x"30b2",x"2fa3",x"3756",x"36eb",x"38a6",x"ba54",x"3207",x"3998",x"3099",x"2fa8",x"3761",x"3712",x"38b5",x"ba3e",x"32bc",x"3994",x"3095"),
(x"304c",x"389f",x"36eb",x"3bba",x"3376",x"2f14",x"3924",x"2afe",x"305b",x"3885",x"36eb",x"3bef",x"ad09",x"2e69",x"3924",x"2a8f",x"3052",x"3886",x"3712",x"3bf0",x"2a00",x"2f46",x"3920",x"2a91"),
(x"3030",x"3914",x"3711",x"38a4",x"ba69",x"309a",x"399a",x"2fec",x"303a",x"3911",x"36eb",x"3884",x"ba69",x"3249",x"399d",x"2fe2",x"2fed",x"390e",x"36eb",x"360d",x"bb5a",x"2ef3",x"399b",x"2fd2"),
(x"2e81",x"38a5",x"36eb",x"bacb",x"b812",x"3064",x"39a0",x"309b",x"2e6a",x"38b0",x"36eb",x"bbcf",x"3174",x"3043",x"39a1",x"3095",x"2e81",x"38af",x"3712",x"bbe0",x"ae5e",x"30a3",x"399d",x"3093"),
(x"2ea1",x"3883",x"370f",x"b891",x"3a72",x"30f5",x"3974",x"2c2c",x"2e9d",x"3886",x"36eb",x"b86e",x"3a87",x"313e",x"3978",x"2c22",x"2efa",x"3888",x"36eb",x"35e4",x"3b4d",x"31a2",x"3977",x"2c09"),
(x"2fa8",x"3761",x"3712",x"38b5",x"ba3e",x"32bc",x"3994",x"3095",x"2fa3",x"3756",x"36eb",x"38a6",x"ba54",x"3207",x"3998",x"3099",x"2f52",x"3756",x"36eb",x"b996",x"b95e",x"33ec",x"3999",x"308f"),
(x"305b",x"3885",x"36eb",x"3bef",x"ad09",x"2e69",x"3924",x"2a8f",x"3046",x"386d",x"36eb",x"3b75",x"b5a2",x"2d46",x"3925",x"2a2a",x"3041",x"386e",x"3710",x"3b6b",x"b5ba",x"2efe",x"3920",x"2a2b"),
(x"2fe3",x"390e",x"3718",x"38ae",x"ba78",x"2b7c",x"3998",x"2fdf",x"2fed",x"390e",x"36eb",x"360d",x"bb5a",x"2ef3",x"399b",x"2fd2",x"2fd8",x"3909",x"36eb",x"3be6",x"b08e",x"2c41",x"399b",x"2fcd"),
(x"2e6a",x"38b0",x"36eb",x"bbcf",x"3174",x"3043",x"39a1",x"3095",x"2e90",x"38ba",x"36eb",x"b6fe",x"3b25",x"2ea4",x"39a1",x"308f",x"2e99",x"38b7",x"3714",x"b972",x"39bb",x"30de",x"399d",x"308e"),
(x"2ec4",x"3925",x"3710",x"2828",x"a60a",x"3bfe",x"395a",x"38b8",x"2ed8",x"3913",x"3713",x"b0f4",x"99bc",x"3be7",x"3959",x"38c2",x"2e95",x"3910",x"3711",x"acd1",x"a504",x"3bf9",x"395d",x"38c4"),
(x"2e95",x"3932",x"3714",x"2eb0",x"a8fa",x"3bf3",x"395e",x"38b1",x"2eca",x"3935",x"3714",x"2946",x"9ffc",x"3bfe",x"395a",x"38af",x"2ec4",x"3925",x"3710",x"2828",x"a60a",x"3bfe",x"395a",x"38b8"),
(x"2eb5",x"3942",x"3712",x"a587",x"a08e",x"3bff",x"395c",x"38a8",x"2eca",x"3935",x"3714",x"2946",x"9ffc",x"3bfe",x"395a",x"38af",x"2e95",x"3932",x"3714",x"2eb0",x"a8fa",x"3bf3",x"395e",x"38b1"),
(x"2eb5",x"3942",x"3712",x"a587",x"a08e",x"3bff",x"395c",x"38a8",x"2edf",x"393d",x"3712",x"2953",x"a7ae",x"3bfd",x"3959",x"38aa",x"2eca",x"3935",x"3714",x"2946",x"9ffc",x"3bfe",x"395a",x"38af"),
(x"2f1a",x"3951",x"3715",x"a0ea",x"aafd",x"3bfc",x"3956",x"389f",x"2f3d",x"3949",x"3714",x"231d",x"ab5f",x"3bfc",x"3953",x"38a3",x"2f06",x"3944",x"3714",x"a8bf",x"ac22",x"3bfa",x"3957",x"38a7"),
(x"2f91",x"3956",x"3715",x"27e2",x"a9b5",x"3bfc",x"394e",x"389b",x"2fa3",x"394d",x"3715",x"270a",x"2779",x"3bfe",x"394d",x"38a1",x"2f3d",x"3949",x"3714",x"231d",x"ab5f",x"3bfc",x"3953",x"38a3"),
(x"300a",x"3951",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3946",x"389e",x"3004",x"394a",x"3716",x"24bc",x"2ceb",x"3bf9",x"3946",x"38a2",x"2fa3",x"394d",x"3715",x"270a",x"2779",x"3bfe",x"394d",x"38a1"),
(x"3046",x"3945",x"3715",x"a266",x"1d87",x"3bff",x"393e",x"38a4",x"302c",x"393d",x"3714",x"a8e0",x"a99e",x"3bfc",x"3941",x"38a9",x"3004",x"394a",x"3716",x"24bc",x"2ceb",x"3bf9",x"3946",x"38a2"),
(x"3061",x"3933",x"3715",x"a891",x"27ce",x"3bfd",x"3939",x"38ae",x"3036",x"3932",x"3714",x"a538",x"29ab",x"3bfd",x"393f",x"38af",x"302c",x"393d",x"3714",x"a8e0",x"a99e",x"3bfc",x"3941",x"38a9"),
(x"3061",x"3933",x"3715",x"a891",x"27ce",x"3bfd",x"3939",x"38ae",x"3058",x"3922",x"3717",x"ad04",x"a793",x"3bf8",x"393a",x"38b8",x"3026",x"3929",x"3715",x"ac67",x"a8a5",x"3bf9",x"3941",x"38b4"),
(x"3030",x"3914",x"3711",x"a8d9",x"252b",x"3bfe",x"393f",x"38c0",x"3006",x"3928",x"3714",x"aa45",x"ab10",x"3bfa",x"3945",x"38b5",x"3026",x"3929",x"3715",x"ac67",x"a8a5",x"3bf9",x"3941",x"38b4"),
(x"2f5e",x"3928",x"3711",x"abef",x"28a8",x"3bfa",x"3950",x"38b6",x"2f85",x"392d",x"3710",x"a352",x"2e7e",x"3bf5",x"394e",x"38b3",x"2fd7",x"392c",x"3711",x"aa66",x"3318",x"3bca",x"3949",x"38b3"),
(x"2f89",x"3910",x"3713",x"b41f",x"2c3a",x"3bb6",x"394d",x"38c4",x"2f73",x"3913",x"3711",x"b40c",x"a6bb",x"3bbc",x"394f",x"38c1",x"2fe3",x"390e",x"3718",x"ab65",x"3528",x"3b8f",x"3947",x"38c4"),
(x"2f8e",x"3906",x"3714",x"ade0",x"24c2",x"3bf6",x"394d",x"38c9",x"2fcc",x"3909",x"3718",x"b420",x"9418",x"3bba",x"3948",x"38c7",x"2fc7",x"38f6",x"3715",x"a7ae",x"24ea",x"3bfe",x"3949",x"38d2"),
(x"2f8e",x"3906",x"3714",x"ade0",x"24c2",x"3bf6",x"394d",x"38c9",x"2f89",x"3910",x"3713",x"b41f",x"2c3a",x"3bb6",x"394d",x"38c4",x"2fcc",x"3909",x"3718",x"b420",x"9418",x"3bba",x"3948",x"38c7"),
(x"2f5e",x"3928",x"3711",x"abef",x"28a8",x"3bfa",x"3950",x"38b6",x"2f51",x"3919",x"3710",x"a856",x"29ab",x"3bfc",x"3951",x"38bf",x"2f45",x"3921",x"3710",x"aa8d",x"a973",x"3bfb",x"3952",x"38ba"),
(x"3006",x"3928",x"3714",x"aa45",x"ab10",x"3bfa",x"3945",x"38b5",x"3030",x"3914",x"3711",x"a8d9",x"252b",x"3bfe",x"393f",x"38c0",x"2f51",x"3919",x"3710",x"a856",x"29ab",x"3bfc",x"3951",x"38bf"),
(x"2f82",x"390f",x"36eb",x"bbf6",x"aa70",x"2d61",x"394f",x"2c30",x"2f89",x"3910",x"3713",x"bbc2",x"b3a4",x"298a",x"394a",x"2c28",x"2f8e",x"3906",x"3714",x"bbf3",x"2e23",x"2b27",x"394a",x"2c3b"),
(x"2f8e",x"3906",x"3714",x"bbf3",x"2e23",x"2b27",x"394a",x"2c3b",x"2f6c",x"38ee",x"36eb",x"b46a",x"3b91",x"316a",x"394e",x"2c76",x"2f82",x"390f",x"36eb",x"bbf6",x"aa70",x"2d61",x"394f",x"2c30"),
(x"3a25",x"3c7f",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0",x"3a26",x"3c69",x"3710",x"3bcf",x"2680",x"32dc",x"39f4",x"33ca",x"3a20",x"3c69",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa"),
(x"3a1f",x"3c7f",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a20",x"3c69",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa",x"3a19",x"3c69",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392"),
(x"3a18",x"3c7f",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a19",x"3c69",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392",x"3a14",x"3c69",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387"),
(x"3a10",x"3c7f",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a14",x"3c69",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387",x"3a0d",x"3c69",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b"),
(x"3a09",x"3c7f",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"39fc",x"3c80",x"3713",x"af5f",x"3bdb",x"30c1",x"3bc0",x"39a6",x"3a03",x"3c81",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bbd",x"39a7"),
(x"3a09",x"3c81",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a11",x"3c81",x"374a",x"b547",x"b37e",x"3b50",x"3bb7",x"399b",x"3a10",x"3c7f",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b"),
(x"39fc",x"3c69",x"3710",x"ba72",x"9a8d",x"38bc",x"39f2",x"333e",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e",x"3a02",x"3c68",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352"),
(x"3a02",x"3c96",x"3711",x"bbe1",x"a6cf",x"3179",x"3be9",x"39fb",x"3a04",x"3c96",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7",x"3a03",x"3c81",x"370e",x"bbc2",x"ab4f",x"338c",x"3bf9",x"39fa"),
(x"3a08",x"3c96",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a0f",x"3c96",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a11",x"3c81",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed"),
(x"3a0f",x"3c96",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a17",x"3c96",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3be8",x"39eb",x"3a19",x"3c82",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a1d",x"3c96",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a21",x"3c81",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6",x"3a19",x"3c82",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a24",x"3c96",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a25",x"3c81",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3",x"3a21",x"3c81",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6"),
(x"3a2a",x"3c96",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a2d",x"3c81",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a25",x"3c81",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3"),
(x"3a2d",x"3c81",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a2a",x"3c96",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a2f",x"3c96",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"3a25",x"3c81",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a2d",x"3c81",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a",x"3a25",x"3c7f",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c"),
(x"3a0d",x"3c69",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b",x"3a07",x"3c69",x"373c",x"bac4",x"2853",x"3841",x"39f2",x"336a",x"3a09",x"3c7f",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369"),
(x"3a11",x"3c81",x"374a",x"b547",x"b37e",x"3b50",x"3bb7",x"399b",x"3a19",x"3c82",x"374d",x"3243",x"b807",x"3abb",x"3bb5",x"3999",x"3a18",x"3c7f",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998"),
(x"3a18",x"3c7f",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998",x"3a19",x"3c82",x"374d",x"3243",x"b807",x"3abb",x"3bb5",x"3999",x"3a21",x"3c81",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a25",x"3c81",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a1f",x"3c7f",x"3733",x"3800",x"ba99",x"3436",x"3bb7",x"3993",x"3a21",x"3c81",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a2a",x"3c96",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a20",x"3c97",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b",x"3a26",x"3c97",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3a24",x"3c96",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a1a",x"3c97",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e",x"3a20",x"3c97",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b"),
(x"3a1d",x"3c96",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e",x"3a15",x"3c97",x"374b",x"aaab",x"39a7",x"39a5",x"3b22",x"3871",x"3a1a",x"3c97",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e"),
(x"3a17",x"3c96",x"3751",x"2fda",x"39a6",x"3994",x"3b24",x"3871",x"3a15",x"3c97",x"374b",x"aaab",x"39a7",x"39a5",x"3b22",x"3871",x"3a1d",x"3c96",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e"),
(x"3a0f",x"3c96",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a0f",x"3c97",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873",x"3a15",x"3c97",x"374b",x"aaab",x"39a7",x"39a5",x"3b22",x"3871"),
(x"3a08",x"3c96",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a09",x"3c98",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875",x"3a0f",x"3c97",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873"),
(x"3a04",x"3c96",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879",x"3a01",x"3c97",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879",x"3a09",x"3c98",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875"),
(x"3a02",x"3c96",x"3711",x"b40d",x"bb3a",x"3585",x"3b18",x"387b",x"3a01",x"3c97",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879",x"3a04",x"3c96",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879"),
(x"3a02",x"3c96",x"3711",x"b40d",x"bb3a",x"3585",x"3b18",x"387b",x"39fb",x"3c97",x"3713",x"aedc",x"bb7b",x"3565",x"3b16",x"387a",x"3a01",x"3c97",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879"),
(x"3a02",x"3c96",x"3711",x"315a",x"2baa",x"3bdf",x"3a19",x"3349",x"3a03",x"3c81",x"370e",x"34eb",x"a6e9",x"3b9c",x"3a06",x"334b",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3a24",x"3cae",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a27",x"3cae",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9",x"3a26",x"3c97",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4"),
(x"3a24",x"3cae",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a20",x"3c97",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a21",x"3cae",x"373a",x"3acd",x"a5ae",x"3834",x"3a2d",x"33a3"),
(x"3a20",x"3c97",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a1a",x"3c97",x"3746",x"38a5",x"a839",x"3a81",x"3a1a",x"338e",x"3a1a",x"3cae",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a15",x"3c97",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a14",x"3cae",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385",x"3a1a",x"3cae",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a0f",x"3c97",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a0d",x"3cad",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378",x"3a14",x"3cae",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385"),
(x"3a09",x"3c98",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a07",x"3cae",x"373c",x"baa1",x"a6bb",x"3879",x"3a2d",x"3366",x"3a0d",x"3cad",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378"),
(x"3a09",x"3c98",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a01",x"3c97",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"3a00",x"3cad",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c"),
(x"3a01",x"3c97",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"39fb",x"3c97",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"39fc",x"3cae",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340"),
(x"3475",x"3c8f",x"3710",x"0000",x"0000",x"3c00",x"3a13",x"2451",x"3485",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"3485",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"3485",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"349b",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"349b",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f"),
(x"349b",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"34bb",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2643",x"34bb",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643"),
(x"34bb",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643",x"34bb",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2643",x"34cb",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"34cb",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3",x"34e9",x"3c9d",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"278b",x"34e9",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b"),
(x"34e9",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b",x"34e9",x"3c9d",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"278b",x"3501",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"3501",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a",x"351b",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"351b",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878"),
(x"351b",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"353f",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"353f",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"353f",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"3555",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"3555",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949"),
(x"3555",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"357d",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"357d",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"357d",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"3592",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20",x"3592",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"363b",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"363b",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2c3f",x"36f7",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"363b",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"362c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"362c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"362c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"3592",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20",x"3592",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"35f5",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b84",x"35fd",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2ba0",x"35fd",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"35e4",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35fd",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0",x"35f3",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"35d3",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35f3",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d",x"35f1",x"3ca0",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"35f5",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b84",x"35e4",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35fd",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"35e4",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35d3",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35f3",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"35d3",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35bd",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"35f1",x"3c76",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"35bd",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"359e",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"35bd",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35f1",x"3ca0",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"3587",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"29f9",x"358a",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"2a04",x"3593",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"36f7",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d",x"3710",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2dbb",x"3710",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"380a",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b",x"37b8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2ee7",x"37b8",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"37b8",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7",x"37b8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2ee7",x"37a8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"37a8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9",x"378c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"378c",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"378c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"376c",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2e5e",x"376c",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"376c",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e",x"376c",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2e5e",x"3752",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"36f7",x"3cb2",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e",x"3716",x"3cb1",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"36df",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"3716",x"3cb1",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"372e",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0",x"36dc",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"36df",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"3716",x"3c65",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4",x"36f7",x"3c65",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"36dc",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"372e",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3716",x"3c65",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"3753",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2e32",x"3742",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"375f",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"3742",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"372e",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3754",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"3753",x"3cad",x"3710",x"0000",x"0000",x"3c00",x"3a2c",x"2e32",x"3760",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2e49",x"375f",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"3742",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"375f",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47",x"3754",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"36cb",x"3c9d",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2d40",x"36c2",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2d2f",x"36c4",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"36cb",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"2d40",x"3705",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"36c4",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"3705",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"3713",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"36dc",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"3705",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36c4",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33",x"36dc",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"3713",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"36dc",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e",x"372e",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"372e",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"36dc",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"3713",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"3713",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3754",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33",x"3752",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"3713",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"3716",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5",x"3752",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"3710",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb",x"3710",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2dbb",x"3716",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"3752",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"3752",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30",x"3716",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"3813",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"3813",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac",x"380a",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"382a",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"382a",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2ffc",x"3813",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"382a",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3885",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30a2",x"3885",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"388c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"388c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"3885",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"38bf",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38bf",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"3109",x"38d5",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130"),
(x"38bf",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38b2",x"3c7d",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b2",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"38b2",x"3c7d",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b0",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"38b0",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38b0",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"388c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"388c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"3872",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"3877",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088",x"386d",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3076"),
(x"3885",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"3894",x"3c67",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc",x"3877",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088"),
(x"386d",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"3076",x"3877",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3872",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080"),
(x"3877",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3894",x"3caf",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"3885",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"3894",x"3caf",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"38b7",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"388c",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"388c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"38b7",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"3894",x"3c67",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"38d8",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3135",x"38c7",x"3c6c",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38d4",x"3c73",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d"),
(x"38d8",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3135",x"38d9",x"3ca6",x"3710",x"0000",x"0000",x"3c00",x"3a26",x"3136",x"38d4",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d"),
(x"38c7",x"3cab",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38d4",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d",x"38c9",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a"),
(x"38c7",x"3c6c",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38b7",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38c9",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a"),
(x"388c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"388c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"38b0",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"388c",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae",x"38b2",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"38b0",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38b2",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"38b7",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"388c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae"),
(x"38b7",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38b2",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"388c",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"38f6",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"38f6",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b",x"38d5",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130"),
(x"3915",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"3915",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"31a2",x"38f6",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b"),
(x"3915",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"392f",x"3cab",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"31d0",x"392f",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"393f",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"393f",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed",x"392f",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"3953",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"3953",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211",x"393f",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"395a",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"395a",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d",x"3953",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211"),
(x"395d",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"395d",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"3222",x"395a",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d"),
(x"395d",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"3963",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"322d",x"3963",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3972",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3972",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248",x"3963",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3985",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3985",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"3269",x"3972",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248"),
(x"3985",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3994",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3284",x"3994",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3999",x"3cac",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"3999",x"3c6a",x"3710",x"96f6",x"9f93",x"3c00",x"39f3",x"328d",x"3994",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3999",x"3cac",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39fb",x"3c97",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e"),
(x"39f5",x"3cae",x"3710",x"b60a",x"25b5",x"3b67",x"3a2d",x"3331",x"39fc",x"3cae",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340",x"39fb",x"3c97",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d"),
(x"3999",x"3c6a",x"3710",x"96f6",x"9f93",x"3c00",x"39f3",x"328d",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e",x"39fc",x"3c69",x"3710",x"ba72",x"9a8d",x"38bc",x"39f2",x"333e"),
(x"3a0d",x"3cad",x"374b",x"a412",x"3bfd",x"2963",x"3bce",x"3a59",x"3a07",x"3cae",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a1a",x"3cae",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e"),
(x"3a07",x"3cae",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a00",x"3cad",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"3a21",x"3cae",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60"),
(x"3a00",x"3cad",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"39fc",x"3cae",x"3718",x"135f",x"3bfd",x"299e",x"3bd8",x"3a52",x"3a24",x"3cae",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62"),
(x"39fc",x"3cae",x"3718",x"135f",x"3bfd",x"299e",x"3bd8",x"3a52",x"39f5",x"3cae",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f",x"3a27",x"3cae",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63"),
(x"3a19",x"3c69",x"3749",x"209b",x"bc00",x"135f",x"3a90",x"3a5e",x"3a07",x"3c69",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a8e",x"3a57",x"3a0d",x"3c69",x"374b",x"1481",x"bbff",x"269a",x"3a91",x"3a59"),
(x"3a20",x"3c69",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a02",x"3c68",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55",x"3a07",x"3c69",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a8e",x"3a57"),
(x"3a26",x"3c69",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63",x"39fc",x"3c69",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53",x"3a02",x"3c68",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55"),
(x"34e9",x"3c7a",x"36da",x"b699",x"bb49",x"0000",x"3a6e",x"3b90",x"34e9",x"3c7a",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90",x"3501",x"3c78",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94"),
(x"3872",x"3c78",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"3872",x"3c78",x"3710",x"b9d1",x"397d",x"0000",x"3a95",x"3a08",x"386c",x"3c74",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c"),
(x"3813",x"3c97",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"3813",x"3c97",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5",x"380a",x"3c97",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9"),
(x"34cb",x"3c7e",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34cb",x"3c7e",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89",x"34e9",x"3c7a",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90"),
(x"39fc",x"3c69",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"39fc",x"3c69",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53",x"3a26",x"3c69",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63"),
(x"3885",x"3c7c",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"3885",x"3c7c",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00",x"3872",x"3c78",x"3710",x"b9d1",x"397d",x"0000",x"3a95",x"3a08"),
(x"375f",x"3ca7",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"375f",x"3ca7",x"3710",x"3bc1",x"b3d7",x"068d",x"3aa1",x"3a26",x"3760",x"3ca9",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28"),
(x"34bb",x"3c7f",x"36da",x"b13f",x"bbe4",x"0000",x"3a6e",x"3b86",x"34bb",x"3c7f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86",x"34cb",x"3c7e",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89"),
(x"388c",x"3c7e",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"388c",x"3c7e",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd",x"3885",x"3c7c",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00"),
(x"380a",x"3c97",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"380a",x"3c97",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9",x"37b8",x"3c94",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b"),
(x"349b",x"3c80",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"349b",x"3c80",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80",x"34bb",x"3c7f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86"),
(x"388c",x"3c80",x"36da",x"b967",x"b9e6",x"0000",x"3a8a",x"39fb",x"388c",x"3c80",x"3710",x"bb52",x"b671",x"0000",x"3a95",x"39fb",x"388c",x"3c7e",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd"),
(x"37b8",x"3c94",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"37b8",x"3c94",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b",x"37a8",x"3c95",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e"),
(x"3485",x"3c82",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"3485",x"3c82",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b",x"349b",x"3c80",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80"),
(x"3885",x"3c81",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"3885",x"3c81",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf",x"388c",x"3c80",x"3710",x"bb52",x"b671",x"0000",x"3a87",x"3bb2"),
(x"37a8",x"3c95",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"37a8",x"3c95",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e",x"378c",x"3c99",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14"),
(x"3a2f",x"3c96",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"385a",x"3a2f",x"3c96",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"3861",x"3a26",x"3c97",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3475",x"3c87",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3475",x"3c87",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77",x"3485",x"3c82",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b"),
(x"3753",x"3c6a",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3753",x"3c6a",x"3710",x"38fe",x"ba3f",x"8000",x"3a87",x"3b4e",x"3760",x"3c6d",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52"),
(x"378c",x"3c99",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"378c",x"3c99",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14",x"376c",x"3c9c",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a"),
(x"382a",x"3c81",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"382a",x"3c81",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d",x"3885",x"3c81",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf"),
(x"376c",x"3c9c",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"376c",x"3c9c",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a",x"3752",x"3ca1",x"3710",x"3bfd",x"aac2",x"0000",x"3aa1",x"3a21"),
(x"3999",x"3c6a",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"3999",x"3c6a",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d",x"39fc",x"3c69",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53"),
(x"3813",x"3c7f",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"3813",x"3c7f",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84",x"382a",x"3c81",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d"),
(x"3753",x"3cad",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3753",x"3cad",x"3710",x"37e4",x"3af5",x"868d",x"3aa1",x"3a2b",x"3742",x"3cae",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f"),
(x"380a",x"3c7f",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"380a",x"3c7f",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81",x"3813",x"3c7f",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84"),
(x"3742",x"3cae",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"3742",x"3cae",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f",x"372e",x"3cae",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32"),
(x"3760",x"3c6d",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"3760",x"3c6d",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52",x"375f",x"3c70",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54"),
(x"372e",x"3cae",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"372e",x"3cae",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32",x"3716",x"3cb1",x"3710",x"32c2",x"3bd1",x"0000",x"3aa1",x"3a37"),
(x"37b8",x"3c82",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"37b8",x"3c82",x"3710",x"2df5",x"bbf7",x"0000",x"3a87",x"3b6f",x"380a",x"3c7f",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81"),
(x"3716",x"3cb1",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"3716",x"3cb1",x"3710",x"32c2",x"3bd1",x"0000",x"3aa1",x"3a37",x"36f7",x"3cb2",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d"),
(x"37a8",x"3c82",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"37a8",x"3c82",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c",x"37b8",x"3c82",x"3710",x"2df5",x"bbf7",x"0000",x"3a87",x"3b6f"),
(x"36f7",x"3cb2",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"36f7",x"3cb2",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d",x"36e3",x"3caf",x"3710",x"bb17",x"3766",x"068d",x"3aa1",x"3a41"),
(x"378c",x"3c7e",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"378c",x"3c7e",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66",x"37a8",x"3c82",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c"),
(x"36e3",x"3caf",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36e3",x"3caf",x"3710",x"bb17",x"3766",x"068d",x"3aa1",x"3a41",x"36df",x"3cac",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44"),
(x"376c",x"3c7b",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"376c",x"3c7b",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f",x"378c",x"3c7e",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66"),
(x"36df",x"3cac",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36df",x"3cac",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44",x"36dc",x"3ca9",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47"),
(x"3a26",x"3c97",x"36da",x"3bff",x"a4d0",x"0000",x"3a18",x"33f3",x"3a26",x"3c97",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4",x"3a27",x"3cae",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9"),
(x"39f5",x"3cae",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"39f5",x"3cae",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f",x"3999",x"3cac",x"3710",x"b329",x"3bcb",x"868d",x"3bd9",x"3a2b"),
(x"3752",x"3c75",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"3752",x"3c75",x"3710",x"3be0",x"b1a3",x"868d",x"3a87",x"3b59",x"376c",x"3c7b",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f"),
(x"36dc",x"3ca9",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36dc",x"3ca9",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47",x"36c4",x"3ca2",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d"),
(x"3999",x"3cac",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"3999",x"3cac",x"3710",x"b329",x"3bcb",x"868d",x"3bd9",x"3a2b",x"3994",x"3cac",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29"),
(x"3742",x"3c68",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"3742",x"3c68",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b",x"3753",x"3c6a",x"3710",x"38fe",x"ba3f",x"8000",x"3a87",x"3b4e"),
(x"36c4",x"3ca2",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36c4",x"3ca2",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d",x"36c2",x"3c9f",x"3710",x"bafe",x"b7c2",x"0000",x"3aa1",x"3a50"),
(x"3994",x"3cac",x"36da",x"b458",x"3bb2",x"068d",x"3be3",x"3a29",x"3994",x"3cac",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29",x"3985",x"3ca7",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22"),
(x"372e",x"3c68",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"372e",x"3c68",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47",x"3742",x"3c68",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b"),
(x"36c2",x"3c9f",x"36da",x"bbe7",x"b0ec",x"8000",x"3a97",x"3a50",x"36c2",x"3c9f",x"3710",x"bafe",x"b7c2",x"0000",x"3aa1",x"3a50",x"36cb",x"3c9d",x"3710",x"b86c",x"baaa",x"0000",x"3aa1",x"3a52"),
(x"3985",x"3ca7",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3985",x"3ca7",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22",x"3972",x"3ca2",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a"),
(x"3716",x"3c65",x"36da",x"32c2",x"bbd1",x"8000",x"3a7c",x"3b42",x"3716",x"3c65",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42",x"372e",x"3c68",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47"),
(x"36cb",x"3c9d",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"36cb",x"3c9d",x"3710",x"b86c",x"baaa",x"0000",x"3aa1",x"3a52",x"3705",x"3c9a",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d"),
(x"3972",x"3ca2",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3972",x"3ca2",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a",x"3963",x"3ca2",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14"),
(x"36f7",x"3c65",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"36f7",x"3c65",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c",x"3716",x"3c65",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42"),
(x"3705",x"3c9a",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"3705",x"3c9a",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d",x"3713",x"3c99",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60"),
(x"3963",x"3ca2",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"3963",x"3ca2",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14",x"395d",x"3ca4",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11"),
(x"36e3",x"3c67",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36e3",x"3c67",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38",x"36f7",x"3c65",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c"),
(x"3713",x"3c99",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3713",x"3c99",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60",x"3716",x"3c98",x"3710",x"bbad",x"3480",x"0000",x"3aa1",x"3a61"),
(x"395d",x"3ca4",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"395d",x"3ca4",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11",x"395a",x"3ca7",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e"),
(x"36df",x"3c6a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36df",x"3c6a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35",x"36e3",x"3c67",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38"),
(x"3716",x"3c98",x"36da",x"bbb8",x"b42d",x"0000",x"3a54",x"39ec",x"3716",x"3c98",x"3710",x"bbad",x"3480",x"0000",x"3a5f",x"39ec",x"3710",x"3c96",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee"),
(x"395a",x"3ca7",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"395a",x"3ca7",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e",x"3953",x"3cac",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09"),
(x"36dc",x"3c6d",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36dc",x"3c6d",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33",x"36df",x"3c6a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35"),
(x"3710",x"3c96",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"3710",x"3c96",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee",x"36f7",x"3c95",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3"),
(x"3475",x"3c8f",x"36da",x"baeb",x"3803",x"8000",x"3a6e",x"3b70",x"3475",x"3c8f",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70",x"3475",x"3c87",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77"),
(x"3953",x"3cac",x"36da",x"39a8",x"39a7",x"0a8d",x"3be3",x"3a09",x"3953",x"3cac",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09",x"393f",x"3cae",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01"),
(x"36c4",x"3c74",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36c4",x"3c74",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c",x"36dc",x"3c6d",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33"),
(x"363b",x"3c95",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"363b",x"3c95",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16",x"362c",x"3c96",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19"),
(x"3994",x"3c6b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3994",x"3c6b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b",x"3999",x"3c6a",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d"),
(x"393f",x"3cae",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"393f",x"3cae",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01",x"392f",x"3cab",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa"),
(x"36c2",x"3c77",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36c2",x"3c77",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a",x"36c4",x"3c74",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c"),
(x"36f7",x"3c95",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"36f7",x"3c95",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3",x"363b",x"3c95",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16"),
(x"3985",x"3c6f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3985",x"3c6f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25",x"3994",x"3c6b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b"),
(x"3752",x"3ca1",x"36da",x"3be0",x"31a3",x"868d",x"3a97",x"3a21",x"3752",x"3ca1",x"3710",x"3bfd",x"aac2",x"0000",x"3aa1",x"3a21",x"3754",x"3ca4",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23"),
(x"36cb",x"3c79",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"36cb",x"3c79",x"3710",x"b922",x"3a22",x"0000",x"3a87",x"3b28",x"36c2",x"3c77",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a"),
(x"362c",x"3c96",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"362c",x"3c96",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19",x"35f7",x"3c9e",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25"),
(x"3972",x"3c74",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3972",x"3c74",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d",x"3985",x"3c6f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25"),
(x"392f",x"3cab",x"36da",x"b73b",x"3b22",x"068d",x"3be3",x"39fa",x"392f",x"3cab",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa",x"3915",x"3c9e",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec"),
(x"3705",x"3c7c",x"36da",x"b676",x"3b51",x"0000",x"3a7c",x"3b1d",x"3705",x"3c7c",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d",x"36cb",x"3c79",x"3710",x"b922",x"3a22",x"0000",x"3a87",x"3b28"),
(x"35f7",x"3c9e",x"36da",x"3a05",x"3944",x"8000",x"3a54",x"3a25",x"35f7",x"3c9e",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25",x"35f1",x"3ca0",x"3710",x"3bf9",x"ad20",x"0000",x"3a5f",x"3a27"),
(x"3963",x"3c74",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"3963",x"3c74",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17",x"3972",x"3c74",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d"),
(x"3754",x"3ca4",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"3754",x"3ca4",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23",x"375f",x"3ca7",x"3710",x"3bc1",x"b3d7",x"068d",x"3aa1",x"3a26"),
(x"3713",x"3c7e",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3713",x"3c7e",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a",x"3705",x"3c7c",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d"),
(x"35f1",x"3ca0",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f1",x"3ca0",x"3710",x"3bf9",x"ad20",x"0000",x"3a5f",x"3a27",x"35f3",x"3ca2",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28"),
(x"395d",x"3c72",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"395d",x"3c72",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14",x"3963",x"3c74",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17"),
(x"3915",x"3c9e",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"3915",x"3c9e",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec",x"38f6",x"3c96",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de"),
(x"3716",x"3c7f",x"36da",x"bbad",x"b480",x"0000",x"3a7c",x"3b19",x"3716",x"3c7f",x"3710",x"bbb8",x"342d",x"0000",x"3a87",x"3b19",x"3713",x"3c7e",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a"),
(x"35f3",x"3ca2",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35f3",x"3ca2",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28",x"35fd",x"3ca5",x"3710",x"3bf0",x"aff4",x"868d",x"3a5f",x"3a2b"),
(x"395a",x"3c6f",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"395a",x"3c6f",x"3710",x"3b46",x"b6a7",x"8000",x"3a85",x"3a12",x"395d",x"3c72",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14"),
(x"38f6",x"3c96",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"38f6",x"3c96",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de",x"38d5",x"3c94",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1"),
(x"3710",x"3c80",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"3710",x"3c80",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f",x"3716",x"3c7f",x"3710",x"bbb8",x"342d",x"0000",x"3b06",x"3a11"),
(x"35fd",x"3ca5",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35fd",x"3ca5",x"3710",x"3bf0",x"aff4",x"868d",x"3a5f",x"3a2b",x"35fd",x"3ca7",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d"),
(x"3953",x"3c6a",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"3953",x"3c6a",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d",x"395a",x"3c6f",x"3710",x"3b46",x"b6a7",x"8000",x"3a85",x"3a12"),
(x"38d5",x"3c94",x"36da",x"1987",x"3c00",x"0000",x"3be3",x"39d1",x"38d5",x"3c94",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1",x"38bf",x"3c96",x"3710",x"35f3",x"3b6c",x"0000",x"3bd9",x"39c8"),
(x"36f7",x"3c81",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"36f7",x"3c81",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a",x"3710",x"3c80",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f"),
(x"35fd",x"3ca7",x"36da",x"3b87",x"3567",x"8000",x"3a54",x"3a2d",x"35fd",x"3ca7",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d",x"35f5",x"3ca8",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e"),
(x"393f",x"3c68",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"393f",x"3c68",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05",x"3953",x"3c6a",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d"),
(x"38bf",x"3c96",x"36da",x"3489",x"3bab",x"0000",x"3be3",x"39c8",x"38bf",x"3c96",x"3710",x"35f3",x"3b6c",x"0000",x"3bd9",x"39c8",x"38b2",x"3c99",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2"),
(x"362c",x"3c80",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"362c",x"3c80",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4",x"363b",x"3c81",x"3710",x"3439",x"bbb7",x"0000",x"3b06",x"39e7"),
(x"35f5",x"3ca8",x"36da",x"364b",x"3b5a",x"8000",x"3a54",x"3a2e",x"35f5",x"3ca8",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e",x"35e4",x"3ca8",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32"),
(x"392f",x"3c6b",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"392f",x"3c6b",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff",x"393f",x"3c68",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05"),
(x"38b2",x"3c99",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38b2",x"3c99",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2",x"38b0",x"3c9c",x"3710",x"3ba6",x"b4ac",x"0000",x"3bd9",x"39c0"),
(x"363b",x"3c81",x"36da",x"34bd",x"bba4",x"0000",x"3afb",x"39e7",x"363b",x"3c81",x"3710",x"3439",x"bbb7",x"0000",x"3b06",x"39e7",x"36f7",x"3c81",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a"),
(x"35e4",x"3ca8",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35e4",x"3ca8",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32",x"35d3",x"3ca7",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35"),
(x"3754",x"3c72",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"3754",x"3c72",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57",x"3752",x"3c75",x"3710",x"3be0",x"b1a3",x"868d",x"3a87",x"3b59"),
(x"38b0",x"3c9c",x"36da",x"3bfc",x"2b27",x"0000",x"3be3",x"39c0",x"38b0",x"3c9c",x"3710",x"3ba6",x"b4ac",x"0000",x"3bd9",x"39c0",x"38b2",x"3c9e",x"3710",x"399c",x"b9b3",x"8000",x"3bd9",x"39be"),
(x"35f7",x"3c78",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"35f7",x"3c78",x"3710",x"3a05",x"b944",x"8000",x"3b06",x"39d8",x"362c",x"3c80",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4"),
(x"35d3",x"3ca7",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35d3",x"3ca7",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35",x"35bd",x"3ca8",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39"),
(x"3915",x"3c79",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"3915",x"3c79",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1",x"392f",x"3c6b",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff"),
(x"38b2",x"3c9e",x"36da",x"3a58",x"b8de",x"0000",x"3a7d",x"3ac5",x"38b2",x"3c9e",x"3710",x"399c",x"b9b3",x"8000",x"3a87",x"3ac5",x"38bd",x"3ca0",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9"),
(x"35f1",x"3c76",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f1",x"3c76",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6",x"35f7",x"3c78",x"3710",x"3a05",x"b944",x"8000",x"3b06",x"39d8"),
(x"35bd",x"3ca8",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"35bd",x"3ca8",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39",x"359e",x"3ca5",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40"),
(x"375f",x"3c70",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"375f",x"3c70",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54",x"3754",x"3c72",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57"),
(x"38bd",x"3ca0",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38bd",x"3ca0",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9",x"38c9",x"3ca1",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace"),
(x"35f3",x"3c75",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35f3",x"3c75",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5",x"35f1",x"3c76",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6"),
(x"359e",x"3ca5",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"359e",x"3ca5",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40",x"358a",x"3c9f",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45"),
(x"38f6",x"3c80",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"38f6",x"3c80",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4",x"3915",x"3c79",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1"),
(x"38c9",x"3ca1",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38c9",x"3ca1",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace",x"38d4",x"3ca4",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2"),
(x"35fd",x"3c71",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35fd",x"3c71",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2",x"35f3",x"3c75",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5"),
(x"358a",x"3c9f",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"358a",x"3c9f",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45",x"3587",x"3c9a",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49"),
(x"38d5",x"3c82",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38d5",x"3c82",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7",x"38f6",x"3c80",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4"),
(x"38d4",x"3ca4",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38d4",x"3ca4",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2",x"38d9",x"3ca6",x"3710",x"3bfc",x"ab00",x"0000",x"3a87",x"3ad5"),
(x"3a26",x"3c69",x"36da",x"3bff",x"26b5",x"0000",x"39f5",x"33fa",x"3a26",x"3c69",x"3710",x"3bcf",x"2680",x"32dc",x"39f4",x"33ca",x"3a25",x"3c7f",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0"),
(x"35fd",x"3c6f",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35fd",x"3c6f",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0",x"35fd",x"3c71",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2"),
(x"3587",x"3c9a",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"3587",x"3c9a",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49",x"3593",x"3c95",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d"),
(x"38bf",x"3c80",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38bf",x"3c80",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf",x"38d5",x"3c82",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7"),
(x"38d9",x"3ca6",x"36da",x"3b88",x"b564",x"0000",x"3a7d",x"3ad5",x"38d9",x"3ca6",x"3710",x"3bfc",x"ab00",x"0000",x"3a87",x"3ad5",x"38d8",x"3ca7",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6"),
(x"35f5",x"3c6e",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35f5",x"3c6e",x"3710",x"364b",x"bb5a",x"8000",x"3b06",x"39ce",x"35fd",x"3c6f",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0"),
(x"3593",x"3c95",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3593",x"3c95",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d",x"3592",x"3c93",x"3710",x"ba08",x"3941",x"0000",x"3a5f",x"3a4f"),
(x"38b2",x"3c7d",x"36da",x"3af2",x"b7f0",x"0000",x"3a7b",x"39c9",x"38b2",x"3c7d",x"3710",x"3a0a",x"b93e",x"8000",x"3a85",x"39c9",x"38bf",x"3c80",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf"),
(x"38d8",x"3ca7",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38d8",x"3ca7",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6",x"38c7",x"3cab",x"3710",x"3649",x"3b5b",x"0000",x"3a87",x"3add"),
(x"35e4",x"3c6e",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35e4",x"3c6e",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb",x"35f5",x"3c6e",x"3710",x"364b",x"bb5a",x"8000",x"3b06",x"39ce"),
(x"3592",x"3c93",x"36da",x"bba4",x"34bb",x"0000",x"3a6e",x"3b35",x"3592",x"3c93",x"3710",x"ba08",x"3941",x"0000",x"3a79",x"3b35",x"357d",x"3c93",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39"),
(x"38b0",x"3c7b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b0",x"3c7b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d",x"38b2",x"3c7d",x"3710",x"3a0a",x"b93e",x"8000",x"3a95",x"3a50"),
(x"38c7",x"3cab",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38c7",x"3cab",x"3710",x"3649",x"3b5b",x"0000",x"3a87",x"3add",x"38b7",x"3cae",x"3710",x"32f6",x"3bce",x"0000",x"3a87",x"3ae4"),
(x"35d3",x"3c70",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35d3",x"3c70",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8",x"35e4",x"3c6e",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb"),
(x"357d",x"3c93",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"357d",x"3c93",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39",x"3555",x"3c94",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41"),
(x"38b2",x"3c79",x"36da",x"399d",x"39b3",x"8000",x"3a8a",x"3a4c",x"38b2",x"3c79",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c",x"38b0",x"3c7b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d"),
(x"38b7",x"3cae",x"36da",x"3528",x"3b92",x"0000",x"3a7d",x"3ae4",x"38b7",x"3cae",x"3710",x"32f6",x"3bce",x"0000",x"3a87",x"3ae4",x"3894",x"3caf",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1"),
(x"35bd",x"3c6e",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"35bd",x"3c6e",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3",x"35d3",x"3c70",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8"),
(x"3555",x"3c94",x"36da",x"345a",x"3bb2",x"0000",x"3a6e",x"3b41",x"3555",x"3c94",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41",x"353f",x"3c97",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46"),
(x"38bd",x"3c76",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38bd",x"3c76",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47",x"38b2",x"3c79",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c"),
(x"3894",x"3caf",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"3894",x"3caf",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1",x"3877",x"3cac",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc"),
(x"359e",x"3c71",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"359e",x"3c71",x"3710",x"b80b",x"bae7",x"868d",x"3b06",x"39bd",x"35bd",x"3c6e",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3"),
(x"353f",x"3c97",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"353f",x"3c97",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46",x"351b",x"3c9c",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e"),
(x"38c9",x"3c75",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38c9",x"3c75",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43",x"38bd",x"3c76",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47"),
(x"3877",x"3cac",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"3877",x"3cac",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc",x"386d",x"3ca8",x"3710",x"bba8",x"34a3",x"868d",x"3a87",x"3b01"),
(x"358a",x"3c77",x"36da",x"bbad",x"b482",x"868d",x"3afb",x"39b7",x"358a",x"3c77",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7",x"359e",x"3c71",x"3710",x"b80b",x"bae7",x"868d",x"3b06",x"39bd"),
(x"351b",x"3c9c",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"351b",x"3c9c",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e",x"3501",x"3c9e",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53"),
(x"38d4",x"3c73",x"36da",x"38a8",x"3a80",x"8000",x"3a8a",x"3a3e",x"38d4",x"3c73",x"3710",x"37f2",x"3af1",x"8000",x"3a95",x"3a3e",x"38c9",x"3c75",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43"),
(x"386d",x"3ca8",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"386d",x"3ca8",x"3710",x"bba8",x"34a3",x"868d",x"3a87",x"3b01",x"386c",x"3ca2",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05"),
(x"3587",x"3c7c",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"3587",x"3c7c",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3",x"358a",x"3c77",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7"),
(x"3501",x"3c9e",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"3501",x"3c9e",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53",x"34e9",x"3c9d",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57"),
(x"38d9",x"3c71",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d9",x"3c71",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c",x"38d4",x"3c73",x"3710",x"37f2",x"3af1",x"8000",x"3a95",x"3a3e"),
(x"386c",x"3ca2",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"386c",x"3ca2",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05",x"3872",x"3c9f",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08"),
(x"3593",x"3c81",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3593",x"3c81",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af",x"3587",x"3c7c",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3"),
(x"34e9",x"3c9d",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"34e9",x"3c9d",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57",x"34cb",x"3c98",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e"),
(x"38d8",x"3c6f",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38d8",x"3c6f",x"3710",x"3be4",x"b12f",x"0000",x"3a95",x"3a3b",x"38d9",x"3c71",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c"),
(x"3872",x"3c9f",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"3872",x"3c9f",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08",x"3885",x"3c9a",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10"),
(x"3592",x"3c83",x"36da",x"ba08",x"b941",x"8000",x"3afb",x"39ae",x"3592",x"3c83",x"3710",x"bba4",x"b4bb",x"0000",x"3b06",x"39ae",x"3593",x"3c81",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af"),
(x"34cb",x"3c98",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34cb",x"3c98",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e",x"34bb",x"3c97",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61"),
(x"38c7",x"3c6c",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38c7",x"3c6c",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34",x"38d8",x"3c6f",x"3710",x"3be4",x"b12f",x"0000",x"3a95",x"3a3b"),
(x"3885",x"3c9a",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"3885",x"3c9a",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10",x"388c",x"3c98",x"3710",x"bbfd",x"a9ab",x"0000",x"3a87",x"3b13"),
(x"357d",x"3c83",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"357d",x"3c83",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae",x"3592",x"3c83",x"3710",x"bba4",x"b4bb",x"0000",x"3a79",x"3bb2"),
(x"34bb",x"3c97",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"34bb",x"3c97",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61",x"349b",x"3c96",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67"),
(x"38b7",x"3c68",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"38b7",x"3c68",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d",x"38c7",x"3c6c",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34"),
(x"388c",x"3c98",x"36da",x"bb54",x"b669",x"0000",x"3a97",x"39c6",x"388c",x"3c98",x"3710",x"bbfd",x"a9ab",x"0000",x"3aa1",x"39c6",x"388c",x"3c96",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8"),
(x"3555",x"3c82",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"3555",x"3c82",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6",x"357d",x"3c83",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae"),
(x"349b",x"3c96",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"349b",x"3c96",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67",x"3485",x"3c94",x"3710",x"b92c",x"3a1a",x"868d",x"3a79",x"3b6c"),
(x"3894",x"3c67",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"3894",x"3c67",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20",x"38b7",x"3c68",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d"),
(x"388c",x"3c96",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"388c",x"3c96",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8",x"3885",x"3c95",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca"),
(x"353f",x"3c7f",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"353f",x"3c7f",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2",x"3555",x"3c82",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6"),
(x"3485",x"3c94",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"3485",x"3c94",x"3710",x"b92c",x"3a1a",x"868d",x"3a79",x"3b6c",x"3475",x"3c8f",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70"),
(x"3877",x"3c6a",x"36da",x"b8aa",x"ba7f",x"8000",x"3a8a",x"3a15",x"3877",x"3c6a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15",x"3894",x"3c67",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20"),
(x"3760",x"3ca9",x"36da",x"3bfa",x"2cac",x"068d",x"3a97",x"3a28",x"3760",x"3ca9",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28",x"3753",x"3cad",x"3710",x"37e4",x"3af5",x"868d",x"3aa1",x"3a2b"),
(x"3a2d",x"3c81",x"36da",x"3bfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"3a2d",x"3c81",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a2f",x"3c96",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"351b",x"3c7a",x"36da",x"350e",x"bb96",x"0000",x"3a6e",x"3b9a",x"351b",x"3c7a",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a",x"353f",x"3c7f",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2"),
(x"3a27",x"3cae",x"36da",x"a3ae",x"3bff",x"0000",x"3be3",x"3a63",x"3a27",x"3cae",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63",x"39f5",x"3cae",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f"),
(x"386d",x"3c6f",x"36da",x"bba8",x"b4a3",x"068d",x"3a8a",x"3a10",x"386d",x"3c6f",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10",x"3877",x"3c6a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15"),
(x"3885",x"3c95",x"36da",x"b304",x"3bce",x"0000",x"3a97",x"39ca",x"3885",x"3c95",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca",x"382a",x"3c96",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed"),
(x"3501",x"3c78",x"36da",x"ada8",x"bbf8",x"0000",x"3a6e",x"3b94",x"3501",x"3c78",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94",x"351b",x"3c7a",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a"),
(x"386c",x"3c74",x"36da",x"bb38",x"36e2",x"068d",x"3a8a",x"3a0c",x"386c",x"3c74",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c",x"386d",x"3c6f",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10"),
(x"382a",x"3c96",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"382a",x"3c96",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed",x"3813",x"3c97",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5"),
(x"3a25",x"3c7f",x"36da",x"367a",x"bb50",x"0000",x"3bc0",x"3984",x"3a25",x"3c7f",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c",x"3a2d",x"3c81",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a"),
(x"3a1f",x"3c7f",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a25",x"3c7f",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0",x"3a20",x"3c69",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa"),
(x"3a18",x"3c7f",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a1f",x"3c7f",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a19",x"3c69",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392"),
(x"3a10",x"3c7f",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a18",x"3c7f",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a14",x"3c69",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387"),
(x"3a09",x"3c7f",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a10",x"3c7f",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a0d",x"3c69",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b"),
(x"3a09",x"3c81",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a09",x"3c7f",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"3a03",x"3c81",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bbd",x"39a7"),
(x"3a09",x"3c7f",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"3a09",x"3c81",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a10",x"3c7f",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b"),
(x"3a08",x"3c96",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a09",x"3c81",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1",x"3a04",x"3c96",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7"),
(x"3a03",x"3c81",x"370e",x"bbc2",x"ab4f",x"338c",x"3bf9",x"39fa",x"3a04",x"3c96",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7",x"3a09",x"3c81",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1"),
(x"3a09",x"3c81",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1",x"3a08",x"3c96",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a11",x"3c81",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed"),
(x"3a11",x"3c81",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed",x"3a0f",x"3c96",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a19",x"3c82",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a17",x"3c96",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3be8",x"39eb",x"3a1d",x"3c96",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a19",x"3c82",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a1d",x"3c96",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a24",x"3c96",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a21",x"3c81",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6"),
(x"3a24",x"3c96",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a2a",x"3c96",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a25",x"3c81",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3"),
(x"3a1f",x"3c7f",x"3733",x"3800",x"ba99",x"3436",x"3bb7",x"3993",x"3a25",x"3c81",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a25",x"3c7f",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c"),
(x"3a02",x"3c68",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352",x"3a09",x"3c7f",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a07",x"3c69",x"373c",x"bac4",x"2853",x"3841",x"39f2",x"336a"),
(x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e",x"3a09",x"3c7f",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a02",x"3c68",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352"),
(x"3a10",x"3c7f",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b",x"3a11",x"3c81",x"374a",x"b547",x"b37e",x"3b50",x"3bb7",x"399b",x"3a18",x"3c7f",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998"),
(x"3a1f",x"3c7f",x"3733",x"3800",x"ba99",x"3436",x"3bb7",x"3993",x"3a18",x"3c7f",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998",x"3a21",x"3c81",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a2f",x"3c96",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"3861",x"3a2a",x"3c96",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a26",x"3c97",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3a2a",x"3c96",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a24",x"3c96",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a20",x"3c97",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b"),
(x"3a24",x"3c96",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a1d",x"3c96",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e",x"3a1a",x"3c97",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e"),
(x"3a17",x"3c96",x"3751",x"2fda",x"39a6",x"3994",x"3b24",x"3871",x"3a0f",x"3c96",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a15",x"3c97",x"374b",x"aaab",x"39a7",x"39a5",x"3b22",x"3871"),
(x"3a0f",x"3c96",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a08",x"3c96",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a0f",x"3c97",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873"),
(x"3a08",x"3c96",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a04",x"3c96",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879",x"3a09",x"3c98",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875"),
(x"39fb",x"3c97",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"3a02",x"3c96",x"3711",x"315a",x"2baa",x"3bdf",x"3a19",x"3349",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3a20",x"3c97",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a24",x"3cae",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a26",x"3c97",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4"),
(x"3a21",x"3cae",x"373a",x"3acd",x"a5ae",x"3834",x"3a2d",x"33a3",x"3a20",x"3c97",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a1a",x"3cae",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a1a",x"3c97",x"3746",x"38a5",x"a839",x"3a81",x"3a1a",x"338e",x"3a15",x"3c97",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a1a",x"3cae",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a15",x"3c97",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a0f",x"3c97",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a14",x"3cae",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385"),
(x"3a0f",x"3c97",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a09",x"3c98",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a0d",x"3cad",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378"),
(x"3a07",x"3cae",x"373c",x"baa1",x"a6bb",x"3879",x"3a2d",x"3366",x"3a09",x"3c98",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a00",x"3cad",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c"),
(x"3a00",x"3cad",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c",x"3a01",x"3c97",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"39fc",x"3cae",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340"),
(x"3475",x"3c87",x"3710",x"0000",x"0000",x"3c00",x"3a0c",x"2451",x"3475",x"3c8f",x"3710",x"0000",x"0000",x"3c00",x"3a13",x"2451",x"3485",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"3485",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1",x"3485",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"349b",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f"),
(x"349b",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f",x"349b",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"34bb",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643"),
(x"34cb",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"26b3",x"34bb",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643",x"34cb",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"34cb",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"26b3",x"34cb",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3",x"34e9",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b"),
(x"3501",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"281a",x"34e9",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b",x"3501",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"3501",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"281a",x"3501",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a",x"351b",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878"),
(x"351b",x"3c7a",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878",x"351b",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"353f",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"353f",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb",x"353f",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"3555",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949"),
(x"3555",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949",x"3555",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"357d",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"357d",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7",x"357d",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"3592",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"36f7",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2d8d",x"363b",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"36f7",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"363b",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2c3f",x"363b",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"362c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"362c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23",x"362c",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"3592",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"35e4",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35f5",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b84",x"35fd",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"35d3",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35e4",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35f3",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"35bd",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35d3",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35f1",x"3ca0",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"35fd",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2ba0",x"35f5",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b84",x"35fd",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"35fd",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0",x"35e4",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35f3",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"35f3",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d",x"35d3",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35f1",x"3c76",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"35f1",x"3c76",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76",x"35bd",x"3c6e",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"359e",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"35bd",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"36f7",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2d8d",x"36f7",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d",x"3710",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"380a",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2f8b",x"380a",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b",x"37b8",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"37a8",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ec9",x"37b8",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7",x"37a8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"37a8",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ec9",x"37a8",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9",x"378c",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"378c",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97",x"378c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"376c",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"3752",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"376c",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e",x"3752",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"36e3",x"3caf",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"2d6a",x"36f7",x"3cb2",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e",x"36df",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"36df",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63",x"3716",x"3cb1",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"36dc",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"36e3",x"3c67",x"3710",x"0000",x"0000",x"3c00",x"39f0",x"2d6a",x"36df",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"36f7",x"3c65",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"36df",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"36dc",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"3716",x"3c65",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"3760",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2e49",x"3753",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2e32",x"375f",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"375f",x"3c70",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47",x"3742",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"3754",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"3742",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"3753",x"3cad",x"3710",x"0000",x"0000",x"3c00",x"3a2c",x"2e32",x"375f",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"372e",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0",x"3742",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"3754",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"3705",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36cb",x"3c9d",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2d40",x"36c4",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"36c2",x"3c77",x"3710",x"0000",x"0000",x"3c00",x"39fe",x"2d2f",x"36cb",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"2d40",x"36c4",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"36c4",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33",x"3705",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"36dc",x"3c6d",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"3713",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3705",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36dc",x"3ca9",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"3754",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33",x"3713",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"372e",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"3754",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33",x"372e",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3713",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"3716",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5",x"3713",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3752",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"3754",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33",x"3713",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"3752",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"3716",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5",x"3710",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb",x"3716",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"3716",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5",x"3752",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"3716",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"380a",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2f8b",x"3813",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"380a",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"3813",x"3c97",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"382a",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3813",x"3c7f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"382a",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2ffc",x"382a",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3885",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"3885",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30a2",x"388c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"3885",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"38d5",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130",x"38bf",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38d5",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130"),
(x"38bf",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"3109",x"38bf",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38b2",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"38b2",x"3c99",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1",x"38b2",x"3c7d",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b0",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38b0",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed",x"38b0",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"388c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"386c",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3075",x"3872",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"386d",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3076"),
(x"3872",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"3885",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"3877",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088"),
(x"386c",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3075",x"386d",x"3ca8",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"3076",x"3872",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080"),
(x"3872",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080",x"3877",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3885",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"3885",x"3c9a",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2",x"3894",x"3caf",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"388c",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"3885",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"388c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"3894",x"3c67",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"38d9",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"3136",x"38d8",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3135",x"38d4",x"3c73",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d"),
(x"38c7",x"3cab",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38d8",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3135",x"38d4",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d"),
(x"38b7",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38c7",x"3cab",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38c9",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a"),
(x"38d4",x"3c73",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d",x"38c7",x"3c6c",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38c9",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a"),
(x"38b2",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"388c",x"3c7e",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"38b0",x"3c7b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"388c",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"388c",x"3c98",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae",x"38b0",x"3c9c",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38c9",x"3c75",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a",x"38b7",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38bd",x"3c76",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3107"),
(x"38d5",x"3c94",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130",x"38f6",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"38d5",x"3c82",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130"),
(x"38f6",x"3c96",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"3915",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"38f6",x"3c80",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b"),
(x"3915",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"31a2",x"3915",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"392f",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"392f",x"3cab",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"31d0",x"393f",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"392f",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"393f",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"3953",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"393f",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"3953",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"395a",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"3953",x"3c6a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211"),
(x"395a",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"395d",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"395a",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d"),
(x"395d",x"3c72",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"3222",x"395d",x"3ca4",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"3963",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3963",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"322d",x"3972",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3963",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3972",x"3ca2",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3985",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3972",x"3c74",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248"),
(x"3985",x"3c6f",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"3269",x"3985",x"3ca7",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3994",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3994",x"3cac",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3284",x"3999",x"3cac",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"3994",x"3c6b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3999",x"3c6a",x"3710",x"96f6",x"9f93",x"3c00",x"39f3",x"328d",x"3999",x"3cac",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39fc",x"3c80",x"3713",x"ac10",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3999",x"3cac",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39f5",x"3cae",x"3710",x"b60a",x"25b5",x"3b67",x"3a2d",x"3331",x"39fb",x"3c97",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d"),
(x"3a14",x"3cae",x"374f",x"a8f4",x"3bfa",x"ac2a",x"3bcd",x"3a5c",x"3a0d",x"3cad",x"374b",x"a412",x"3bfd",x"2963",x"3bce",x"3a59",x"3a1a",x"3cae",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e"),
(x"3a1a",x"3cae",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e",x"3a07",x"3cae",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a21",x"3cae",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60"),
(x"3a21",x"3cae",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60",x"3a00",x"3cad",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"3a24",x"3cae",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62"),
(x"3a24",x"3cae",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62",x"39fc",x"3cae",x"3718",x"135f",x"3bfd",x"299e",x"3bd8",x"3a52",x"3a27",x"3cae",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63"),
(x"3a14",x"3c69",x"374e",x"a81b",x"bbe6",x"b0f3",x"3a92",x"3a5c",x"3a19",x"3c69",x"3749",x"209b",x"bc00",x"135f",x"3a90",x"3a5e",x"3a0d",x"3c69",x"374b",x"1481",x"bbff",x"269a",x"3a91",x"3a59"),
(x"3a19",x"3c69",x"3749",x"209b",x"bc00",x"135f",x"3a90",x"3a5e",x"3a20",x"3c69",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a07",x"3c69",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a8e",x"3a57"),
(x"3a20",x"3c69",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a26",x"3c69",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63",x"3a02",x"3c68",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55"),
(x"3501",x"3c78",x"36da",x"ada8",x"bbf8",x"0000",x"3a6e",x"3b94",x"34e9",x"3c7a",x"36da",x"b699",x"bb49",x"0000",x"3a6e",x"3b90",x"3501",x"3c78",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94"),
(x"386c",x"3c74",x"36da",x"bb38",x"36e2",x"068d",x"3a8a",x"3a0c",x"3872",x"3c78",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"386c",x"3c74",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c"),
(x"380a",x"3c97",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"3813",x"3c97",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"380a",x"3c97",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9"),
(x"34e9",x"3c7a",x"36da",x"b699",x"bb49",x"0000",x"3a6e",x"3b90",x"34cb",x"3c7e",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34e9",x"3c7a",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90"),
(x"3a26",x"3c69",x"36da",x"1e3f",x"bc00",x"0000",x"3a7b",x"3a63",x"39fc",x"3c69",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"3a26",x"3c69",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63"),
(x"3872",x"3c78",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"3885",x"3c7c",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"3872",x"3c78",x"3710",x"b9d1",x"397d",x"0000",x"3a95",x"3a08"),
(x"3760",x"3ca9",x"36da",x"3bfa",x"2cac",x"068d",x"3a97",x"3a28",x"375f",x"3ca7",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"3760",x"3ca9",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28"),
(x"34cb",x"3c7e",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34bb",x"3c7f",x"36da",x"b13f",x"bbe4",x"0000",x"3a6e",x"3b86",x"34cb",x"3c7e",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89"),
(x"3885",x"3c7c",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"388c",x"3c7e",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"3885",x"3c7c",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00"),
(x"37b8",x"3c94",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"380a",x"3c97",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"37b8",x"3c94",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b"),
(x"34bb",x"3c7f",x"36da",x"b13f",x"bbe4",x"0000",x"3a6e",x"3b86",x"349b",x"3c80",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"34bb",x"3c7f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86"),
(x"388c",x"3c7e",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"388c",x"3c80",x"36da",x"b967",x"b9e6",x"0000",x"3a8a",x"39fb",x"388c",x"3c7e",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd"),
(x"37a8",x"3c95",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"37b8",x"3c94",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"37a8",x"3c95",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e"),
(x"349b",x"3c80",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"3485",x"3c82",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"349b",x"3c80",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80"),
(x"388c",x"3c80",x"36da",x"b967",x"b9e6",x"0000",x"3a7c",x"3bb2",x"3885",x"3c81",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"388c",x"3c80",x"3710",x"bb52",x"b671",x"0000",x"3a87",x"3bb2"),
(x"378c",x"3c99",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"37a8",x"3c95",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"378c",x"3c99",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14"),
(x"3a26",x"3c97",x"36da",x"3311",x"3bcd",x"0000",x"3b16",x"385d",x"3a2f",x"3c96",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"385a",x"3a26",x"3c97",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3485",x"3c82",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"3475",x"3c87",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3485",x"3c82",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b"),
(x"3760",x"3c6d",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"3753",x"3c6a",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3760",x"3c6d",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52"),
(x"376c",x"3c9c",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"378c",x"3c99",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"376c",x"3c9c",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a"),
(x"3885",x"3c81",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"382a",x"3c81",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"3885",x"3c81",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf"),
(x"3752",x"3ca1",x"36da",x"3be0",x"31a3",x"868d",x"3a97",x"3a21",x"376c",x"3c9c",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"3752",x"3ca1",x"3710",x"3bfd",x"aac2",x"0000",x"3aa1",x"3a21"),
(x"39fc",x"3c69",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"3999",x"3c6a",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"39fc",x"3c69",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53"),
(x"382a",x"3c81",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"3813",x"3c7f",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"382a",x"3c81",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d"),
(x"3742",x"3cae",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"3753",x"3cad",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3742",x"3cae",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f"),
(x"3813",x"3c7f",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"380a",x"3c7f",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"3813",x"3c7f",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84"),
(x"372e",x"3cae",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"3742",x"3cae",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"372e",x"3cae",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32"),
(x"375f",x"3c70",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"3760",x"3c6d",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"375f",x"3c70",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54"),
(x"3716",x"3cb1",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"372e",x"3cae",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"3716",x"3cb1",x"3710",x"32c2",x"3bd1",x"0000",x"3aa1",x"3a37"),
(x"380a",x"3c7f",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"37b8",x"3c82",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"380a",x"3c7f",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81"),
(x"36f7",x"3cb2",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"3716",x"3cb1",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"36f7",x"3cb2",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d"),
(x"37b8",x"3c82",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"37a8",x"3c82",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"37b8",x"3c82",x"3710",x"2df5",x"bbf7",x"0000",x"3a87",x"3b6f"),
(x"36e3",x"3caf",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36f7",x"3cb2",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"36e3",x"3caf",x"3710",x"bb17",x"3766",x"068d",x"3aa1",x"3a41"),
(x"37a8",x"3c82",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"378c",x"3c7e",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"37a8",x"3c82",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c"),
(x"36df",x"3cac",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36e3",x"3caf",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36df",x"3cac",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44"),
(x"378c",x"3c7e",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"376c",x"3c7b",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"378c",x"3c7e",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66"),
(x"36dc",x"3ca9",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36df",x"3cac",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36dc",x"3ca9",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47"),
(x"3a27",x"3cae",x"36da",x"3bff",x"a4d0",x"0000",x"3a2c",x"33f9",x"3a26",x"3c97",x"36da",x"3bff",x"a4d0",x"0000",x"3a18",x"33f3",x"3a27",x"3cae",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9"),
(x"3999",x"3cac",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"39f5",x"3cae",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"3999",x"3cac",x"3710",x"b329",x"3bcb",x"868d",x"3bd9",x"3a2b"),
(x"376c",x"3c7b",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"3752",x"3c75",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"376c",x"3c7b",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f"),
(x"36c4",x"3ca2",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36dc",x"3ca9",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36c4",x"3ca2",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d"),
(x"3994",x"3cac",x"36da",x"b458",x"3bb2",x"068d",x"3be3",x"3a29",x"3999",x"3cac",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"3994",x"3cac",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29"),
(x"3753",x"3c6a",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3742",x"3c68",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"3753",x"3c6a",x"3710",x"38fe",x"ba3f",x"8000",x"3a87",x"3b4e"),
(x"36c2",x"3c9f",x"36da",x"bbe7",x"b0ec",x"8000",x"3a97",x"3a50",x"36c4",x"3ca2",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36c2",x"3c9f",x"3710",x"bafe",x"b7c2",x"0000",x"3aa1",x"3a50"),
(x"3985",x"3ca7",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3994",x"3cac",x"36da",x"b458",x"3bb2",x"068d",x"3be3",x"3a29",x"3985",x"3ca7",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22"),
(x"3742",x"3c68",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"372e",x"3c68",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"3742",x"3c68",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b"),
(x"36cb",x"3c9d",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"36c2",x"3c9f",x"36da",x"bbe7",x"b0ec",x"8000",x"3a97",x"3a50",x"36cb",x"3c9d",x"3710",x"b86c",x"baaa",x"0000",x"3aa1",x"3a52"),
(x"3972",x"3ca2",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3985",x"3ca7",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3972",x"3ca2",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a"),
(x"372e",x"3c68",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"3716",x"3c65",x"36da",x"32c2",x"bbd1",x"8000",x"3a7c",x"3b42",x"372e",x"3c68",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47"),
(x"3705",x"3c9a",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"36cb",x"3c9d",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"3705",x"3c9a",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d"),
(x"3963",x"3ca2",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"3972",x"3ca2",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3963",x"3ca2",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14"),
(x"3716",x"3c65",x"36da",x"32c2",x"bbd1",x"8000",x"3a7c",x"3b42",x"36f7",x"3c65",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"3716",x"3c65",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42"),
(x"3713",x"3c99",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3705",x"3c9a",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"3713",x"3c99",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60"),
(x"395d",x"3ca4",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"3963",x"3ca2",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"395d",x"3ca4",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11"),
(x"36f7",x"3c65",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"36e3",x"3c67",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36f7",x"3c65",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c"),
(x"3716",x"3c98",x"36da",x"bbb8",x"b42d",x"0000",x"3a97",x"3a61",x"3713",x"3c99",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3716",x"3c98",x"3710",x"bbad",x"3480",x"0000",x"3aa1",x"3a61"),
(x"395a",x"3ca7",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"395d",x"3ca4",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"395a",x"3ca7",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e"),
(x"36e3",x"3c67",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36df",x"3c6a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36e3",x"3c67",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38"),
(x"3710",x"3c96",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"3716",x"3c98",x"36da",x"bbb8",x"b42d",x"0000",x"3a54",x"39ec",x"3710",x"3c96",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee"),
(x"3953",x"3cac",x"36da",x"39a8",x"39a7",x"0a8d",x"3be3",x"3a09",x"395a",x"3ca7",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"3953",x"3cac",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09"),
(x"36df",x"3c6a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36dc",x"3c6d",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36df",x"3c6a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35"),
(x"36f7",x"3c95",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"3710",x"3c96",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"36f7",x"3c95",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3"),
(x"3475",x"3c87",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3475",x"3c8f",x"36da",x"baeb",x"3803",x"8000",x"3a6e",x"3b70",x"3475",x"3c87",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77"),
(x"393f",x"3cae",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"3953",x"3cac",x"36da",x"39a8",x"39a7",x"0a8d",x"3be3",x"3a09",x"393f",x"3cae",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01"),
(x"36dc",x"3c6d",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36c4",x"3c74",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36dc",x"3c6d",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33"),
(x"362c",x"3c96",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"363b",x"3c95",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"362c",x"3c96",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19"),
(x"3999",x"3c6a",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"3994",x"3c6b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3999",x"3c6a",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d"),
(x"392f",x"3cab",x"36da",x"b73b",x"3b22",x"068d",x"3be3",x"39fa",x"393f",x"3cae",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"392f",x"3cab",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa"),
(x"36c4",x"3c74",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36c2",x"3c77",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36c4",x"3c74",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c"),
(x"363b",x"3c95",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"36f7",x"3c95",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"363b",x"3c95",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16"),
(x"3994",x"3c6b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3985",x"3c6f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3994",x"3c6b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b"),
(x"3754",x"3ca4",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"3752",x"3ca1",x"36da",x"3be0",x"31a3",x"868d",x"3a97",x"3a21",x"3754",x"3ca4",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23"),
(x"36c2",x"3c77",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36cb",x"3c79",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"36c2",x"3c77",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a"),
(x"35f7",x"3c9e",x"36da",x"3a05",x"3944",x"8000",x"3a54",x"3a25",x"362c",x"3c96",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"35f7",x"3c9e",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25"),
(x"3985",x"3c6f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3972",x"3c74",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3985",x"3c6f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25"),
(x"3915",x"3c9e",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"392f",x"3cab",x"36da",x"b73b",x"3b22",x"068d",x"3be3",x"39fa",x"3915",x"3c9e",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec"),
(x"36cb",x"3c79",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"3705",x"3c7c",x"36da",x"b676",x"3b51",x"0000",x"3a7c",x"3b1d",x"36cb",x"3c79",x"3710",x"b922",x"3a22",x"0000",x"3a87",x"3b28"),
(x"35f1",x"3ca0",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f7",x"3c9e",x"36da",x"3a05",x"3944",x"8000",x"3a54",x"3a25",x"35f1",x"3ca0",x"3710",x"3bf9",x"ad20",x"0000",x"3a5f",x"3a27"),
(x"3972",x"3c74",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3963",x"3c74",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"3972",x"3c74",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d"),
(x"375f",x"3ca7",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"3754",x"3ca4",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"375f",x"3ca7",x"3710",x"3bc1",x"b3d7",x"068d",x"3aa1",x"3a26"),
(x"3705",x"3c7c",x"36da",x"b676",x"3b51",x"0000",x"3a7c",x"3b1d",x"3713",x"3c7e",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3705",x"3c7c",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d"),
(x"35f3",x"3ca2",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35f1",x"3ca0",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f3",x"3ca2",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28"),
(x"3963",x"3c74",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"395d",x"3c72",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"3963",x"3c74",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17"),
(x"38f6",x"3c96",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"3915",x"3c9e",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"38f6",x"3c96",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de"),
(x"3713",x"3c7e",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3716",x"3c7f",x"36da",x"bbad",x"b480",x"0000",x"3a7c",x"3b19",x"3713",x"3c7e",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a"),
(x"35fd",x"3ca5",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35f3",x"3ca2",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35fd",x"3ca5",x"3710",x"3bf0",x"aff4",x"868d",x"3a5f",x"3a2b"),
(x"395d",x"3c72",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"395a",x"3c6f",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"395d",x"3c72",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14"),
(x"38d5",x"3c94",x"36da",x"1987",x"3c00",x"0000",x"3be3",x"39d1",x"38f6",x"3c96",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"38d5",x"3c94",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1"),
(x"3716",x"3c7f",x"36da",x"bbad",x"b480",x"0000",x"3afb",x"3a11",x"3710",x"3c80",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"3716",x"3c7f",x"3710",x"bbb8",x"342d",x"0000",x"3b06",x"3a11"),
(x"35fd",x"3ca7",x"36da",x"3b87",x"3567",x"8000",x"3a54",x"3a2d",x"35fd",x"3ca5",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35fd",x"3ca7",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d"),
(x"395a",x"3c6f",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"3953",x"3c6a",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"395a",x"3c6f",x"3710",x"3b46",x"b6a7",x"8000",x"3a85",x"3a12"),
(x"38bf",x"3c96",x"36da",x"3489",x"3bab",x"0000",x"3be3",x"39c8",x"38d5",x"3c94",x"36da",x"1987",x"3c00",x"0000",x"3be3",x"39d1",x"38bf",x"3c96",x"3710",x"35f3",x"3b6c",x"0000",x"3bd9",x"39c8"),
(x"3710",x"3c80",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"36f7",x"3c81",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"3710",x"3c80",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f"),
(x"35f5",x"3ca8",x"36da",x"364b",x"3b5a",x"8000",x"3a54",x"3a2e",x"35fd",x"3ca7",x"36da",x"3b87",x"3567",x"8000",x"3a54",x"3a2d",x"35f5",x"3ca8",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e"),
(x"3953",x"3c6a",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"393f",x"3c68",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"3953",x"3c6a",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d"),
(x"38b2",x"3c99",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38bf",x"3c96",x"36da",x"3489",x"3bab",x"0000",x"3be3",x"39c8",x"38b2",x"3c99",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2"),
(x"363b",x"3c81",x"36da",x"34bd",x"bba4",x"0000",x"3afb",x"39e7",x"362c",x"3c80",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"363b",x"3c81",x"3710",x"3439",x"bbb7",x"0000",x"3b06",x"39e7"),
(x"35e4",x"3ca8",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35f5",x"3ca8",x"36da",x"364b",x"3b5a",x"8000",x"3a54",x"3a2e",x"35e4",x"3ca8",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32"),
(x"393f",x"3c68",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"392f",x"3c6b",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"393f",x"3c68",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05"),
(x"38b0",x"3c9c",x"36da",x"3bfc",x"2b27",x"0000",x"3be3",x"39c0",x"38b2",x"3c99",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38b0",x"3c9c",x"3710",x"3ba6",x"b4ac",x"0000",x"3bd9",x"39c0"),
(x"36f7",x"3c81",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"363b",x"3c81",x"36da",x"34bd",x"bba4",x"0000",x"3afb",x"39e7",x"36f7",x"3c81",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a"),
(x"35d3",x"3ca7",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35e4",x"3ca8",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35d3",x"3ca7",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35"),
(x"3752",x"3c75",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"3754",x"3c72",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"3752",x"3c75",x"3710",x"3be0",x"b1a3",x"868d",x"3a87",x"3b59"),
(x"38b2",x"3c9e",x"36da",x"3a58",x"b8de",x"0000",x"3be3",x"39be",x"38b0",x"3c9c",x"36da",x"3bfc",x"2b27",x"0000",x"3be3",x"39c0",x"38b2",x"3c9e",x"3710",x"399c",x"b9b3",x"8000",x"3bd9",x"39be"),
(x"362c",x"3c80",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"35f7",x"3c78",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"362c",x"3c80",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4"),
(x"35bd",x"3ca8",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"35d3",x"3ca7",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35bd",x"3ca8",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39"),
(x"392f",x"3c6b",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"3915",x"3c79",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"392f",x"3c6b",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff"),
(x"38bd",x"3ca0",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38b2",x"3c9e",x"36da",x"3a58",x"b8de",x"0000",x"3a7d",x"3ac5",x"38bd",x"3ca0",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9"),
(x"35f7",x"3c78",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"35f1",x"3c76",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f7",x"3c78",x"3710",x"3a05",x"b944",x"8000",x"3b06",x"39d8"),
(x"359e",x"3ca5",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"35bd",x"3ca8",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"359e",x"3ca5",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40"),
(x"3754",x"3c72",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"375f",x"3c70",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"3754",x"3c72",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57"),
(x"38c9",x"3ca1",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38bd",x"3ca0",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38c9",x"3ca1",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace"),
(x"35f1",x"3c76",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f3",x"3c75",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35f1",x"3c76",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6"),
(x"358a",x"3c9f",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"359e",x"3ca5",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"358a",x"3c9f",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45"),
(x"3915",x"3c79",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"38f6",x"3c80",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"3915",x"3c79",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1"),
(x"38d4",x"3ca4",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38c9",x"3ca1",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38d4",x"3ca4",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2"),
(x"35f3",x"3c75",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35fd",x"3c71",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35f3",x"3c75",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5"),
(x"3587",x"3c9a",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"358a",x"3c9f",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"3587",x"3c9a",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49"),
(x"38f6",x"3c80",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"38d5",x"3c82",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38f6",x"3c80",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4"),
(x"38d9",x"3ca6",x"36da",x"3b88",x"b564",x"0000",x"3a7d",x"3ad5",x"38d4",x"3ca4",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38d9",x"3ca6",x"3710",x"3bfc",x"ab00",x"0000",x"3a87",x"3ad5"),
(x"3a25",x"3c7f",x"36da",x"3bff",x"26b5",x"0000",x"3a09",x"33f0",x"3a26",x"3c69",x"36da",x"3bff",x"26b5",x"0000",x"39f5",x"33fa",x"3a25",x"3c7f",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0"),
(x"35fd",x"3c71",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35fd",x"3c6f",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35fd",x"3c71",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2"),
(x"3593",x"3c95",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3587",x"3c9a",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"3593",x"3c95",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d"),
(x"38d5",x"3c82",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38bf",x"3c80",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38d5",x"3c82",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7"),
(x"38d8",x"3ca7",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38d9",x"3ca6",x"36da",x"3b88",x"b564",x"0000",x"3a7d",x"3ad5",x"38d8",x"3ca7",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6"),
(x"35fd",x"3c6f",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35f5",x"3c6e",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35fd",x"3c6f",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0"),
(x"3592",x"3c93",x"36da",x"bba4",x"34bb",x"0000",x"3a54",x"3a4f",x"3593",x"3c95",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3592",x"3c93",x"3710",x"ba08",x"3941",x"0000",x"3a5f",x"3a4f"),
(x"38bf",x"3c80",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38b2",x"3c7d",x"36da",x"3af2",x"b7f0",x"0000",x"3a7b",x"39c9",x"38bf",x"3c80",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf"),
(x"38c7",x"3cab",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38d8",x"3ca7",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38c7",x"3cab",x"3710",x"3649",x"3b5b",x"0000",x"3a87",x"3add"),
(x"35f5",x"3c6e",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35e4",x"3c6e",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35f5",x"3c6e",x"3710",x"364b",x"bb5a",x"8000",x"3b06",x"39ce"),
(x"357d",x"3c93",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"3592",x"3c93",x"36da",x"bba4",x"34bb",x"0000",x"3a6e",x"3b35",x"357d",x"3c93",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39"),
(x"38b2",x"3c7d",x"36da",x"3af2",x"b7f0",x"0000",x"3a8a",x"3a50",x"38b0",x"3c7b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b2",x"3c7d",x"3710",x"3a0a",x"b93e",x"8000",x"3a95",x"3a50"),
(x"38b7",x"3cae",x"36da",x"3528",x"3b92",x"0000",x"3a7d",x"3ae4",x"38c7",x"3cab",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38b7",x"3cae",x"3710",x"32f6",x"3bce",x"0000",x"3a87",x"3ae4"),
(x"35e4",x"3c6e",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35d3",x"3c70",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35e4",x"3c6e",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb"),
(x"3555",x"3c94",x"36da",x"345a",x"3bb2",x"0000",x"3a6e",x"3b41",x"357d",x"3c93",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"3555",x"3c94",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41"),
(x"38b0",x"3c7b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b2",x"3c79",x"36da",x"399d",x"39b3",x"8000",x"3a8a",x"3a4c",x"38b0",x"3c7b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d"),
(x"3894",x"3caf",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"38b7",x"3cae",x"36da",x"3528",x"3b92",x"0000",x"3a7d",x"3ae4",x"3894",x"3caf",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1"),
(x"35d3",x"3c70",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35bd",x"3c6e",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"35d3",x"3c70",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8"),
(x"353f",x"3c97",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"3555",x"3c94",x"36da",x"345a",x"3bb2",x"0000",x"3a6e",x"3b41",x"353f",x"3c97",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46"),
(x"38b2",x"3c79",x"36da",x"399d",x"39b3",x"8000",x"3a8a",x"3a4c",x"38bd",x"3c76",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38b2",x"3c79",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c"),
(x"3877",x"3cac",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"3894",x"3caf",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"3877",x"3cac",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc"),
(x"35bd",x"3c6e",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"359e",x"3c71",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"35bd",x"3c6e",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3"),
(x"351b",x"3c9c",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"353f",x"3c97",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"351b",x"3c9c",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e"),
(x"38bd",x"3c76",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38c9",x"3c75",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38bd",x"3c76",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47"),
(x"386d",x"3ca8",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"3877",x"3cac",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"386d",x"3ca8",x"3710",x"bba8",x"34a3",x"868d",x"3a87",x"3b01"),
(x"359e",x"3c71",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"358a",x"3c77",x"36da",x"bbad",x"b482",x"868d",x"3afb",x"39b7",x"359e",x"3c71",x"3710",x"b80b",x"bae7",x"868d",x"3b06",x"39bd"),
(x"3501",x"3c9e",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"351b",x"3c9c",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"3501",x"3c9e",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53"),
(x"38c9",x"3c75",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38d4",x"3c73",x"36da",x"38a8",x"3a80",x"8000",x"3a8a",x"3a3e",x"38c9",x"3c75",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43"),
(x"386c",x"3ca2",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"386d",x"3ca8",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"386c",x"3ca2",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05"),
(x"358a",x"3c77",x"36da",x"bbad",x"b482",x"868d",x"3afb",x"39b7",x"3587",x"3c7c",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"358a",x"3c77",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7"),
(x"34e9",x"3c9d",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"3501",x"3c9e",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"34e9",x"3c9d",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57"),
(x"38d4",x"3c73",x"36da",x"38a8",x"3a80",x"8000",x"3a8a",x"3a3e",x"38d9",x"3c71",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d4",x"3c73",x"3710",x"37f2",x"3af1",x"8000",x"3a95",x"3a3e"),
(x"3872",x"3c9f",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"386c",x"3ca2",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"3872",x"3c9f",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08"),
(x"3587",x"3c7c",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"3593",x"3c81",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3587",x"3c7c",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3"),
(x"34cb",x"3c98",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34e9",x"3c9d",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"34cb",x"3c98",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e"),
(x"38d9",x"3c71",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d8",x"3c6f",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38d9",x"3c71",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c"),
(x"3885",x"3c9a",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"3872",x"3c9f",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"3885",x"3c9a",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10"),
(x"3593",x"3c81",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3592",x"3c83",x"36da",x"ba08",x"b941",x"8000",x"3afb",x"39ae",x"3593",x"3c81",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af"),
(x"34bb",x"3c97",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"34cb",x"3c98",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34bb",x"3c97",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61"),
(x"38d8",x"3c6f",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38c7",x"3c6c",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38d8",x"3c6f",x"3710",x"3be4",x"b12f",x"0000",x"3a95",x"3a3b"),
(x"388c",x"3c98",x"36da",x"bb54",x"b669",x"0000",x"3a7d",x"3b13",x"3885",x"3c9a",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"388c",x"3c98",x"3710",x"bbfd",x"a9ab",x"0000",x"3a87",x"3b13"),
(x"3592",x"3c83",x"36da",x"ba08",x"b941",x"8000",x"3a6e",x"3bb2",x"357d",x"3c83",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"3592",x"3c83",x"3710",x"bba4",x"b4bb",x"0000",x"3a79",x"3bb2"),
(x"349b",x"3c96",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"34bb",x"3c97",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"349b",x"3c96",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67"),
(x"38c7",x"3c6c",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38b7",x"3c68",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"38c7",x"3c6c",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34"),
(x"388c",x"3c96",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"388c",x"3c98",x"36da",x"bb54",x"b669",x"0000",x"3a97",x"39c6",x"388c",x"3c96",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8"),
(x"357d",x"3c83",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"3555",x"3c82",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"357d",x"3c83",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae"),
(x"3485",x"3c94",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"349b",x"3c96",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"3485",x"3c94",x"3710",x"b92c",x"3a1a",x"868d",x"3a79",x"3b6c"),
(x"38b7",x"3c68",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"3894",x"3c67",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"38b7",x"3c68",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d"),
(x"3885",x"3c95",x"36da",x"b304",x"3bce",x"0000",x"3a97",x"39ca",x"388c",x"3c96",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"3885",x"3c95",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca"),
(x"3555",x"3c82",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"353f",x"3c7f",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"3555",x"3c82",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6"),
(x"3475",x"3c8f",x"36da",x"baeb",x"3803",x"8000",x"3a6e",x"3b70",x"3485",x"3c94",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"3475",x"3c8f",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70"),
(x"3894",x"3c67",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"3877",x"3c6a",x"36da",x"b8aa",x"ba7f",x"8000",x"3a8a",x"3a15",x"3894",x"3c67",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20"),
(x"3753",x"3cad",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3760",x"3ca9",x"36da",x"3bfa",x"2cac",x"068d",x"3a97",x"3a28",x"3753",x"3cad",x"3710",x"37e4",x"3af5",x"868d",x"3aa1",x"3a2b"),
(x"3a2f",x"3c96",x"36da",x"3bfe",x"a8f0",x"0000",x"3be9",x"39cf",x"3a2d",x"3c81",x"36da",x"3bfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"3a2f",x"3c96",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"353f",x"3c7f",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"351b",x"3c7a",x"36da",x"350e",x"bb96",x"0000",x"3a6e",x"3b9a",x"353f",x"3c7f",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2"),
(x"39f5",x"3cae",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"3a27",x"3cae",x"36da",x"a3ae",x"3bff",x"0000",x"3be3",x"3a63",x"39f5",x"3cae",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f"),
(x"3877",x"3c6a",x"36da",x"b8aa",x"ba7f",x"8000",x"3a8a",x"3a15",x"386d",x"3c6f",x"36da",x"bba8",x"b4a3",x"068d",x"3a8a",x"3a10",x"3877",x"3c6a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15"),
(x"382a",x"3c96",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"3885",x"3c95",x"36da",x"b304",x"3bce",x"0000",x"3a97",x"39ca",x"382a",x"3c96",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed"),
(x"351b",x"3c7a",x"36da",x"350e",x"bb96",x"0000",x"3a6e",x"3b9a",x"3501",x"3c78",x"36da",x"ada8",x"bbf8",x"0000",x"3a6e",x"3b94",x"351b",x"3c7a",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a"),
(x"386d",x"3c6f",x"36da",x"bba8",x"b4a3",x"068d",x"3a8a",x"3a10",x"386c",x"3c74",x"36da",x"bb38",x"36e2",x"068d",x"3a8a",x"3a0c",x"386d",x"3c6f",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10"),
(x"3813",x"3c97",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"382a",x"3c96",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"3813",x"3c97",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5"),
(x"3a2d",x"3c81",x"36da",x"367a",x"bb50",x"0000",x"3bbd",x"3982",x"3a25",x"3c7f",x"36da",x"367a",x"bb50",x"0000",x"3bc0",x"3984",x"3a2d",x"3c81",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a"),
(x"38b2",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"38b7",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38bd",x"3ca0",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3107"),
(x"3592",x"3c93",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20",x"3593",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"359e",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"358a",x"3c77",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2a0e",x"3593",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27"),
(x"359e",x"3c71",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"3593",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"3972",x"3540",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3972",x"3540",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d",x"3985",x"352f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25"),
(x"362c",x"35ca",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"362c",x"35ca",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19",x"35f7",x"35e8",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25"),
(x"36cb",x"3555",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"36cb",x"3555",x"3710",x"b922",x"3a22",x"868d",x"3a87",x"3b28",x"36c2",x"354d",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a"),
(x"3752",x"35f7",x"36da",x"3bdf",x"31a3",x"8000",x"3a97",x"3a21",x"3752",x"35f7",x"3710",x"3bfd",x"aabe",x"0000",x"3aa1",x"3a21",x"3754",x"3600",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23"),
(x"3985",x"352f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3985",x"352f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25",x"3994",x"351b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b"),
(x"36f7",x"35c6",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"36f7",x"35c6",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3",x"363b",x"35c5",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16"),
(x"36c2",x"354d",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36c2",x"354d",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a",x"36c4",x"3540",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c"),
(x"393f",x"362a",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"393f",x"362a",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01",x"392f",x"361d",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa"),
(x"3994",x"351b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3994",x"351b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b",x"3999",x"3519",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d"),
(x"363b",x"35c5",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"363b",x"35c5",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16",x"362c",x"35ca",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19"),
(x"36c4",x"3540",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36c4",x"3540",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c",x"36dc",x"3527",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33"),
(x"3953",x"3620",x"36da",x"39a8",x"39a7",x"068d",x"3be3",x"3a09",x"3953",x"3620",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09",x"393f",x"362a",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01"),
(x"3475",x"35af",x"36da",x"baeb",x"3803",x"068d",x"3a6e",x"3b70",x"3475",x"35af",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70",x"3475",x"358c",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77"),
(x"3710",x"35ca",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"3710",x"35ca",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee",x"36f7",x"35c6",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3"),
(x"36dc",x"3527",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36dc",x"3527",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33",x"36df",x"351a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35"),
(x"395a",x"360e",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"395a",x"360e",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e",x"3953",x"3620",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09"),
(x"3716",x"35cf",x"36da",x"bbb8",x"b42d",x"0000",x"3a54",x"39ec",x"3716",x"35cf",x"3710",x"bbad",x"3480",x"0000",x"3a5f",x"39ec",x"3710",x"35ca",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee"),
(x"36df",x"351a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36df",x"351a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35",x"36e3",x"350c",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38"),
(x"395d",x"3602",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"395d",x"3602",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11",x"395a",x"360e",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e"),
(x"3713",x"35d4",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3713",x"35d4",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60",x"3716",x"35cf",x"3710",x"bbad",x"3480",x"0000",x"3aa1",x"3a61"),
(x"36e3",x"350c",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36e3",x"350c",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38",x"36f7",x"3503",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c"),
(x"3963",x"35fa",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"3963",x"35fa",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14",x"395d",x"3602",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11"),
(x"3705",x"35db",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"3705",x"35db",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d",x"3713",x"35d4",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60"),
(x"36f7",x"3503",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"36f7",x"3503",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c",x"3716",x"3507",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42"),
(x"3972",x"35fb",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3972",x"35fb",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a",x"3963",x"35fa",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14"),
(x"36cb",x"35e6",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"36cb",x"35e6",x"3710",x"b86c",x"baa9",x"0000",x"3aa1",x"3a52",x"3705",x"35db",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d"),
(x"3716",x"3507",x"36da",x"32c2",x"bbd1",x"0000",x"3a7c",x"3b42",x"3716",x"3507",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42",x"372e",x"3511",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47"),
(x"3985",x"360c",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3985",x"360c",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22",x"3972",x"35fb",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a"),
(x"36c2",x"35ef",x"36da",x"bbe7",x"b0ec",x"868d",x"3a97",x"3a50",x"36c2",x"35ef",x"3710",x"baff",x"b7c2",x"0000",x"3aa1",x"3a50",x"36cb",x"35e6",x"3710",x"b86c",x"baa9",x"0000",x"3aa1",x"3a52"),
(x"372e",x"3511",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"372e",x"3511",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47",x"3742",x"3511",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b"),
(x"3994",x"3620",x"36da",x"b458",x"3bb2",x"0000",x"3be3",x"3a29",x"3994",x"3620",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29",x"3985",x"360c",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22"),
(x"36c4",x"35fb",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36c4",x"35fb",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d",x"36c2",x"35ef",x"3710",x"baff",x"b7c2",x"0000",x"3aa1",x"3a50"),
(x"3742",x"3511",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"3742",x"3511",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b",x"3753",x"3518",x"3710",x"38fe",x"ba3f",x"868d",x"3a87",x"3b4e"),
(x"3999",x"3622",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"3999",x"3622",x"3710",x"b328",x"3bcb",x"0000",x"3bd9",x"3a2b",x"3994",x"3620",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29"),
(x"36dc",x"3615",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36dc",x"3615",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47",x"36c4",x"35fb",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d"),
(x"3752",x"3544",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"3752",x"3544",x"3710",x"3be0",x"b1a3",x"0000",x"3a87",x"3b59",x"376c",x"355c",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f"),
(x"39f5",x"3627",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"39f5",x"3627",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f",x"3999",x"3622",x"3710",x"b328",x"3bcb",x"0000",x"3bd9",x"3a2b"),
(x"3a26",x"35cd",x"36da",x"3bff",x"a4d0",x"0000",x"3a18",x"33f3",x"3a26",x"35cd",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4",x"3a27",x"3629",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9"),
(x"36df",x"3621",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36df",x"3621",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44",x"36dc",x"3615",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47"),
(x"376c",x"355c",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"376c",x"355c",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f",x"378c",x"3568",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66"),
(x"36e3",x"362f",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36e3",x"362f",x"3710",x"bb17",x"3766",x"0000",x"3aa1",x"3a41",x"36df",x"3621",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44"),
(x"378c",x"3568",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"378c",x"3568",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66",x"37a8",x"3578",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c"),
(x"36f7",x"3638",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"36f7",x"3638",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d",x"36e3",x"362f",x"3710",x"bb17",x"3766",x"0000",x"3aa1",x"3a41"),
(x"37a8",x"3578",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"37a8",x"3578",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c",x"37b8",x"357b",x"3710",x"2df3",x"bbf7",x"0000",x"3a87",x"3b6f"),
(x"3716",x"3634",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"3716",x"3634",x"3710",x"32c1",x"3bd1",x"0000",x"3aa1",x"3a37",x"36f7",x"3638",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d"),
(x"37b8",x"357b",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"37b8",x"357b",x"3710",x"2df3",x"bbf7",x"0000",x"3a87",x"3b6f",x"380a",x"356e",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81"),
(x"372e",x"362a",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"372e",x"362a",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32",x"3716",x"3634",x"3710",x"32c1",x"3bd1",x"0000",x"3aa1",x"3a37"),
(x"3760",x"3526",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"3760",x"3526",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52",x"375f",x"3530",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54"),
(x"3742",x"362a",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"3742",x"362a",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f",x"372e",x"362a",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32"),
(x"380a",x"356e",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"380a",x"356e",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81",x"3813",x"356c",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84"),
(x"3753",x"3623",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3753",x"3623",x"3710",x"37e4",x"3af5",x"8000",x"3aa1",x"3a2b",x"3742",x"362a",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f"),
(x"3813",x"356c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"3813",x"356c",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84",x"382a",x"3574",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d"),
(x"3999",x"3519",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"3999",x"3519",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d",x"39fc",x"3513",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53"),
(x"376c",x"35e0",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"376c",x"35e0",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a",x"3752",x"35f7",x"3710",x"3bfd",x"aabe",x"0000",x"3aa1",x"3a21"),
(x"382a",x"3574",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"382a",x"3574",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d",x"3885",x"3575",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf"),
(x"378c",x"35d3",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"378c",x"35d3",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14",x"376c",x"35e0",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a"),
(x"3753",x"3518",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3753",x"3518",x"3710",x"38fe",x"ba3f",x"868d",x"3a87",x"3b4e",x"3760",x"3526",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52"),
(x"3475",x"358c",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3475",x"358c",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77",x"3485",x"357a",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b"),
(x"3a2f",x"35c9",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"385a",x"3a2f",x"35c9",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"3861",x"3a26",x"35cd",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"37a8",x"35c3",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"37a8",x"35c3",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e",x"378c",x"35d3",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14"),
(x"3885",x"3575",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"3885",x"3575",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf",x"388c",x"3572",x"3710",x"bb52",x"b671",x"0000",x"3a87",x"3bb2"),
(x"3485",x"357a",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"3485",x"357a",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b",x"349b",x"3571",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80"),
(x"37b8",x"35c0",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"37b8",x"35c0",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b",x"37a8",x"35c3",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e"),
(x"388c",x"3572",x"36da",x"b967",x"b9e6",x"0000",x"3a8a",x"39fb",x"388c",x"3572",x"3710",x"bb52",x"b671",x"0000",x"3a95",x"39fb",x"388c",x"356a",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd"),
(x"349b",x"3571",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"349b",x"3571",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80",x"34bb",x"356f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86"),
(x"380a",x"35cd",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"380a",x"35cd",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9",x"37b8",x"35c0",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b"),
(x"388c",x"356a",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"388c",x"356a",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd",x"3885",x"3562",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00"),
(x"34bb",x"356f",x"36da",x"b140",x"bbe4",x"0000",x"3a6e",x"3b86",x"34bb",x"356f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86",x"34cb",x"356b",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89"),
(x"375f",x"360b",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"375f",x"360b",x"3710",x"3bc1",x"b3d8",x"0000",x"3aa1",x"3a26",x"3760",x"3615",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28"),
(x"3885",x"3562",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"3885",x"3562",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00",x"3872",x"3550",x"3710",x"b9d1",x"397d",x"068d",x"3a95",x"3a08"),
(x"39fc",x"3513",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"39fc",x"3513",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53",x"3a26",x"3514",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63"),
(x"34cb",x"356b",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34cb",x"356b",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89",x"34e9",x"3558",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90"),
(x"3813",x"35cf",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"3813",x"35cf",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5",x"380a",x"35cd",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9"),
(x"3872",x"3550",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"3872",x"3550",x"3710",x"b9d1",x"397d",x"068d",x"3a95",x"3a08",x"386c",x"3541",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c"),
(x"34e9",x"3558",x"36da",x"b698",x"bb49",x"0000",x"3a6e",x"3b90",x"34e9",x"3558",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90",x"3501",x"3552",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94"),
(x"3a26",x"3514",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63",x"39fc",x"3513",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53",x"3a02",x"3513",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55"),
(x"3a20",x"3513",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a02",x"3513",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55",x"3a07",x"3513",x"373c",x"0cea",x"bbfe",x"27bb",x"3a8e",x"3a57"),
(x"3a19",x"3514",x"3749",x"208e",x"bc00",x"128d",x"3a90",x"3a5e",x"3a07",x"3513",x"373c",x"0cea",x"bbfe",x"27bb",x"3a8e",x"3a57",x"3a0d",x"3514",x"374b",x"1481",x"bbff",x"26a1",x"3a91",x"3a59"),
(x"39fc",x"3627",x"3718",x"135f",x"3bfd",x"29a1",x"3bd8",x"3a52",x"39f5",x"3627",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f",x"3a27",x"3629",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63"),
(x"3a00",x"3627",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"39fc",x"3627",x"3718",x"135f",x"3bfd",x"29a1",x"3bd8",x"3a52",x"3a24",x"3629",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62"),
(x"3a07",x"3628",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a00",x"3627",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"3a21",x"3629",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60"),
(x"3a0d",x"3627",x"374b",x"a412",x"3bfd",x"2966",x"3bce",x"3a59",x"3a07",x"3628",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a1a",x"3628",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e"),
(x"3999",x"3519",x"3710",x"975f",x"9f93",x"3c00",x"39f3",x"328d",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e",x"39fc",x"3513",x"3710",x"ba72",x"9a8d",x"38bc",x"39f2",x"333e"),
(x"39f5",x"3627",x"3710",x"b60a",x"25b5",x"3b67",x"3a2d",x"3331",x"39fc",x"3627",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340",x"39fb",x"35cc",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d"),
(x"3999",x"3622",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39fb",x"35cc",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3999",x"3622",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"3999",x"3519",x"3710",x"975f",x"9f93",x"3c00",x"39f3",x"328d",x"3994",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3985",x"360c",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3994",x"3620",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3284",x"3994",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3985",x"360c",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3985",x"352f",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"3269",x"3972",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248"),
(x"3972",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3972",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248",x"3963",x"3541",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"395d",x"3602",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"3963",x"35fa",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"322d",x"3963",x"3541",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"395d",x"3602",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"395d",x"3539",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"3222",x"395a",x"352d",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d"),
(x"395a",x"360e",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"395a",x"352d",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d",x"3953",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211"),
(x"3953",x"3620",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"3953",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211",x"393f",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"393f",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"393f",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed",x"392f",x"351e",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"3915",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"392f",x"361d",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"31d0",x"392f",x"351e",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"3915",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"3915",x"3554",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"31a2",x"38f6",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b"),
(x"38f6",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"38f6",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b",x"38d5",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130"),
(x"38b7",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38b2",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"388c",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"38b2",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"38b7",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"388c",x"356a",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae"),
(x"388c",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae",x"38b2",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"38b0",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"388c",x"356a",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"388c",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"38b0",x"355b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"38c7",x"351f",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38b7",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38c9",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a"),
(x"38c7",x"361c",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38d4",x"35ff",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d",x"38c9",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a"),
(x"38d8",x"360d",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3135",x"38d9",x"3608",x"3710",x"0000",x"0000",x"3c00",x"3a26",x"3136",x"38d4",x"35ff",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d"),
(x"38d8",x"352e",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3135",x"38c7",x"351f",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38d4",x"353c",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d"),
(x"388c",x"356a",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"38b7",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"3894",x"350e",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"3894",x"362d",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"38b7",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"388c",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"3877",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3894",x"362d",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"3885",x"35da",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"386d",x"3610",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"3076",x"3877",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3872",x"35eb",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080"),
(x"3885",x"3562",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"3894",x"350e",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc",x"3877",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088"),
(x"3872",x"3550",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"3877",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088",x"386d",x"352c",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3076"),
(x"38b0",x"355b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"388c",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"388c",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"38b2",x"3565",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b0",x"355b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"38b0",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38bf",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38b2",x"3565",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b2",x"35d6",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"38bf",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38bf",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"3109",x"38d5",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130"),
(x"388c",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"388c",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"30ad",x"3885",x"3575",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"382a",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3885",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30a2",x"3885",x"3575",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"382a",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"382a",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2ffc",x"3813",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"3813",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"3813",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac",x"380a",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"3752",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"3752",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30",x"3716",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"3710",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb",x"3710",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2dbb",x"3716",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"3713",x"3567",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"3716",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5",x"3752",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"3713",x"35d4",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3754",x"3600",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33",x"3752",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"372e",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"36dc",x"3527",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"3713",x"3567",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"3713",x"35d4",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"36dc",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e",x"372e",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"3705",x"35db",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36c4",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33",x"36dc",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"3705",x"3560",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"3713",x"3567",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"36dc",x"3527",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"36cb",x"3555",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"2d40",x"3705",x"3560",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"36c4",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"36cb",x"35e6",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2d40",x"36c2",x"35ef",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2d2f",x"36c4",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"3742",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"375f",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47",x"3754",x"3600",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"3753",x"3623",x"3710",x"0000",x"0000",x"3c00",x"3a2c",x"2e32",x"3760",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2e49",x"375f",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"3742",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"372e",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3754",x"353b",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"3753",x"3518",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2e32",x"3742",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"375f",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"36dc",x"3527",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"372e",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3716",x"3507",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"36df",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"3716",x"3507",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4",x"36f7",x"3503",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"3716",x"3634",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"372e",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0",x"36dc",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"36f7",x"3638",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e",x"3716",x"3634",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"36df",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"376c",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e",x"376c",x"355c",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2e5e",x"3752",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"378c",x"3568",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"376c",x"355c",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2e5e",x"376c",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"37a8",x"3578",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9",x"378c",x"3568",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"378c",x"35d3",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"37b8",x"35c0",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7",x"37b8",x"357b",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2ee7",x"37a8",x"3578",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"380a",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b",x"37b8",x"357b",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2ee7",x"37b8",x"35c0",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"36f7",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d",x"3710",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2dbb",x"3710",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"3587",x"35d9",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"29f9",x"358a",x"35ee",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"2a04",x"3593",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"35bd",x"3610",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35f1",x"35f1",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"35bd",x"352b",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"359e",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"35d3",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35bd",x"352b",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"35f1",x"354a",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"35e4",x"352a",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35d3",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35f3",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"35f5",x"3528",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b84",x"35e4",x"352a",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35fd",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"35d3",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35f3",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d",x"35f1",x"35f1",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"35e4",x"3612",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35fd",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0",x"35f3",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"35f5",x"3613",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b84",x"35fd",x"360e",x"3710",x"868d",x"0000",x"3c00",x"3a27",x"2ba0",x"35fd",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"3592",x"357c",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20",x"3592",x"35bf",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"362c",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"363b",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"362c",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"362c",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"363b",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"363b",x"35c5",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2c3f",x"36f7",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"357d",x"35bd",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"3592",x"35bf",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20",x"3592",x"357c",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"3555",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"357d",x"35bd",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"357d",x"357e",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"353f",x"35cd",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"3555",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"3555",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949"),
(x"351b",x"35e2",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"353f",x"35cd",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"353f",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"3501",x"35e9",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a",x"351b",x"35e2",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"351b",x"3559",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878"),
(x"34e9",x"3558",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b",x"34e9",x"35e3",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"278b",x"3501",x"35e9",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"34cb",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3",x"34e9",x"35e3",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"278b",x"34e9",x"3558",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b"),
(x"34bb",x"356f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643",x"34bb",x"35cc",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2643",x"34cb",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"349b",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"34bb",x"35cc",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2643",x"34bb",x"356f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643"),
(x"3485",x"35c1",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"349b",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"349b",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f"),
(x"3475",x"35af",x"3710",x"0000",x"0000",x"3c00",x"3a13",x"2451",x"3485",x"35c1",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"3485",x"357a",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"3a01",x"35ce",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"39fb",x"35cc",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"39fc",x"3627",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340"),
(x"3a09",x"35cf",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a01",x"35ce",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"3a00",x"3627",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c"),
(x"3a09",x"35cf",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a07",x"3628",x"373c",x"baa1",x"a6bb",x"3879",x"3a2d",x"3366",x"3a0d",x"3627",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378"),
(x"3a0f",x"35cf",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a0d",x"3627",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378",x"3a14",x"3628",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385"),
(x"3a15",x"35ce",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a14",x"3628",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385",x"3a1a",x"3628",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a20",x"35ce",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a1a",x"35ce",x"3746",x"38a5",x"a839",x"3a81",x"3a1a",x"338e",x"3a1a",x"3628",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a24",x"3629",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a20",x"35ce",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a21",x"3629",x"373a",x"3acd",x"a5ae",x"3834",x"3a2d",x"33a3"),
(x"3a24",x"3629",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a27",x"3629",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9",x"3a26",x"35cd",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4"),
(x"3a02",x"35c9",x"3711",x"315a",x"2baa",x"3bdf",x"3a19",x"3349",x"3a03",x"3574",x"370e",x"34eb",x"a6e9",x"3b9c",x"3a06",x"334b",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3a02",x"35c9",x"3711",x"b40d",x"bb3a",x"3584",x"3b18",x"387b",x"39fb",x"35cc",x"3713",x"aedc",x"bb7b",x"3565",x"3b16",x"387a",x"3a01",x"35ce",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879"),
(x"3a02",x"35c9",x"3711",x"b40d",x"bb3a",x"3584",x"3b18",x"387b",x"3a01",x"35ce",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879",x"3a04",x"35c9",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879"),
(x"3a04",x"35c9",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879",x"3a01",x"35ce",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3879",x"3a09",x"35cf",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875"),
(x"3a08",x"35c8",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a09",x"35cf",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875",x"3a0f",x"35cf",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873"),
(x"3a0f",x"35c8",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a0f",x"35cf",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873",x"3a15",x"35ce",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"3871"),
(x"3a17",x"35c8",x"3751",x"2fd8",x"39a6",x"3994",x"3b24",x"3871",x"3a15",x"35ce",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"3871",x"3a1d",x"35c8",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e"),
(x"3a1d",x"35c8",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e",x"3a15",x"35ce",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"3871",x"3a1a",x"35ce",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e"),
(x"3a24",x"35c8",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a1a",x"35ce",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e",x"3a20",x"35ce",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b"),
(x"3a2a",x"35c8",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a20",x"35ce",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b",x"3a26",x"35cd",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3a25",x"3577",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a1f",x"356e",x"3733",x"3800",x"ba99",x"3437",x"3bb7",x"3993",x"3a21",x"3577",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a18",x"356e",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998",x"3a19",x"3577",x"374d",x"3243",x"b807",x"3abb",x"3bb5",x"3999",x"3a21",x"3577",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a11",x"3577",x"374a",x"b548",x"b37e",x"3b50",x"3bb7",x"399b",x"3a19",x"3577",x"374d",x"3243",x"b807",x"3abb",x"3bb5",x"3999",x"3a18",x"356e",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998"),
(x"3a0d",x"3514",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b",x"3a07",x"3513",x"373c",x"bac4",x"2853",x"3841",x"39f2",x"336a",x"3a09",x"356e",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369"),
(x"3a25",x"3577",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a2d",x"3576",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a",x"3a25",x"356e",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c"),
(x"3a2d",x"3576",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a2a",x"35c8",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a2f",x"35c9",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"3a2a",x"35c8",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a2d",x"3576",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a25",x"3577",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3"),
(x"3a24",x"35c8",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a25",x"3577",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3",x"3a21",x"3577",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6"),
(x"3a1d",x"35c8",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a21",x"3577",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6",x"3a19",x"3577",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a0f",x"35c8",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a17",x"35c8",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3be8",x"39eb",x"3a19",x"3577",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a08",x"35c8",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a0f",x"35c8",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a11",x"3577",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed"),
(x"3a02",x"35c9",x"3711",x"bbe1",x"a6cf",x"3179",x"3be9",x"39fb",x"3a04",x"35c9",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7",x"3a03",x"3574",x"370e",x"bbc2",x"ab4f",x"338c",x"3bf9",x"39fa"),
(x"39fc",x"3513",x"3710",x"ba72",x"9a8d",x"38bc",x"39f2",x"333e",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e",x"3a02",x"3513",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352"),
(x"3a09",x"3575",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a11",x"3577",x"374a",x"b548",x"b37e",x"3b50",x"3bb7",x"399b",x"3a10",x"356e",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b"),
(x"3a09",x"356e",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"39fc",x"3571",x"3713",x"af5f",x"3bdb",x"30c1",x"3bc0",x"39a6",x"3a03",x"3574",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bbd",x"39a7"),
(x"3a10",x"356e",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a14",x"3513",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387",x"3a0d",x"3514",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b"),
(x"3a18",x"356e",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a19",x"3514",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392",x"3a14",x"3513",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387"),
(x"3a1f",x"356e",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a20",x"3513",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa",x"3a19",x"3514",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392"),
(x"3a25",x"356e",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0",x"3a26",x"3514",x"3710",x"3bcf",x"2680",x"32dc",x"39f4",x"33ca",x"3a20",x"3513",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa"),
(x"392f",x"361d",x"36da",x"b73b",x"3b22",x"8000",x"3be3",x"39fa",x"392f",x"361d",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa",x"3915",x"35e8",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec"),
(x"3705",x"3560",x"36da",x"b675",x"3b51",x"0000",x"3a7c",x"3b1d",x"3705",x"3560",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d",x"36cb",x"3555",x"3710",x"b922",x"3a22",x"868d",x"3a87",x"3b28"),
(x"35f7",x"35e8",x"36da",x"3a05",x"3943",x"8000",x"3a54",x"3a25",x"35f7",x"35e8",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25",x"35f1",x"35f1",x"3710",x"3bf9",x"ad21",x"0000",x"3a5f",x"3a27"),
(x"3963",x"3541",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"3963",x"3541",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17",x"3972",x"3540",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d"),
(x"3754",x"3600",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"3754",x"3600",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23",x"375f",x"360b",x"3710",x"3bc1",x"b3d8",x"0000",x"3aa1",x"3a26"),
(x"3713",x"3567",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3713",x"3567",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a",x"3705",x"3560",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d"),
(x"35f1",x"35f1",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f1",x"35f1",x"3710",x"3bf9",x"ad21",x"0000",x"3a5f",x"3a27",x"35f3",x"35f7",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28"),
(x"395d",x"3539",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"395d",x"3539",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14",x"3963",x"3541",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17"),
(x"3915",x"35e8",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"3915",x"35e8",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec",x"38f6",x"35ca",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de"),
(x"3716",x"356c",x"36da",x"bbad",x"b480",x"0000",x"3a7c",x"3b19",x"3716",x"356c",x"3710",x"bbb8",x"342e",x"0000",x"3a87",x"3b19",x"3713",x"3567",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a"),
(x"35f3",x"35f7",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35f3",x"35f7",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28",x"35fd",x"3605",x"3710",x"3bf0",x"aff4",x"068d",x"3a5f",x"3a2b"),
(x"395a",x"352d",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"395a",x"352d",x"3710",x"3b46",x"b6a7",x"868d",x"3a85",x"3a12",x"395d",x"3539",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14"),
(x"38f6",x"35ca",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"38f6",x"35ca",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de",x"38d5",x"35c2",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1"),
(x"3710",x"3571",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"3710",x"3571",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f",x"3716",x"356c",x"3710",x"bbb8",x"342e",x"0000",x"3b06",x"3a11"),
(x"35fd",x"3605",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35fd",x"3605",x"3710",x"3bf0",x"aff4",x"068d",x"3a5f",x"3a2b",x"35fd",x"360e",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d"),
(x"3953",x"351b",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"3953",x"351b",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d",x"395a",x"352d",x"3710",x"3b46",x"b6a7",x"868d",x"3a85",x"3a12"),
(x"38d5",x"35c2",x"36da",x"1953",x"3c00",x"0000",x"3be3",x"39d1",x"38d5",x"35c2",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1",x"38bf",x"35c9",x"3710",x"35f3",x"3b6d",x"0000",x"3bd9",x"39c8"),
(x"36f7",x"3576",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"36f7",x"3576",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a",x"3710",x"3571",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f"),
(x"35fd",x"360e",x"36da",x"3b87",x"3567",x"068d",x"3a54",x"3a2d",x"35fd",x"360e",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d",x"35f5",x"3613",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e"),
(x"393f",x"3511",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"393f",x"3511",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05",x"3953",x"351b",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d"),
(x"38bf",x"35c9",x"36da",x"3489",x"3bac",x"0000",x"3be3",x"39c8",x"38bf",x"35c9",x"3710",x"35f3",x"3b6d",x"0000",x"3bd9",x"39c8",x"38b2",x"35d6",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2"),
(x"362c",x"3571",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"362c",x"3571",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4",x"363b",x"3576",x"3710",x"3439",x"bbb7",x"868d",x"3b06",x"39e7"),
(x"35f5",x"3613",x"36da",x"364b",x"3b5a",x"868d",x"3a54",x"3a2e",x"35f5",x"3613",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e",x"35e4",x"3612",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32"),
(x"392f",x"351e",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"392f",x"351e",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff",x"393f",x"3511",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05"),
(x"38b2",x"35d6",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38b2",x"35d6",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2",x"38b0",x"35e0",x"3710",x"3ba6",x"b4ab",x"0000",x"3bd9",x"39c0"),
(x"363b",x"3576",x"36da",x"34be",x"bba4",x"0000",x"3afb",x"39e7",x"363b",x"3576",x"3710",x"3439",x"bbb7",x"868d",x"3b06",x"39e7",x"36f7",x"3576",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a"),
(x"35e4",x"3612",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35e4",x"3612",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32",x"35d3",x"360b",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35"),
(x"3754",x"353b",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"3754",x"353b",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57",x"3752",x"3544",x"3710",x"3be0",x"b1a3",x"0000",x"3a87",x"3b59"),
(x"38b0",x"35e0",x"36da",x"3bfc",x"2b2b",x"0000",x"3be3",x"39c0",x"38b0",x"35e0",x"3710",x"3ba6",x"b4ab",x"0000",x"3bd9",x"39c0",x"38b2",x"35e8",x"3710",x"399c",x"b9b3",x"8000",x"3bd9",x"39be"),
(x"35f7",x"3553",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"35f7",x"3553",x"3710",x"3a05",x"b943",x"0000",x"3b06",x"39d8",x"362c",x"3571",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4"),
(x"35d3",x"360b",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35d3",x"360b",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35",x"35bd",x"3610",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39"),
(x"3915",x"3554",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"3915",x"3554",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1",x"392f",x"351e",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff"),
(x"38b2",x"35e8",x"36da",x"3a58",x"b8de",x"0000",x"3a7d",x"3ac5",x"38b2",x"35e8",x"3710",x"399c",x"b9b3",x"8000",x"3a87",x"3ac5",x"38bd",x"35f3",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9"),
(x"35f1",x"354a",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f1",x"354a",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6",x"35f7",x"3553",x"3710",x"3a05",x"b943",x"0000",x"3b06",x"39d8"),
(x"35bd",x"3610",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"35bd",x"3610",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39",x"359e",x"3605",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40"),
(x"375f",x"3530",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"375f",x"3530",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54",x"3754",x"353b",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57"),
(x"38bd",x"35f3",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38bd",x"35f3",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9",x"38c9",x"35f7",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace"),
(x"35f3",x"3544",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35f3",x"3544",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5",x"35f1",x"354a",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6"),
(x"359e",x"3605",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"359e",x"3605",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40",x"358a",x"35ee",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45"),
(x"38f6",x"3572",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"38f6",x"3572",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4",x"3915",x"3554",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1"),
(x"38c9",x"35f7",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38c9",x"35f7",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace",x"38d4",x"35ff",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2"),
(x"35fd",x"3536",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35fd",x"3536",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2",x"35f3",x"3544",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5"),
(x"358a",x"35ee",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"358a",x"35ee",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45",x"3587",x"35d9",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49"),
(x"38d5",x"3579",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38d5",x"3579",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7",x"38f6",x"3572",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4"),
(x"38d4",x"35ff",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38d4",x"35ff",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2",x"38d9",x"3608",x"3710",x"3bfc",x"ab00",x"868d",x"3a87",x"3ad5"),
(x"3a26",x"3514",x"36da",x"3bff",x"26b5",x"0000",x"39f5",x"33fa",x"3a26",x"3514",x"3710",x"3bcf",x"2680",x"32dc",x"39f4",x"33ca",x"3a25",x"356e",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0"),
(x"35fd",x"352d",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35fd",x"352d",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0",x"35fd",x"3536",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2"),
(x"3587",x"35d9",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"3587",x"35d9",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49",x"3593",x"35c7",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d"),
(x"38bf",x"3572",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38bf",x"3572",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf",x"38d5",x"3579",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7"),
(x"38d9",x"3608",x"36da",x"3b87",x"b565",x"0000",x"3a7d",x"3ad5",x"38d9",x"3608",x"3710",x"3bfc",x"ab00",x"868d",x"3a87",x"3ad5",x"38d8",x"360d",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6"),
(x"35f5",x"3528",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35f5",x"3528",x"3710",x"364b",x"bb5a",x"068d",x"3b06",x"39ce",x"35fd",x"352d",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0"),
(x"3593",x"35c7",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3593",x"35c7",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d",x"3592",x"35bf",x"3710",x"ba08",x"3941",x"0000",x"3a5f",x"3a4f"),
(x"38b2",x"3565",x"36da",x"3af2",x"b7f0",x"0000",x"3a7b",x"39c9",x"38b2",x"3565",x"3710",x"3a0a",x"b93e",x"8000",x"3a85",x"39c9",x"38bf",x"3572",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf"),
(x"38d8",x"360d",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38d8",x"360d",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6",x"38c7",x"361c",x"3710",x"364a",x"3b5b",x"0000",x"3a87",x"3add"),
(x"35e4",x"352a",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35e4",x"352a",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb",x"35f5",x"3528",x"3710",x"364b",x"bb5a",x"068d",x"3b06",x"39ce"),
(x"3592",x"35bf",x"36da",x"bba4",x"34bb",x"0000",x"3a6e",x"3b35",x"3592",x"35bf",x"3710",x"ba08",x"3941",x"0000",x"3a79",x"3b35",x"357d",x"35bd",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39"),
(x"38b0",x"355b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b0",x"355b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d",x"38b2",x"3565",x"3710",x"3a0a",x"b93e",x"8000",x"3a95",x"3a50"),
(x"38c7",x"361c",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38c7",x"361c",x"3710",x"364a",x"3b5b",x"0000",x"3a87",x"3add",x"38b7",x"362a",x"3710",x"32f7",x"3bce",x"8000",x"3a87",x"3ae4"),
(x"35d3",x"3530",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35d3",x"3530",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8",x"35e4",x"352a",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb"),
(x"357d",x"35bd",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"357d",x"35bd",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39",x"3555",x"35c2",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41"),
(x"38b2",x"3553",x"36da",x"399c",x"39b3",x"8000",x"3a8a",x"3a4c",x"38b2",x"3553",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c",x"38b0",x"355b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d"),
(x"38b7",x"362a",x"36da",x"3528",x"3b92",x"068d",x"3a7d",x"3ae4",x"38b7",x"362a",x"3710",x"32f7",x"3bce",x"8000",x"3a87",x"3ae4",x"3894",x"362d",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1"),
(x"35bd",x"352b",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"35bd",x"352b",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3",x"35d3",x"3530",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8"),
(x"3555",x"35c2",x"36da",x"345b",x"3bb2",x"0000",x"3a6e",x"3b41",x"3555",x"35c2",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41",x"353f",x"35cd",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46"),
(x"38bd",x"3548",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38bd",x"3548",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47",x"38b2",x"3553",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c"),
(x"3894",x"362d",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"3894",x"362d",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1",x"3877",x"3621",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc"),
(x"359e",x"3536",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"359e",x"3536",x"3710",x"b80b",x"bae7",x"8000",x"3b06",x"39bd",x"35bd",x"352b",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3"),
(x"353f",x"35cd",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"353f",x"35cd",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46",x"351b",x"35e2",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e"),
(x"38c9",x"3544",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38c9",x"3544",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43",x"38bd",x"3548",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47"),
(x"3877",x"3621",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"3877",x"3621",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc",x"386d",x"3610",x"3710",x"bba8",x"34a3",x"0000",x"3a87",x"3b01"),
(x"358a",x"354d",x"36da",x"bbad",x"b481",x"8000",x"3afb",x"39b7",x"358a",x"354d",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7",x"359e",x"3536",x"3710",x"b80b",x"bae7",x"8000",x"3b06",x"39bd"),
(x"351b",x"35e2",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"351b",x"35e2",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e",x"3501",x"35e9",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53"),
(x"38d4",x"353c",x"36da",x"38a8",x"3a80",x"0000",x"3a8a",x"3a3e",x"38d4",x"353c",x"3710",x"37f2",x"3af1",x"0000",x"3a95",x"3a3e",x"38c9",x"3544",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43"),
(x"386d",x"3610",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"386d",x"3610",x"3710",x"bba8",x"34a3",x"0000",x"3a87",x"3b01",x"386c",x"35fa",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05"),
(x"3587",x"3562",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"3587",x"3562",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3",x"358a",x"354d",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7"),
(x"3501",x"35e9",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"3501",x"35e9",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53",x"34e9",x"35e3",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57"),
(x"38d9",x"3533",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d9",x"3533",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c",x"38d4",x"353c",x"3710",x"37f2",x"3af1",x"0000",x"3a95",x"3a3e"),
(x"386c",x"35fa",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"386c",x"35fa",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05",x"3872",x"35eb",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08"),
(x"3593",x"3574",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3593",x"3574",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af",x"3587",x"3562",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3"),
(x"34e9",x"35e3",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"34e9",x"35e3",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57",x"34cb",x"35d1",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e"),
(x"38d8",x"352e",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38d8",x"352e",x"3710",x"3be4",x"b12f",x"8a8d",x"3a95",x"3a3b",x"38d9",x"3533",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c"),
(x"3872",x"35eb",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"3872",x"35eb",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08",x"3885",x"35da",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10"),
(x"3592",x"357c",x"36da",x"ba08",x"b941",x"8000",x"3afb",x"39ae",x"3592",x"357c",x"3710",x"bba4",x"b4bb",x"0000",x"3b06",x"39ae",x"3593",x"3574",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af"),
(x"34cb",x"35d1",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34cb",x"35d1",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e",x"34bb",x"35cc",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61"),
(x"38c7",x"351f",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38c7",x"351f",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34",x"38d8",x"352e",x"3710",x"3be4",x"b12f",x"8a8d",x"3a95",x"3a3b"),
(x"3885",x"35da",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"3885",x"35da",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10",x"388c",x"35d1",x"3710",x"bbfd",x"a9ab",x"0000",x"3a87",x"3b13"),
(x"357d",x"357e",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"357d",x"357e",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae",x"3592",x"357c",x"3710",x"bba4",x"b4bb",x"0000",x"3a79",x"3bb2"),
(x"34bb",x"35cc",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"34bb",x"35cc",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61",x"349b",x"35ca",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67"),
(x"38b7",x"3511",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"38b7",x"3511",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d",x"38c7",x"351f",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34"),
(x"388c",x"35d1",x"36da",x"bb54",x"b669",x"0000",x"3a97",x"39c6",x"388c",x"35d1",x"3710",x"bbfd",x"a9ab",x"0000",x"3aa1",x"39c6",x"388c",x"35c9",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8"),
(x"3555",x"3579",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"3555",x"3579",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6",x"357d",x"357e",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae"),
(x"349b",x"35ca",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"349b",x"35ca",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67",x"3485",x"35c1",x"3710",x"b92c",x"3a1a",x"8000",x"3a79",x"3b6c"),
(x"3894",x"350e",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"3894",x"350e",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20",x"38b7",x"3511",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d"),
(x"388c",x"35c9",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"388c",x"35c9",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8",x"3885",x"35c6",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca"),
(x"353f",x"356e",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"353f",x"356e",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2",x"3555",x"3579",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6"),
(x"3485",x"35c1",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"3485",x"35c1",x"3710",x"b92c",x"3a1a",x"8000",x"3a79",x"3b6c",x"3475",x"35af",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70"),
(x"3877",x"351a",x"36da",x"b8aa",x"ba7f",x"068d",x"3a8a",x"3a15",x"3877",x"351a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15",x"3894",x"350e",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20"),
(x"3760",x"3615",x"36da",x"3bfa",x"2cac",x"8a8d",x"3a97",x"3a28",x"3760",x"3615",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28",x"3753",x"3623",x"3710",x"37e4",x"3af5",x"8000",x"3aa1",x"3a2b"),
(x"3a2d",x"3576",x"36da",x"3bfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"3a2d",x"3576",x"3710",x"3bde",x"a849",x"31a9",x"3bf8",x"39db",x"3a2f",x"35c9",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"351b",x"3559",x"36da",x"350e",x"bb96",x"068d",x"3a6e",x"3b9a",x"351b",x"3559",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a",x"353f",x"356e",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2"),
(x"3a27",x"3629",x"36da",x"a3ae",x"3bff",x"0000",x"3be3",x"3a63",x"3a27",x"3629",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63",x"39f5",x"3627",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f"),
(x"386d",x"352c",x"36da",x"bba8",x"b4a3",x"8000",x"3a8a",x"3a10",x"386d",x"352c",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10",x"3877",x"351a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15"),
(x"3885",x"35c6",x"36da",x"b305",x"3bce",x"0000",x"3a97",x"39ca",x"3885",x"35c6",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca",x"382a",x"35c7",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed"),
(x"3501",x"3552",x"36da",x"ada6",x"bbf8",x"8000",x"3a6e",x"3b94",x"3501",x"3552",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94",x"351b",x"3559",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a"),
(x"386c",x"3541",x"36da",x"bb38",x"36e2",x"8000",x"3a8a",x"3a0c",x"386c",x"3541",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c",x"386d",x"352c",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10"),
(x"382a",x"35c7",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"382a",x"35c7",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed",x"3813",x"35cf",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5"),
(x"3a25",x"356e",x"36da",x"367a",x"bb50",x"0000",x"3bc0",x"3984",x"3a25",x"356e",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c",x"3a2d",x"3576",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a"),
(x"3a1f",x"356e",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a25",x"356e",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0",x"3a20",x"3513",x"3732",x"3b18",x"2439",x"3763",x"39f3",x"33aa"),
(x"3a18",x"356e",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a1f",x"356e",x"3733",x"3b23",x"2518",x"3737",x"3a06",x"339f",x"3a19",x"3514",x"3749",x"3871",x"2587",x"3aa6",x"39f3",x"3392"),
(x"3a10",x"356e",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a18",x"356e",x"3748",x"36c9",x"29dc",x"3b3c",x"3a06",x"3388",x"3a14",x"3513",x"374e",x"2fa2",x"2997",x"3bef",x"39f2",x"3387"),
(x"3a09",x"356e",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a10",x"356e",x"3749",x"b4de",x"2b76",x"3b9b",x"3a06",x"337b",x"3a0d",x"3514",x"374b",x"b745",x"2966",x"3b1e",x"39f2",x"337b"),
(x"3a09",x"3575",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a09",x"356e",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"3a03",x"3574",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bbd",x"39a7"),
(x"3a09",x"356e",x"373b",x"b7a6",x"3a67",x"35ca",x"3bba",x"399e",x"3a09",x"3575",x"373a",x"baf6",x"2b34",x"37d2",x"3bb9",x"399f",x"3a10",x"356e",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b"),
(x"3a08",x"35c8",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a09",x"3575",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1",x"3a04",x"35c9",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7"),
(x"3a03",x"3574",x"370e",x"bbc2",x"ab4f",x"338c",x"3bf9",x"39fa",x"3a04",x"35c9",x"3727",x"bbc5",x"a901",x"3377",x"3be8",x"39f7",x"3a09",x"3575",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1"),
(x"3a09",x"3575",x"373a",x"ba80",x"a874",x"38a7",x"3bf8",x"39f1",x"3a08",x"35c8",x"373e",x"bb1c",x"a938",x"374b",x"3be8",x"39f2",x"3a11",x"3577",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed"),
(x"3a11",x"3577",x"374a",x"b575",x"a7e2",x"3b84",x"3bf7",x"39ed",x"3a0f",x"35c8",x"374d",x"b891",x"aa52",x"3a8d",x"3be8",x"39ee",x"3a19",x"3577",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a17",x"35c8",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3be8",x"39eb",x"3a1d",x"35c8",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a19",x"3577",x"374d",x"3400",x"aa73",x"3bbc",x"3bf7",x"39ea"),
(x"3a1d",x"35c8",x"374d",x"3802",x"a90b",x"3aea",x"3be8",x"39e8",x"3a24",x"35c8",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a21",x"3577",x"3744",x"3962",x"a91e",x"39e8",x"3bf7",x"39e6"),
(x"3a24",x"35c8",x"373f",x"3a93",x"a694",x"388c",x"3be8",x"39e4",x"3a2a",x"35c8",x"3725",x"3b3f",x"a65f",x"36c3",x"3be8",x"39de",x"3a25",x"3577",x"3738",x"3aa3",x"a5dc",x"3875",x"3bf7",x"39e3"),
(x"3a1f",x"356e",x"3733",x"3800",x"ba99",x"3437",x"3bb7",x"3993",x"3a25",x"3577",x"3738",x"36f3",x"bae7",x"3422",x"3bb5",x"3992",x"3a25",x"356e",x"3710",x"3700",x"bb23",x"2f05",x"3bba",x"398c"),
(x"3a02",x"3513",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352",x"3a09",x"356e",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a07",x"3513",x"373c",x"bac4",x"2853",x"3841",x"39f2",x"336a"),
(x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e",x"3a09",x"356e",x"373b",x"b9d7",x"2404",x"3976",x"3a05",x"3369",x"3a02",x"3513",x"3724",x"bb1f",x"1a24",x"3747",x"39f2",x"3352"),
(x"3a10",x"356e",x"3749",x"b3aa",x"a4af",x"3bc3",x"3bb8",x"399b",x"3a11",x"3577",x"374a",x"b548",x"b37e",x"3b50",x"3bb7",x"399b",x"3a18",x"356e",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998"),
(x"3a1f",x"356e",x"3733",x"3800",x"ba99",x"3437",x"3bb7",x"3993",x"3a18",x"356e",x"3748",x"2918",x"b8de",x"3a57",x"3bb7",x"3998",x"3a21",x"3577",x"3744",x"37e0",x"ba17",x"36be",x"3bb4",x"3995"),
(x"3a2f",x"35c9",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"3861",x"3a2a",x"35c8",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a26",x"35cd",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3a2a",x"35c8",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3865",x"3a24",x"35c8",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a20",x"35ce",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"386b"),
(x"3a24",x"35c8",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"386a",x"3a1d",x"35c8",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"386e",x"3a1a",x"35ce",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"386e"),
(x"3a17",x"35c8",x"3751",x"2fd8",x"39a6",x"3994",x"3b24",x"3871",x"3a0f",x"35c8",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a15",x"35ce",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"3871"),
(x"3a0f",x"35c8",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3873",x"3a08",x"35c8",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a0f",x"35cf",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3873"),
(x"3a08",x"35c8",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3876",x"3a04",x"35c9",x"3727",x"bada",x"b46b",x"36f8",x"3b1b",x"3879",x"3a09",x"35cf",x"373e",x"ba28",x"9e0a",x"391a",x"3b1e",x"3875"),
(x"39fb",x"35cc",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d",x"3a02",x"35c9",x"3711",x"315a",x"2baa",x"3bdf",x"3a19",x"3349",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3a20",x"35ce",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a24",x"3629",x"372b",x"3b86",x"a8a8",x"3564",x"3a2d",x"33b1",x"3a26",x"35cd",x"3710",x"3bed",x"a7ae",x"3024",x"3a19",x"33c4"),
(x"3a21",x"3629",x"373a",x"3acd",x"a5ae",x"3834",x"3a2d",x"33a3",x"3a20",x"35ce",x"3739",x"3abd",x"a8b5",x"384c",x"3a1a",x"339e",x"3a1a",x"3628",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a1a",x"35ce",x"3746",x"38a5",x"a839",x"3a81",x"3a1a",x"338e",x"3a15",x"35ce",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a1a",x"3628",x"3749",x"38cd",x"a812",x"3a64",x"3a2d",x"3391"),
(x"3a15",x"35ce",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a1a",x"3385",x"3a0f",x"35cf",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a14",x"3628",x"374f",x"32be",x"a89e",x"3bd0",x"3a2d",x"3385"),
(x"3a0f",x"35cf",x"3749",x"b771",x"a91b",x"3b13",x"3a1a",x"3379",x"3a09",x"35cf",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a0d",x"3627",x"374b",x"b6cb",x"a758",x"3b3d",x"3a2d",x"3378"),
(x"3a07",x"3628",x"373c",x"baa1",x"a6bb",x"3879",x"3a2d",x"3366",x"3a09",x"35cf",x"373e",x"ba21",x"a786",x"3921",x"3a1a",x"336a",x"3a00",x"3627",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c"),
(x"3a00",x"3627",x"3722",x"ba6c",x"a860",x"38c2",x"3a2d",x"334c",x"3a01",x"35ce",x"371c",x"b9f4",x"a495",x"3957",x"3a1a",x"334a",x"39fc",x"3627",x"3718",x"b8fc",x"a86a",x"3a40",x"3a2d",x"3340"),
(x"3475",x"358c",x"3710",x"0000",x"0000",x"3c00",x"3a0c",x"2451",x"3475",x"35af",x"3710",x"0000",x"0000",x"3c00",x"3a13",x"2451",x"3485",x"357a",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"3485",x"357a",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"24c1",x"3485",x"35c1",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"24c1",x"349b",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f"),
(x"349b",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"255f",x"349b",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"255f",x"34bb",x"356f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643"),
(x"34cb",x"356b",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"26b3",x"34bb",x"356f",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2643",x"34cb",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"34cb",x"356b",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"26b3",x"34cb",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"26b3",x"34e9",x"3558",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b"),
(x"3501",x"3552",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"281a",x"34e9",x"3558",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"278b",x"3501",x"35e9",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"3501",x"3552",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"281a",x"3501",x"35e9",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"281a",x"351b",x"3559",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878"),
(x"351b",x"3559",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2878",x"351b",x"35e2",x"3710",x"0000",x"0000",x"3c00",x"3a1e",x"2878",x"353f",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"353f",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"28fb",x"353f",x"35cd",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"28fb",x"3555",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949"),
(x"3555",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2949",x"3555",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2949",x"357d",x"357e",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"357d",x"357e",x"3710",x"0000",x"0000",x"3c00",x"3a09",x"29d7",x"357d",x"35bd",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"29d7",x"3592",x"357c",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"36f7",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2d8d",x"363b",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"36f7",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"363b",x"35c5",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2c3f",x"363b",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2c3f",x"362c",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"362c",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2c23",x"362c",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2c23",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b",x"3592",x"35bf",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"35e4",x"3612",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35f5",x"3613",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b84",x"35fd",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"35d3",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35e4",x"3612",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2b48",x"35f3",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"35bd",x"3610",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35d3",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2b0a",x"35f1",x"35f1",x"3710",x"0000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"35fd",x"352d",x"3710",x"868d",x"0000",x"3c00",x"39f7",x"2ba0",x"35f5",x"3528",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b84",x"35fd",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"35fd",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2ba0",x"35e4",x"352a",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2b48",x"35f3",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"35f3",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2b7d",x"35d3",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2b0a",x"35f1",x"354a",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"35f1",x"354a",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2b76",x"35bd",x"352b",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"2aba",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"359e",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"35bd",x"3610",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"2aba",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"36f7",x"3576",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2d8d",x"36f7",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2d8d",x"3710",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"380a",x"35cd",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2f8b",x"380a",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b",x"37b8",x"35c0",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"37a8",x"35c3",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ec9",x"37b8",x"35c0",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ee7",x"37a8",x"3578",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"37a8",x"35c3",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"2ec9",x"37a8",x"3578",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"2ec9",x"378c",x"35d3",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"378c",x"35d3",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2e97",x"378c",x"3568",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2e97",x"376c",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"3752",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"376c",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"2e5e",x"3752",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"36e3",x"362f",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"2d6a",x"36f7",x"3638",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e",x"36df",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"36df",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"2d63",x"3716",x"3634",x"3710",x"0000",x"0000",x"3c00",x"3a2f",x"2dc4",x"36dc",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"36e3",x"350c",x"3710",x"0000",x"0000",x"3c00",x"39f0",x"2d6a",x"36df",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"36f7",x"3503",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"36df",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2d63",x"36dc",x"3527",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e",x"3716",x"3507",x"3710",x"0000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"3760",x"3526",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2e49",x"3753",x"3518",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"2e32",x"375f",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"375f",x"3530",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"2e47",x"3742",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2e14",x"3754",x"353b",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"3742",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"3753",x"3623",x"3710",x"0000",x"0000",x"3c00",x"3a2c",x"2e32",x"375f",x"360b",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"372e",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0",x"3742",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2e14",x"3754",x"3600",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"3705",x"35db",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36cb",x"35e6",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2d40",x"36c4",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"36c2",x"354d",x"3710",x"0000",x"0000",x"3c00",x"39fe",x"2d2f",x"36cb",x"3555",x"3710",x"0000",x"0000",x"3c00",x"3a00",x"2d40",x"36c4",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"36c4",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"2d33",x"3705",x"3560",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"2da6",x"36dc",x"3527",x"3710",x"0000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"3713",x"35d4",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3705",x"35db",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"2da6",x"36dc",x"3615",x"3710",x"0000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"3754",x"3600",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"2e33",x"3713",x"35d4",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"372e",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"3754",x"353b",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33",x"372e",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"2df0",x"3713",x"3567",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"3716",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5",x"3713",x"35d4",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"2dbf",x"3752",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"3754",x"353b",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"2e33",x"3713",x"3567",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"2dbf",x"3752",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"3716",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5",x"3710",x"3571",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2dbb",x"3716",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"3716",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2dc5",x"3752",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"2e30",x"3716",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"380a",x"35cd",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"2f8b",x"3813",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"380a",x"356e",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"3813",x"35cf",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"2fac",x"382a",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3813",x"356c",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"382a",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"2ffc",x"382a",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2ffc",x"3885",x"3575",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"3885",x"35c6",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30a2",x"388c",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"3885",x"3575",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"38d5",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130",x"38bf",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38d5",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130"),
(x"38bf",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"3109",x"38bf",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"3109",x"38b2",x"35d6",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"38b2",x"35d6",x"3710",x"0000",x"0000",x"3c00",x"3a1b",x"30f1",x"38b2",x"3565",x"3710",x"0000",x"0000",x"3c00",x"3a03",x"30f1",x"38b0",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38b0",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed",x"38b0",x"355b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed",x"388c",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"386c",x"3541",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3075",x"3872",x"3550",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"386d",x"352c",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3076"),
(x"3872",x"3550",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3080",x"3885",x"3562",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"3877",x"351a",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3088"),
(x"386c",x"35fa",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3075",x"386d",x"3610",x"3710",x"0000",x"0000",x"3c00",x"3a28",x"3076",x"3872",x"35eb",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080"),
(x"3872",x"35eb",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3080",x"3877",x"3621",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3088",x"3885",x"35da",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"3885",x"35da",x"3710",x"0000",x"0000",x"3c00",x"3a1c",x"30a2",x"3894",x"362d",x"3710",x"0000",x"0000",x"3c00",x"3a2e",x"30bc",x"388c",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"3885",x"3562",x"3710",x"0000",x"0000",x"3c00",x"3a02",x"30a2",x"388c",x"356a",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"3894",x"350e",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"38d9",x"3533",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"3136",x"38d8",x"352e",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"3135",x"38d4",x"353c",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d"),
(x"38c7",x"361c",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38d8",x"360d",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3135",x"38d4",x"35ff",x"3710",x"0000",x"0000",x"3c00",x"3a24",x"312d"),
(x"38b7",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38c7",x"361c",x"3710",x"0000",x"0000",x"3c00",x"3a2a",x"3117",x"38c9",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a"),
(x"38d4",x"353c",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"312d",x"38c7",x"351f",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"3117",x"38c9",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a"),
(x"38b2",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"388c",x"356a",x"3710",x"0000",x"0000",x"3c00",x"3a04",x"30ae",x"38b0",x"355b",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"388c",x"35c9",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"30ad",x"388c",x"35d1",x"3710",x"0000",x"0000",x"3c00",x"3a1a",x"30ae",x"38b0",x"35e0",x"3710",x"0000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"38c9",x"3544",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"311a",x"38b7",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38bd",x"3548",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3107"),
(x"38d5",x"35c2",x"3710",x"0000",x"0000",x"3c00",x"3a17",x"3130",x"38f6",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"38d5",x"3579",x"3710",x"0000",x"0000",x"3c00",x"3a07",x"3130"),
(x"38f6",x"35ca",x"3710",x"0000",x"0000",x"3c00",x"3a19",x"316b",x"3915",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"38f6",x"3572",x"3710",x"0000",x"0000",x"3c00",x"3a06",x"316b"),
(x"3915",x"3554",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"31a2",x"3915",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"31a2",x"392f",x"351e",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"392f",x"361d",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"31d0",x"393f",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"392f",x"351e",x"3710",x"0000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"393f",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"31ed",x"3953",x"3620",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"393f",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"3953",x"3620",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3211",x"395a",x"360e",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"3953",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3211"),
(x"395a",x"360e",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"321d",x"395d",x"3602",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"395a",x"352d",x"3710",x"0000",x"0000",x"3c00",x"39f7",x"321d"),
(x"395d",x"3539",x"3710",x"0000",x"0000",x"3c00",x"39fa",x"3222",x"395d",x"3602",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"3222",x"3963",x"3541",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3963",x"35fa",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"322d",x"3972",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3963",x"3541",x"3710",x"0000",x"0000",x"3c00",x"39fc",x"322d"),
(x"3972",x"35fb",x"3710",x"0000",x"0000",x"3c00",x"3a23",x"3248",x"3985",x"360c",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3972",x"3540",x"3710",x"0000",x"0000",x"3c00",x"39fb",x"3248"),
(x"3985",x"352f",x"3710",x"0000",x"0000",x"3c00",x"39f8",x"3269",x"3985",x"360c",x"3710",x"0000",x"0000",x"3c00",x"3a27",x"3269",x"3994",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3994",x"3620",x"3710",x"0000",x"0000",x"3c00",x"3a2b",x"3284",x"3999",x"3622",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"3994",x"351b",x"3710",x"0000",x"0000",x"3c00",x"39f3",x"3284"),
(x"3999",x"3519",x"3710",x"975f",x"9f93",x"3c00",x"39f3",x"328d",x"3999",x"3622",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39fc",x"3571",x"3713",x"ac0e",x"a310",x"3bfb",x"3a06",x"333e"),
(x"3999",x"3622",x"3710",x"935f",x"1e0a",x"3c00",x"3a2c",x"328d",x"39f5",x"3627",x"3710",x"b60a",x"25b5",x"3b67",x"3a2d",x"3331",x"39fb",x"35cc",x"3713",x"a9a8",x"a460",x"3bfd",x"3a19",x"333d"),
(x"3a14",x"3628",x"374f",x"a8f4",x"3bfa",x"ac2a",x"3bcd",x"3a5c",x"3a0d",x"3627",x"374b",x"a412",x"3bfd",x"2966",x"3bce",x"3a59",x"3a1a",x"3628",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e"),
(x"3a1a",x"3628",x"3749",x"a2b5",x"3bfe",x"281b",x"3bcf",x"3a5e",x"3a07",x"3628",x"373c",x"a752",x"3bff",x"9bfc",x"3bd1",x"3a56",x"3a21",x"3629",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60"),
(x"3a21",x"3629",x"373a",x"a884",x"3bfe",x"2546",x"3bd1",x"3a60",x"3a00",x"3627",x"3722",x"23fc",x"3bf8",x"2d56",x"3bd6",x"3a54",x"3a24",x"3629",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62"),
(x"3a24",x"3629",x"372b",x"a504",x"3bff",x"9a24",x"3bd4",x"3a62",x"39fc",x"3627",x"3718",x"135f",x"3bfd",x"29a1",x"3bd8",x"3a52",x"3a27",x"3629",x"3710",x"a3ef",x"3bff",x"9818",x"3bd9",x"3a63"),
(x"3a14",x"3513",x"374e",x"a81b",x"bbe6",x"b0f5",x"3a92",x"3a5c",x"3a19",x"3514",x"3749",x"208e",x"bc00",x"128d",x"3a90",x"3a5e",x"3a0d",x"3514",x"374b",x"1481",x"bbff",x"26a1",x"3a91",x"3a59"),
(x"3a19",x"3514",x"3749",x"208e",x"bc00",x"128d",x"3a90",x"3a5e",x"3a20",x"3513",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a07",x"3513",x"373c",x"0cea",x"bbfe",x"27bb",x"3a8e",x"3a57"),
(x"3a20",x"3513",x"3732",x"1f93",x"bc00",x"975f",x"3a8c",x"3a60",x"3a26",x"3514",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63",x"3a02",x"3513",x"3724",x"1c81",x"bbff",x"a1c9",x"3a89",x"3a55"),
(x"3501",x"3552",x"36da",x"ada6",x"bbf8",x"8000",x"3a6e",x"3b94",x"34e9",x"3558",x"36da",x"b698",x"bb49",x"0000",x"3a6e",x"3b90",x"3501",x"3552",x"3710",x"2d0c",x"bbf9",x"0000",x"3a79",x"3b94"),
(x"386c",x"3541",x"36da",x"bb38",x"36e2",x"8000",x"3a8a",x"3a0c",x"3872",x"3550",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"386c",x"3541",x"3710",x"bbdd",x"31e1",x"0000",x"3a95",x"3a0c"),
(x"380a",x"35cd",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"3813",x"35cf",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"380a",x"35cd",x"3710",x"ae12",x"3bf6",x"0000",x"3aa1",x"39f9"),
(x"34e9",x"3558",x"36da",x"b698",x"bb49",x"0000",x"3a6e",x"3b90",x"34cb",x"356b",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34e9",x"3558",x"3710",x"b50d",x"bb97",x"0000",x"3a79",x"3b90"),
(x"3a26",x"3514",x"36da",x"1e3f",x"bc00",x"0000",x"3a7b",x"3a63",x"39fc",x"3513",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"3a26",x"3514",x"3710",x"1f5f",x"bbff",x"a025",x"3a85",x"3a63"),
(x"3872",x"3550",x"36da",x"b903",x"3a3c",x"0000",x"3a8a",x"3a08",x"3885",x"3562",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"3872",x"3550",x"3710",x"b9d1",x"397d",x"068d",x"3a95",x"3a08"),
(x"3760",x"3615",x"36da",x"3bfa",x"2cac",x"8a8d",x"3a97",x"3a28",x"375f",x"360b",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"3760",x"3615",x"3710",x"3b92",x"3528",x"0000",x"3aa1",x"3a28"),
(x"34cb",x"356b",x"36da",x"b501",x"bb99",x"0000",x"3a6e",x"3b89",x"34bb",x"356f",x"36da",x"b140",x"bbe4",x"0000",x"3a6e",x"3b86",x"34cb",x"356b",x"3710",x"b64c",x"bb5a",x"0000",x"3a79",x"3b89"),
(x"3885",x"3562",x"36da",x"b83d",x"3ac8",x"0000",x"3a8a",x"3a00",x"388c",x"356a",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"3885",x"3562",x"3710",x"b7eb",x"3af3",x"0000",x"3a95",x"3a00"),
(x"37b8",x"35c0",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"380a",x"35cd",x"36da",x"ad56",x"3bf8",x"8000",x"3a97",x"39f9",x"37b8",x"35c0",x"3710",x"30d0",x"3be8",x"0000",x"3aa1",x"3a0b"),
(x"34bb",x"356f",x"36da",x"b140",x"bbe4",x"0000",x"3a6e",x"3b86",x"349b",x"3571",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"34bb",x"356f",x"3710",x"b31c",x"bbcc",x"0000",x"3a79",x"3b86"),
(x"388c",x"356a",x"36da",x"bbfd",x"29ab",x"0000",x"3a8a",x"39fd",x"388c",x"3572",x"36da",x"b967",x"b9e6",x"0000",x"3a8a",x"39fb",x"388c",x"356a",x"3710",x"bb54",x"3669",x"0000",x"3a95",x"39fd"),
(x"37a8",x"35c3",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"37b8",x"35c0",x"36da",x"2df3",x"3bf7",x"8000",x"3a97",x"3a0b",x"37a8",x"35c3",x"3710",x"3580",x"3b83",x"0000",x"3aa1",x"3a0e"),
(x"349b",x"3571",x"36da",x"b4a8",x"bba7",x"8000",x"3a6e",x"3b80",x"3485",x"357a",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"349b",x"3571",x"3710",x"b221",x"bbda",x"0000",x"3a79",x"3b80"),
(x"388c",x"3572",x"36da",x"b967",x"b9e6",x"0000",x"3a7c",x"3bb2",x"3885",x"3575",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"388c",x"3572",x"3710",x"bb52",x"b671",x"0000",x"3a87",x"3bb2"),
(x"378c",x"35d3",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"37a8",x"35c3",x"36da",x"33d5",x"3bc1",x"0000",x"3a97",x"3a0e",x"378c",x"35d3",x"3710",x"3688",x"3b4d",x"0000",x"3aa1",x"3a14"),
(x"3a26",x"35cd",x"36da",x"3311",x"3bcd",x"0000",x"3b16",x"385d",x"3a2f",x"35c9",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"385a",x"3a26",x"35cd",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3864"),
(x"3485",x"357a",x"36da",x"b92c",x"ba1a",x"0000",x"3a6e",x"3b7b",x"3475",x"358c",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3485",x"357a",x"3710",x"b819",x"bade",x"8000",x"3a79",x"3b7b"),
(x"3760",x"3526",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"3753",x"3518",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3760",x"3526",x"3710",x"3bfa",x"acac",x"0000",x"3a87",x"3b52"),
(x"376c",x"35e0",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"378c",x"35d3",x"36da",x"373a",x"3b23",x"0000",x"3a97",x"3a14",x"376c",x"35e0",x"3710",x"3899",x"3a8b",x"0000",x"3aa1",x"3a1a"),
(x"3885",x"3575",x"36da",x"b25f",x"bbd7",x"0000",x"3a7c",x"3baf",x"382a",x"3574",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"3885",x"3575",x"3710",x"b305",x"bbce",x"0000",x"3a87",x"3baf"),
(x"3752",x"35f7",x"36da",x"3bdf",x"31a3",x"8000",x"3a97",x"3a21",x"376c",x"35e0",x"36da",x"3787",x"3b0e",x"0000",x"3a97",x"3a1a",x"3752",x"35f7",x"3710",x"3bfd",x"aabe",x"0000",x"3aa1",x"3a21"),
(x"39fc",x"3513",x"36da",x"a104",x"bc00",x"0000",x"3a7b",x"3a53",x"3999",x"3519",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"39fc",x"3513",x"3710",x"9bc8",x"bc00",x"200b",x"3a85",x"3a53"),
(x"382a",x"3574",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b8d",x"3813",x"356c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"382a",x"3574",x"3710",x"2f40",x"bbf2",x"0000",x"3a87",x"3b8d"),
(x"3742",x"362a",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"3753",x"3623",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3742",x"362a",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"3a2f"),
(x"3813",x"356c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a7c",x"3b84",x"380a",x"356e",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"3813",x"356c",x"3710",x"27fc",x"bbfe",x"0000",x"3a87",x"3b84"),
(x"372e",x"362a",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"3742",x"362a",x"36da",x"342c",x"3bb9",x"8000",x"3a97",x"3a2f",x"372e",x"362a",x"3710",x"338a",x"3bc6",x"0000",x"3aa1",x"3a32"),
(x"375f",x"3530",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"3760",x"3526",x"36da",x"3b92",x"b528",x"0000",x"3a7c",x"3b52",x"375f",x"3530",x"3710",x"3b14",x"3774",x"8000",x"3a87",x"3b54"),
(x"3716",x"3634",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"372e",x"362a",x"36da",x"2fc6",x"3bf0",x"0000",x"3a97",x"3a32",x"3716",x"3634",x"3710",x"32c1",x"3bd1",x"0000",x"3aa1",x"3a37"),
(x"380a",x"356e",x"36da",x"ae12",x"bbf6",x"0000",x"3a7c",x"3b81",x"37b8",x"357b",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"380a",x"356e",x"3710",x"ad56",x"bbf8",x"0000",x"3a87",x"3b81"),
(x"36f7",x"3638",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"3716",x"3634",x"36da",x"34b5",x"3ba5",x"0000",x"3a97",x"3a37",x"36f7",x"3638",x"3710",x"b463",x"3bb1",x"8000",x"3aa1",x"3a3d"),
(x"37b8",x"357b",x"36da",x"30d0",x"bbe8",x"0000",x"3a7c",x"3b6f",x"37a8",x"3578",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"37b8",x"357b",x"3710",x"2df3",x"bbf7",x"0000",x"3a87",x"3b6f"),
(x"36e3",x"362f",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36f7",x"3638",x"36da",x"ae6b",x"3bf5",x"0000",x"3a97",x"3a3d",x"36e3",x"362f",x"3710",x"bb17",x"3766",x"0000",x"3aa1",x"3a41"),
(x"37a8",x"3578",x"36da",x"3580",x"bb83",x"0000",x"3a7c",x"3b6c",x"378c",x"3568",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"37a8",x"3578",x"3710",x"33d5",x"bbc1",x"0000",x"3a87",x"3b6c"),
(x"36df",x"3621",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36e3",x"362f",x"36da",x"b9b5",x"399a",x"8000",x"3a97",x"3a41",x"36df",x"3621",x"3710",x"bbc6",x"338f",x"8000",x"3aa1",x"3a44"),
(x"378c",x"3568",x"36da",x"3688",x"bb4d",x"0000",x"3a7c",x"3b66",x"376c",x"355c",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"378c",x"3568",x"3710",x"373a",x"bb23",x"8000",x"3a87",x"3b66"),
(x"36dc",x"3615",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36df",x"3621",x"36da",x"bbbc",x"3412",x"0000",x"3a97",x"3a44",x"36dc",x"3615",x"3710",x"bb3a",x"36d9",x"0000",x"3aa1",x"3a47"),
(x"3a27",x"3629",x"36da",x"3bff",x"a4d0",x"0000",x"3a2c",x"33f9",x"3a26",x"35cd",x"36da",x"3bff",x"a4d0",x"0000",x"3a18",x"33f3",x"3a27",x"3629",x"3710",x"3bea",x"a4d6",x"30a2",x"3a2c",x"33c9"),
(x"3999",x"3622",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"39f5",x"3627",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"3999",x"3622",x"3710",x"b328",x"3bcb",x"0000",x"3bd9",x"3a2b"),
(x"376c",x"355c",x"36da",x"3899",x"ba8b",x"0000",x"3a7c",x"3b5f",x"3752",x"3544",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"376c",x"355c",x"3710",x"3787",x"bb0e",x"0000",x"3a87",x"3b5f"),
(x"36c4",x"35fb",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36dc",x"3615",x"36da",x"bba4",x"34ba",x"0000",x"3a97",x"3a47",x"36c4",x"35fb",x"3710",x"bbc5",x"339b",x"0000",x"3aa1",x"3a4d"),
(x"3994",x"3620",x"36da",x"b458",x"3bb2",x"0000",x"3be3",x"3a29",x"3999",x"3622",x"36da",x"b2b0",x"3bd2",x"0000",x"3be3",x"3a2b",x"3994",x"3620",x"3710",x"b59f",x"3b7d",x"0000",x"3bd9",x"3a29"),
(x"3753",x"3518",x"36da",x"37e4",x"baf5",x"8000",x"3a7c",x"3b4e",x"3742",x"3511",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"3753",x"3518",x"3710",x"38fe",x"ba3f",x"868d",x"3a87",x"3b4e"),
(x"36c2",x"35ef",x"36da",x"bbe7",x"b0ec",x"868d",x"3a97",x"3a50",x"36c4",x"35fb",x"36da",x"bb61",x"362a",x"0000",x"3a97",x"3a4d",x"36c2",x"35ef",x"3710",x"baff",x"b7c2",x"0000",x"3aa1",x"3a50"),
(x"3985",x"360c",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3994",x"3620",x"36da",x"b458",x"3bb2",x"0000",x"3be3",x"3a29",x"3985",x"360c",x"3710",x"b796",x"3b0b",x"0000",x"3bd9",x"3a22"),
(x"3742",x"3511",x"36da",x"30bd",x"bbe9",x"0000",x"3a7c",x"3b4b",x"372e",x"3511",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"3742",x"3511",x"3710",x"342c",x"bbb9",x"0000",x"3a87",x"3b4b"),
(x"36cb",x"35e6",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"36c2",x"35ef",x"36da",x"bbe7",x"b0ec",x"868d",x"3a97",x"3a50",x"36cb",x"35e6",x"3710",x"b86c",x"baa9",x"0000",x"3aa1",x"3a52"),
(x"3972",x"35fb",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3985",x"360c",x"36da",x"b817",x"3adf",x"0000",x"3be3",x"3a22",x"3972",x"35fb",x"3710",x"b0a0",x"3bea",x"0000",x"3bd9",x"3a1a"),
(x"372e",x"3511",x"36da",x"338a",x"bbc6",x"0000",x"3a7c",x"3b47",x"3716",x"3507",x"36da",x"32c2",x"bbd1",x"0000",x"3a7c",x"3b42",x"372e",x"3511",x"3710",x"2fc6",x"bbf0",x"0000",x"3a87",x"3b47"),
(x"3705",x"35db",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"36cb",x"35e6",x"36da",x"b922",x"ba22",x"8000",x"3a97",x"3a52",x"3705",x"35db",x"3710",x"b675",x"bb51",x"0000",x"3aa1",x"3a5d"),
(x"3963",x"35fa",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"3972",x"35fb",x"36da",x"b475",x"3bae",x"0000",x"3be3",x"3a1a",x"3963",x"35fa",x"3710",x"36c5",x"3b3f",x"0000",x"3bd9",x"3a14"),
(x"3716",x"3507",x"36da",x"32c2",x"bbd1",x"0000",x"3a7c",x"3b42",x"36f7",x"3503",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"3716",x"3507",x"3710",x"34b5",x"bba5",x"0000",x"3a87",x"3b42"),
(x"3713",x"35d4",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3705",x"35db",x"36da",x"b599",x"bb7e",x"8000",x"3a97",x"3a5d",x"3713",x"35d4",x"3710",x"ba37",x"b909",x"0000",x"3aa1",x"3a60"),
(x"395d",x"3602",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"3963",x"35fa",x"36da",x"3420",x"3bba",x"8000",x"3be3",x"3a14",x"395d",x"3602",x"3710",x"3ac1",x"3849",x"0000",x"3bd9",x"3a11"),
(x"36f7",x"3503",x"36da",x"b463",x"bbb1",x"8000",x"3a7c",x"3b3c",x"36e3",x"350c",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36f7",x"3503",x"3710",x"ae6b",x"bbf5",x"8000",x"3a87",x"3b3c"),
(x"3716",x"35cf",x"36da",x"bbb8",x"b42d",x"0000",x"3a97",x"3a61",x"3713",x"35d4",x"36da",x"b972",x"b9db",x"8000",x"3a97",x"3a60",x"3716",x"35cf",x"3710",x"bbad",x"3480",x"0000",x"3aa1",x"3a61"),
(x"395a",x"360e",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"395d",x"3602",x"36da",x"399d",x"39b2",x"0000",x"3be3",x"3a11",x"395a",x"360e",x"3710",x"3af1",x"37f3",x"0000",x"3bd9",x"3a0e"),
(x"36e3",x"350c",x"36da",x"bb17",x"b766",x"868d",x"3a7c",x"3b38",x"36df",x"351a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36e3",x"350c",x"3710",x"b9b5",x"b99a",x"0000",x"3a87",x"3b38"),
(x"3710",x"35ca",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"3716",x"35cf",x"36da",x"bbb8",x"b42d",x"0000",x"3a54",x"39ec",x"3710",x"35ca",x"3710",x"b80e",x"3ae5",x"8000",x"3a5f",x"39ee"),
(x"3953",x"3620",x"36da",x"39a8",x"39a7",x"068d",x"3be3",x"3a09",x"395a",x"360e",x"36da",x"3b46",x"36a7",x"0000",x"3be3",x"3a0e",x"3953",x"3620",x"3710",x"3857",x"3ab8",x"0000",x"3bd9",x"3a09"),
(x"36df",x"351a",x"36da",x"bbc6",x"b38f",x"0000",x"3a7c",x"3b35",x"36dc",x"3527",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36df",x"351a",x"3710",x"bbbc",x"b412",x"8000",x"3a87",x"3b35"),
(x"36f7",x"35c6",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"3710",x"35ca",x"36da",x"b8f7",x"3a45",x"0000",x"3a54",x"39ee",x"36f7",x"35c6",x"3710",x"b05b",x"3bec",x"8000",x"3a5f",x"39f3"),
(x"3475",x"358c",x"36da",x"bbab",x"b48e",x"8000",x"3a6e",x"3b77",x"3475",x"35af",x"36da",x"baeb",x"3803",x"068d",x"3a6e",x"3b70",x"3475",x"358c",x"3710",x"baeb",x"b803",x"068d",x"3a79",x"3b77"),
(x"393f",x"362a",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"3953",x"3620",x"36da",x"39a8",x"39a7",x"068d",x"3be3",x"3a09",x"393f",x"362a",x"3710",x"b2bb",x"3bd2",x"0000",x"3bd9",x"3a01"),
(x"36dc",x"3527",x"36da",x"bb3a",x"b6d9",x"8000",x"3a7c",x"3b33",x"36c4",x"3540",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36dc",x"3527",x"3710",x"bba4",x"b4ba",x"0000",x"3a87",x"3b33"),
(x"362c",x"35ca",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"363b",x"35c5",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"362c",x"35ca",x"3710",x"3609",x"3b68",x"8000",x"3a5f",x"3a19"),
(x"3999",x"3519",x"36da",x"b32c",x"bbcb",x"0000",x"3a7b",x"3a2d",x"3994",x"351b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3999",x"3519",x"3710",x"b2ba",x"bbd2",x"0000",x"3a85",x"3a2d"),
(x"392f",x"361d",x"36da",x"b73b",x"3b22",x"8000",x"3be3",x"39fa",x"393f",x"362a",x"36da",x"1cea",x"3c00",x"8000",x"3be3",x"3a01",x"392f",x"361d",x"3710",x"b874",x"3aa4",x"0000",x"3bd9",x"39fa"),
(x"36c4",x"3540",x"36da",x"bbc5",x"b39b",x"068d",x"3a7c",x"3b2c",x"36c2",x"354d",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36c4",x"3540",x"3710",x"bb61",x"b62a",x"0000",x"3a87",x"3b2c"),
(x"363b",x"35c5",x"36da",x"3439",x"3bb7",x"0000",x"3a54",x"3a16",x"36f7",x"35c6",x"36da",x"b12d",x"3be4",x"0000",x"3a54",x"39f3",x"363b",x"35c5",x"3710",x"34bd",x"3ba4",x"0000",x"3a5f",x"3a16"),
(x"3994",x"351b",x"36da",x"b59f",x"bb7d",x"0000",x"3a7b",x"3a2b",x"3985",x"352f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3994",x"351b",x"3710",x"b458",x"bbb2",x"0000",x"3a85",x"3a2b"),
(x"3754",x"3600",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"3752",x"35f7",x"36da",x"3bdf",x"31a3",x"8000",x"3a97",x"3a21",x"3754",x"3600",x"3710",x"3afe",x"b7c4",x"0000",x"3aa1",x"3a23"),
(x"36c2",x"354d",x"36da",x"bafe",x"37c2",x"8000",x"3a7c",x"3b2a",x"36cb",x"3555",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"36c2",x"354d",x"3710",x"bbe7",x"30ec",x"0000",x"3a87",x"3b2a"),
(x"35f7",x"35e8",x"36da",x"3a05",x"3943",x"8000",x"3a54",x"3a25",x"362c",x"35ca",x"36da",x"3550",x"3b8b",x"0000",x"3a54",x"3a19",x"35f7",x"35e8",x"3710",x"3a6a",x"38c7",x"0000",x"3a5f",x"3a25"),
(x"3985",x"352f",x"36da",x"b796",x"bb0b",x"0000",x"3a7b",x"3a25",x"3972",x"3540",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3985",x"352f",x"3710",x"b817",x"badf",x"0000",x"3a85",x"3a25"),
(x"3915",x"35e8",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"392f",x"361d",x"36da",x"b73b",x"3b22",x"8000",x"3be3",x"39fa",x"3915",x"35e8",x"3710",x"b845",x"3ac3",x"0000",x"3bd9",x"39ec"),
(x"36cb",x"3555",x"36da",x"b86c",x"3aaa",x"0000",x"3a7c",x"3b28",x"3705",x"3560",x"36da",x"b675",x"3b51",x"0000",x"3a7c",x"3b1d",x"36cb",x"3555",x"3710",x"b922",x"3a22",x"868d",x"3a87",x"3b28"),
(x"35f1",x"35f1",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f7",x"35e8",x"36da",x"3a05",x"3943",x"8000",x"3a54",x"3a25",x"35f1",x"35f1",x"3710",x"3bf9",x"ad21",x"0000",x"3a5f",x"3a27"),
(x"3972",x"3540",x"36da",x"b0a0",x"bbea",x"0000",x"3a7b",x"3a1d",x"3963",x"3541",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"3972",x"3540",x"3710",x"b475",x"bbae",x"0000",x"3a85",x"3a1d"),
(x"375f",x"360b",x"36da",x"3b14",x"b774",x"8000",x"3a97",x"3a26",x"3754",x"3600",x"36da",x"3ba5",x"b4b5",x"0000",x"3a97",x"3a23",x"375f",x"360b",x"3710",x"3bc1",x"b3d8",x"0000",x"3aa1",x"3a26"),
(x"3705",x"3560",x"36da",x"b675",x"3b51",x"0000",x"3a7c",x"3b1d",x"3713",x"3567",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3705",x"3560",x"3710",x"b599",x"3b7e",x"0000",x"3a87",x"3b1d"),
(x"35f3",x"35f7",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35f1",x"35f1",x"36da",x"3bcd",x"3318",x"0000",x"3a54",x"3a27",x"35f3",x"35f7",x"3710",x"3b36",x"b6ea",x"0000",x"3a5f",x"3a28"),
(x"3963",x"3541",x"36da",x"36c5",x"bb3f",x"0000",x"3a7b",x"3a17",x"395d",x"3539",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"3963",x"3541",x"3710",x"3420",x"bbba",x"0000",x"3a85",x"3a17"),
(x"38f6",x"35ca",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"3915",x"35e8",x"36da",x"b90a",x"3a36",x"0000",x"3be3",x"39ec",x"38f6",x"35ca",x"3710",x"b324",x"3bcc",x"0000",x"3bd9",x"39de"),
(x"3713",x"3567",x"36da",x"ba37",x"3909",x"0000",x"3a7c",x"3b1a",x"3716",x"356c",x"36da",x"bbad",x"b480",x"0000",x"3a7c",x"3b19",x"3713",x"3567",x"3710",x"b972",x"39db",x"0000",x"3a87",x"3b1a"),
(x"35fd",x"3605",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35f3",x"35f7",x"36da",x"3b84",x"b57a",x"0000",x"3a54",x"3a28",x"35fd",x"3605",x"3710",x"3bf0",x"aff4",x"068d",x"3a5f",x"3a2b"),
(x"395d",x"3539",x"36da",x"3ac1",x"b849",x"0000",x"3a7b",x"3a14",x"395a",x"352d",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"395d",x"3539",x"3710",x"399d",x"b9b2",x"0000",x"3a85",x"3a14"),
(x"38d5",x"35c2",x"36da",x"1953",x"3c00",x"0000",x"3be3",x"39d1",x"38f6",x"35ca",x"36da",x"b551",x"3b8b",x"0000",x"3be3",x"39de",x"38d5",x"35c2",x"3710",x"2dde",x"3bf7",x"0000",x"3bd9",x"39d1"),
(x"3716",x"356c",x"36da",x"bbad",x"b480",x"0000",x"3afb",x"3a11",x"3710",x"3571",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"3716",x"356c",x"3710",x"bbb8",x"342e",x"0000",x"3b06",x"3a11"),
(x"35fd",x"360e",x"36da",x"3b87",x"3567",x"068d",x"3a54",x"3a2d",x"35fd",x"3605",x"36da",x"3b91",x"b530",x"8000",x"3a54",x"3a2b",x"35fd",x"360e",x"3710",x"3a08",x"3941",x"0000",x"3a5f",x"3a2d"),
(x"395a",x"352d",x"36da",x"3af1",x"b7f3",x"8000",x"3a7b",x"3a12",x"3953",x"351b",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"395a",x"352d",x"3710",x"3b46",x"b6a7",x"868d",x"3a85",x"3a12"),
(x"38bf",x"35c9",x"36da",x"3489",x"3bac",x"0000",x"3be3",x"39c8",x"38d5",x"35c2",x"36da",x"1953",x"3c00",x"0000",x"3be3",x"39d1",x"38bf",x"35c9",x"3710",x"35f3",x"3b6d",x"0000",x"3bd9",x"39c8"),
(x"3710",x"3571",x"36da",x"b80d",x"bae5",x"8000",x"3afb",x"3a0f",x"36f7",x"3576",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"3710",x"3571",x"3710",x"b8f7",x"ba45",x"0000",x"3b06",x"3a0f"),
(x"35f5",x"3613",x"36da",x"364b",x"3b5a",x"868d",x"3a54",x"3a2e",x"35fd",x"360e",x"36da",x"3b87",x"3567",x"068d",x"3a54",x"3a2d",x"35f5",x"3613",x"3710",x"32d5",x"3bd0",x"8000",x"3a5f",x"3a2e"),
(x"3953",x"351b",x"36da",x"3857",x"bab8",x"8000",x"3a7b",x"3a0d",x"393f",x"3511",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"3953",x"351b",x"3710",x"39a8",x"b9a7",x"0000",x"3a85",x"3a0d"),
(x"38b2",x"35d6",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38bf",x"35c9",x"36da",x"3489",x"3bac",x"0000",x"3be3",x"39c8",x"38b2",x"35d6",x"3710",x"3af2",x"37f0",x"0000",x"3bd9",x"39c2"),
(x"363b",x"3576",x"36da",x"34be",x"bba4",x"0000",x"3afb",x"39e7",x"362c",x"3571",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"363b",x"3576",x"3710",x"3439",x"bbb7",x"868d",x"3b06",x"39e7"),
(x"35e4",x"3612",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35f5",x"3613",x"36da",x"364b",x"3b5a",x"868d",x"3a54",x"3a2e",x"35e4",x"3612",x"3710",x"b3c4",x"3bc2",x"8000",x"3a5f",x"3a32"),
(x"393f",x"3511",x"36da",x"b2bb",x"bbd2",x"0000",x"3a7b",x"3a05",x"392f",x"351e",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"393f",x"3511",x"3710",x"1d04",x"bc00",x"0000",x"3a85",x"3a05"),
(x"38b0",x"35e0",x"36da",x"3bfc",x"2b2b",x"0000",x"3be3",x"39c0",x"38b2",x"35d6",x"36da",x"3a0a",x"393e",x"8000",x"3be3",x"39c2",x"38b0",x"35e0",x"3710",x"3ba6",x"b4ab",x"0000",x"3bd9",x"39c0"),
(x"36f7",x"3576",x"36da",x"b05b",x"bbec",x"0000",x"3afb",x"3a0a",x"363b",x"3576",x"36da",x"34be",x"bba4",x"0000",x"3afb",x"39e7",x"36f7",x"3576",x"3710",x"b12d",x"bbe4",x"0000",x"3b06",x"3a0a"),
(x"35d3",x"360b",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35e4",x"3612",x"36da",x"b0fa",x"3be7",x"0000",x"3a54",x"3a32",x"35d3",x"360b",x"3710",x"1c81",x"3c00",x"0000",x"3a5f",x"3a35"),
(x"3752",x"3544",x"36da",x"3bfd",x"2ac2",x"0000",x"3a7c",x"3b59",x"3754",x"353b",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"3752",x"3544",x"3710",x"3be0",x"b1a3",x"0000",x"3a87",x"3b59"),
(x"38b2",x"35e8",x"36da",x"3a58",x"b8de",x"0000",x"3be3",x"39be",x"38b0",x"35e0",x"36da",x"3bfc",x"2b2b",x"0000",x"3be3",x"39c0",x"38b2",x"35e8",x"3710",x"399c",x"b9b3",x"8000",x"3bd9",x"39be"),
(x"362c",x"3571",x"36da",x"3609",x"bb68",x"8000",x"3afb",x"39e4",x"35f7",x"3553",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"362c",x"3571",x"3710",x"3550",x"bb8b",x"0000",x"3b06",x"39e4"),
(x"35bd",x"3610",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"35d3",x"360b",x"36da",x"b1d2",x"3bdd",x"0000",x"3a54",x"3a35",x"35bd",x"3610",x"3710",x"afcb",x"3bf0",x"8000",x"3a5f",x"3a39"),
(x"392f",x"351e",x"36da",x"b874",x"baa4",x"0000",x"3a7b",x"39ff",x"3915",x"3554",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"392f",x"351e",x"3710",x"b73b",x"bb22",x"0000",x"3a85",x"39ff"),
(x"38bd",x"35f3",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38b2",x"35e8",x"36da",x"3a58",x"b8de",x"0000",x"3a7d",x"3ac5",x"38bd",x"35f3",x"3710",x"3456",x"bbb3",x"0000",x"3a87",x"3ac9"),
(x"35f7",x"3553",x"36da",x"3a6a",x"b8c7",x"0000",x"3afb",x"39d8",x"35f1",x"354a",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f7",x"3553",x"3710",x"3a05",x"b943",x"0000",x"3b06",x"39d8"),
(x"359e",x"3605",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"35bd",x"3610",x"36da",x"2c74",x"3bfb",x"068d",x"3a54",x"3a39",x"359e",x"3605",x"3710",x"b925",x"3a1f",x"0000",x"3a5f",x"3a40"),
(x"3754",x"353b",x"36da",x"3afe",x"37c4",x"0000",x"3a7c",x"3b57",x"375f",x"3530",x"36da",x"3bc1",x"33d7",x"8000",x"3a7c",x"3b54",x"3754",x"353b",x"3710",x"3ba5",x"34b5",x"0000",x"3a87",x"3b57"),
(x"38c9",x"35f7",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38bd",x"35f3",x"36da",x"35fc",x"bb6b",x"0000",x"3a7d",x"3ac9",x"38c9",x"35f7",x"3710",x"34cb",x"bba1",x"0000",x"3a87",x"3ace"),
(x"35f1",x"354a",x"36da",x"3bf9",x"2d21",x"0000",x"3afb",x"39d6",x"35f3",x"3544",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35f1",x"354a",x"3710",x"3bcd",x"b318",x"0000",x"3b06",x"39d6"),
(x"358a",x"35ee",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"359e",x"3605",x"36da",x"b80b",x"3ae7",x"8000",x"3a54",x"3a40",x"358a",x"35ee",x"3710",x"bbad",x"3481",x"0000",x"3a5f",x"3a45"),
(x"3915",x"3554",x"36da",x"b845",x"bac3",x"0000",x"3a7b",x"39f1",x"38f6",x"3572",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"3915",x"3554",x"3710",x"b90a",x"ba36",x"0000",x"3a85",x"39f1"),
(x"38d4",x"35ff",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38c9",x"35f7",x"36da",x"3385",x"bbc6",x"8000",x"3a7d",x"3ace",x"38d4",x"35ff",x"3710",x"38a8",x"ba80",x"8000",x"3a87",x"3ad2"),
(x"35f3",x"3544",x"36da",x"3b36",x"36ea",x"8000",x"3afb",x"39d5",x"35fd",x"3536",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35f3",x"3544",x"3710",x"3b84",x"357a",x"0000",x"3b06",x"39d5"),
(x"3587",x"35d9",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"358a",x"35ee",x"36da",x"bb1e",x"374c",x"8000",x"3a54",x"3a45",x"3587",x"35d9",x"3710",x"bb8b",x"b553",x"0000",x"3a5f",x"3a49"),
(x"38f6",x"3572",x"36da",x"b324",x"bbcc",x"0000",x"3a7b",x"39e4",x"38d5",x"3579",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38f6",x"3572",x"3710",x"b551",x"bb8b",x"0000",x"3a85",x"39e4"),
(x"38d9",x"3608",x"36da",x"3b87",x"b565",x"0000",x"3a7d",x"3ad5",x"38d4",x"35ff",x"36da",x"37f2",x"baf1",x"0000",x"3a7d",x"3ad2",x"38d9",x"3608",x"3710",x"3bfc",x"ab00",x"868d",x"3a87",x"3ad5"),
(x"3a25",x"356e",x"36da",x"3bff",x"26b5",x"0000",x"3a09",x"33f0",x"3a26",x"3514",x"36da",x"3bff",x"26b5",x"0000",x"39f5",x"33fa",x"3a25",x"356e",x"3710",x"3bd6",x"2604",x"3256",x"3a07",x"33c0"),
(x"35fd",x"3536",x"36da",x"3bf0",x"2ff4",x"8000",x"3afb",x"39d2",x"35fd",x"352d",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35fd",x"3536",x"3710",x"3b91",x"3530",x"8000",x"3b06",x"39d2"),
(x"3593",x"35c7",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3587",x"35d9",x"36da",x"bbf7",x"adba",x"8000",x"3a54",x"3a49",x"3593",x"35c7",x"3710",x"bc00",x"15bc",x"0000",x"3a5f",x"3a4d"),
(x"38d5",x"3579",x"36da",x"2dde",x"bbf7",x"0000",x"3a7b",x"39d7",x"38bf",x"3572",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38d5",x"3579",x"3710",x"1987",x"bc00",x"0000",x"3a85",x"39d7"),
(x"38d8",x"360d",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38d9",x"3608",x"36da",x"3b87",x"b565",x"0000",x"3a7d",x"3ad5",x"38d8",x"360d",x"3710",x"3b96",x"350f",x"0000",x"3a87",x"3ad6"),
(x"35fd",x"352d",x"36da",x"3a08",x"b941",x"868d",x"3afb",x"39d0",x"35f5",x"3528",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35fd",x"352d",x"3710",x"3b87",x"b567",x"8000",x"3b06",x"39d0"),
(x"3592",x"35bf",x"36da",x"bba4",x"34bb",x"0000",x"3a54",x"3a4f",x"3593",x"35c7",x"36da",x"bbda",x"b21b",x"0000",x"3a54",x"3a4d",x"3592",x"35bf",x"3710",x"ba08",x"3941",x"0000",x"3a5f",x"3a4f"),
(x"38bf",x"3572",x"36da",x"35f3",x"bb6c",x"0000",x"3a7b",x"39cf",x"38b2",x"3565",x"36da",x"3af2",x"b7f0",x"0000",x"3a7b",x"39c9",x"38bf",x"3572",x"3710",x"3489",x"bbab",x"0000",x"3a85",x"39cf"),
(x"38c7",x"361c",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38d8",x"360d",x"36da",x"3be4",x"312f",x"8000",x"3a7d",x"3ad6",x"38c7",x"361c",x"3710",x"364a",x"3b5b",x"0000",x"3a87",x"3add"),
(x"35f5",x"3528",x"36da",x"32d5",x"bbd0",x"8000",x"3afb",x"39ce",x"35e4",x"352a",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35f5",x"3528",x"3710",x"364b",x"bb5a",x"068d",x"3b06",x"39ce"),
(x"357d",x"35bd",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"3592",x"35bf",x"36da",x"bba4",x"34bb",x"0000",x"3a6e",x"3b35",x"357d",x"35bd",x"3710",x"26c2",x"3bff",x"0000",x"3a79",x"3b39"),
(x"38b2",x"3565",x"36da",x"3af2",x"b7f0",x"0000",x"3a8a",x"3a50",x"38b0",x"355b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b2",x"3565",x"3710",x"3a0a",x"b93e",x"8000",x"3a95",x"3a50"),
(x"38b7",x"362a",x"36da",x"3528",x"3b92",x"068d",x"3a7d",x"3ae4",x"38c7",x"361c",x"36da",x"3654",x"3b58",x"8000",x"3a7d",x"3add",x"38b7",x"362a",x"3710",x"32f7",x"3bce",x"8000",x"3a87",x"3ae4"),
(x"35e4",x"352a",x"36da",x"b3c4",x"bbc2",x"0000",x"3afb",x"39cb",x"35d3",x"3530",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35e4",x"352a",x"3710",x"b0fa",x"bbe7",x"0000",x"3b06",x"39cb"),
(x"3555",x"35c2",x"36da",x"345b",x"3bb2",x"0000",x"3a6e",x"3b41",x"357d",x"35bd",x"36da",x"a8c9",x"3bfe",x"0000",x"3a6e",x"3b39",x"3555",x"35c2",x"3710",x"35eb",x"3b6e",x"0000",x"3a79",x"3b41"),
(x"38b0",x"355b",x"36da",x"3ba6",x"34ac",x"0000",x"3a8a",x"3a4d",x"38b2",x"3553",x"36da",x"399c",x"39b3",x"8000",x"3a8a",x"3a4c",x"38b0",x"355b",x"3710",x"3bfc",x"ab27",x"0000",x"3a95",x"3a4d"),
(x"3894",x"362d",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"38b7",x"362a",x"36da",x"3528",x"3b92",x"068d",x"3a7d",x"3ae4",x"3894",x"362d",x"3710",x"b036",x"3bee",x"0000",x"3a87",x"3af1"),
(x"35d3",x"3530",x"36da",x"1c81",x"bc00",x"0000",x"3afb",x"39c8",x"35bd",x"352b",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"35d3",x"3530",x"3710",x"b1d2",x"bbdd",x"0000",x"3b06",x"39c8"),
(x"353f",x"35cd",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"3555",x"35c2",x"36da",x"345b",x"3bb2",x"0000",x"3a6e",x"3b41",x"353f",x"35cd",x"3710",x"379f",x"3b08",x"0000",x"3a79",x"3b46"),
(x"38b2",x"3553",x"36da",x"399c",x"39b3",x"8000",x"3a8a",x"3a4c",x"38bd",x"3548",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38b2",x"3553",x"3710",x"3a58",x"38de",x"0000",x"3a95",x"3a4c"),
(x"3877",x"3621",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"3894",x"362d",x"36da",x"aa0a",x"3bfd",x"8000",x"3a7d",x"3af1",x"3877",x"3621",x"3710",x"b8aa",x"3a7f",x"8000",x"3a87",x"3afc"),
(x"35bd",x"352b",x"36da",x"afc9",x"bbf0",x"0000",x"3afb",x"39c3",x"359e",x"3536",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"35bd",x"352b",x"3710",x"2c74",x"bbfb",x"0000",x"3b06",x"39c3"),
(x"351b",x"35e2",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"353f",x"35cd",x"36da",x"3746",x"3b1f",x"0000",x"3a6e",x"3b46",x"351b",x"35e2",x"3710",x"350e",x"3b96",x"0000",x"3a79",x"3b4e"),
(x"38bd",x"3548",x"36da",x"3456",x"3bb3",x"0000",x"3a8a",x"3a47",x"38c9",x"3544",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38bd",x"3548",x"3710",x"35fc",x"3b6b",x"0000",x"3a95",x"3a47"),
(x"386d",x"3610",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"3877",x"3621",x"36da",x"b74e",x"3b1d",x"0000",x"3a7d",x"3afc",x"386d",x"3610",x"3710",x"bba8",x"34a3",x"0000",x"3a87",x"3b01"),
(x"359e",x"3536",x"36da",x"b925",x"ba1f",x"8000",x"3afb",x"39bd",x"358a",x"354d",x"36da",x"bbad",x"b481",x"8000",x"3afb",x"39b7",x"359e",x"3536",x"3710",x"b80b",x"bae7",x"8000",x"3b06",x"39bd"),
(x"3501",x"35e9",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"351b",x"35e2",x"36da",x"3664",x"3b55",x"8000",x"3a6e",x"3b4e",x"3501",x"35e9",x"3710",x"ada6",x"3bf8",x"8000",x"3a79",x"3b53"),
(x"38c9",x"3544",x"36da",x"34cb",x"3ba1",x"8000",x"3a8a",x"3a43",x"38d4",x"353c",x"36da",x"38a8",x"3a80",x"0000",x"3a8a",x"3a3e",x"38c9",x"3544",x"3710",x"3385",x"3bc6",x"0000",x"3a95",x"3a43"),
(x"386c",x"35fa",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"386d",x"3610",x"36da",x"bac4",x"3844",x"8000",x"3a7d",x"3b01",x"386c",x"35fa",x"3710",x"bb38",x"b6e2",x"0000",x"3a87",x"3b05"),
(x"358a",x"354d",x"36da",x"bbad",x"b481",x"8000",x"3afb",x"39b7",x"3587",x"3562",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"358a",x"354d",x"3710",x"bb1e",x"b74c",x"8000",x"3b06",x"39b7"),
(x"34e9",x"35e3",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"3501",x"35e9",x"36da",x"2d0c",x"3bf9",x"8000",x"3a6e",x"3b53",x"34e9",x"35e3",x"3710",x"b698",x"3b49",x"0000",x"3a79",x"3b57"),
(x"38d4",x"353c",x"36da",x"38a8",x"3a80",x"0000",x"3a8a",x"3a3e",x"38d9",x"3533",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d4",x"353c",x"3710",x"37f2",x"3af1",x"0000",x"3a95",x"3a3e"),
(x"3872",x"35eb",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"386c",x"35fa",x"36da",x"bbdd",x"b1e1",x"0000",x"3a7d",x"3b05",x"3872",x"35eb",x"3710",x"b902",x"ba3c",x"0000",x"3a87",x"3b08"),
(x"3587",x"3562",x"36da",x"bb8b",x"3553",x"0000",x"3afb",x"39b3",x"3593",x"3574",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3587",x"3562",x"3710",x"bbf7",x"2dba",x"068d",x"3b06",x"39b3"),
(x"34cb",x"35d1",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34e9",x"35e3",x"36da",x"b50d",x"3b97",x"8000",x"3a6e",x"3b57",x"34cb",x"35d1",x"3710",x"b501",x"3b99",x"0000",x"3a79",x"3b5e"),
(x"38d9",x"3533",x"36da",x"3bfc",x"2b00",x"8000",x"3a8a",x"3a3c",x"38d8",x"352e",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38d9",x"3533",x"3710",x"3b88",x"3564",x"0000",x"3a95",x"3a3c"),
(x"3885",x"35da",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"3872",x"35eb",x"36da",x"b9d1",x"b97d",x"8000",x"3a7d",x"3b08",x"3885",x"35da",x"3710",x"b83d",x"bac8",x"0000",x"3a87",x"3b10"),
(x"3593",x"3574",x"36da",x"bc00",x"95bc",x"0000",x"3afb",x"39af",x"3592",x"357c",x"36da",x"ba08",x"b941",x"8000",x"3afb",x"39ae",x"3593",x"3574",x"3710",x"bbda",x"321b",x"0000",x"3b06",x"39af"),
(x"34bb",x"35cc",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"34cb",x"35d1",x"36da",x"b64c",x"3b5a",x"0000",x"3a6e",x"3b5e",x"34bb",x"35cc",x"3710",x"b141",x"3be4",x"0000",x"3a79",x"3b61"),
(x"38d8",x"352e",x"36da",x"3b96",x"b50f",x"0000",x"3a8a",x"3a3b",x"38c7",x"351f",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38d8",x"352e",x"3710",x"3be4",x"b12f",x"8a8d",x"3a95",x"3a3b"),
(x"388c",x"35d1",x"36da",x"bb54",x"b669",x"0000",x"3a7d",x"3b13",x"3885",x"35da",x"36da",x"b7eb",x"baf3",x"0000",x"3a7d",x"3b10",x"388c",x"35d1",x"3710",x"bbfd",x"a9ab",x"0000",x"3a87",x"3b13"),
(x"3592",x"357c",x"36da",x"ba08",x"b941",x"8000",x"3a6e",x"3bb2",x"357d",x"357e",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"3592",x"357c",x"3710",x"bba4",x"b4bb",x"0000",x"3a79",x"3bb2"),
(x"349b",x"35ca",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"34bb",x"35cc",x"36da",x"b31c",x"3bcc",x"0000",x"3a6e",x"3b61",x"349b",x"35ca",x"3710",x"b4a8",x"3ba7",x"0000",x"3a79",x"3b67"),
(x"38c7",x"351f",x"36da",x"364a",x"bb5b",x"0000",x"3a8a",x"3a34",x"38b7",x"3511",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"38c7",x"351f",x"3710",x"3653",x"bb59",x"0000",x"3a95",x"3a34"),
(x"388c",x"35c9",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"388c",x"35d1",x"36da",x"bb54",x"b669",x"0000",x"3a97",x"39c6",x"388c",x"35c9",x"3710",x"b967",x"39e6",x"0000",x"3aa1",x"39c8"),
(x"357d",x"357e",x"36da",x"26bb",x"bbff",x"0000",x"3a6e",x"3bae",x"3555",x"3579",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"357d",x"357e",x"3710",x"a8c9",x"bbfe",x"0000",x"3a79",x"3bae"),
(x"3485",x"35c1",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"349b",x"35ca",x"36da",x"b221",x"3bda",x"8000",x"3a6e",x"3b67",x"3485",x"35c1",x"3710",x"b92c",x"3a1a",x"8000",x"3a79",x"3b6c"),
(x"38b7",x"3511",x"36da",x"32f7",x"bbce",x"0000",x"3a8a",x"3a2d",x"3894",x"350e",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"38b7",x"3511",x"3710",x"3528",x"bb92",x"8000",x"3a95",x"3a2d"),
(x"3885",x"35c6",x"36da",x"b305",x"3bce",x"0000",x"3a97",x"39ca",x"388c",x"35c9",x"36da",x"bb52",x"3671",x"0000",x"3a97",x"39c8",x"3885",x"35c6",x"3710",x"b25f",x"3bd7",x"0000",x"3aa1",x"39ca"),
(x"3555",x"3579",x"36da",x"35eb",x"bb6e",x"0000",x"3a6e",x"3ba6",x"353f",x"356e",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"3555",x"3579",x"3710",x"345a",x"bbb2",x"0000",x"3a79",x"3ba6"),
(x"3475",x"35af",x"36da",x"baeb",x"3803",x"068d",x"3a6e",x"3b70",x"3485",x"35c1",x"36da",x"b819",x"3ade",x"8000",x"3a6e",x"3b6c",x"3475",x"35af",x"3710",x"bbab",x"348e",x"0000",x"3a79",x"3b70"),
(x"3894",x"350e",x"36da",x"b036",x"bbee",x"0000",x"3a8a",x"3a20",x"3877",x"351a",x"36da",x"b8aa",x"ba7f",x"068d",x"3a8a",x"3a15",x"3894",x"350e",x"3710",x"aa0a",x"bbfd",x"0000",x"3a95",x"3a20"),
(x"3753",x"3623",x"36da",x"38fe",x"3a3f",x"8000",x"3a97",x"3a2b",x"3760",x"3615",x"36da",x"3bfa",x"2cac",x"8a8d",x"3a97",x"3a28",x"3753",x"3623",x"3710",x"37e4",x"3af5",x"8000",x"3aa1",x"3a2b"),
(x"3a2f",x"35c9",x"36da",x"3bfe",x"a8f0",x"0000",x"3be9",x"39cf",x"3a2d",x"3576",x"36da",x"3bfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"3a2f",x"35c9",x"3710",x"3b78",x"a99e",x"35b0",x"3be8",x"39da"),
(x"353f",x"356e",x"36da",x"379f",x"bb08",x"0000",x"3a6e",x"3ba2",x"351b",x"3559",x"36da",x"350e",x"bb96",x"068d",x"3a6e",x"3b9a",x"353f",x"356e",x"3710",x"3746",x"bb1f",x"0000",x"3a79",x"3ba2"),
(x"39f5",x"3627",x"36da",x"a49b",x"3bff",x"8000",x"3be3",x"3a4f",x"3a27",x"3629",x"36da",x"a3ae",x"3bff",x"0000",x"3be3",x"3a63",x"39f5",x"3627",x"3710",x"a4e3",x"3bff",x"17c8",x"3bd9",x"3a4f"),
(x"3877",x"351a",x"36da",x"b8aa",x"ba7f",x"068d",x"3a8a",x"3a15",x"386d",x"352c",x"36da",x"bba8",x"b4a3",x"8000",x"3a8a",x"3a10",x"3877",x"351a",x"3710",x"b74e",x"bb1d",x"0000",x"3a95",x"3a15"),
(x"382a",x"35c7",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"3885",x"35c6",x"36da",x"b305",x"3bce",x"0000",x"3a97",x"39ca",x"382a",x"35c7",x"3710",x"30bd",x"3be9",x"0000",x"3aa1",x"39ed"),
(x"351b",x"3559",x"36da",x"350e",x"bb96",x"068d",x"3a6e",x"3b9a",x"3501",x"3552",x"36da",x"ada6",x"bbf8",x"8000",x"3a6e",x"3b94",x"351b",x"3559",x"3710",x"3664",x"bb55",x"8000",x"3a79",x"3b9a"),
(x"386d",x"352c",x"36da",x"bba8",x"b4a3",x"8000",x"3a8a",x"3a10",x"386c",x"3541",x"36da",x"bb38",x"36e2",x"8000",x"3a8a",x"3a0c",x"386d",x"352c",x"3710",x"bac4",x"b844",x"8000",x"3a95",x"3a10"),
(x"3813",x"35cf",x"36da",x"27fc",x"3bfe",x"0000",x"3a97",x"39f5",x"382a",x"35c7",x"36da",x"2f40",x"3bf2",x"0000",x"3a97",x"39ed",x"3813",x"35cf",x"3710",x"a8bf",x"3bfe",x"0000",x"3aa1",x"39f5"),
(x"3a2d",x"3576",x"36da",x"367a",x"bb50",x"0000",x"3bbd",x"3982",x"3a25",x"356e",x"36da",x"367a",x"bb50",x"0000",x"3bc0",x"3984",x"3a2d",x"3576",x"3710",x"3644",x"bb4c",x"2f83",x"3bb7",x"398a"),
(x"38b2",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"30f2",x"38b7",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38bd",x"35f3",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3107"),
(x"3592",x"35bf",x"3710",x"0000",x"0000",x"3c00",x"3a16",x"2a20",x"3593",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"359e",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"358a",x"354d",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2a0e",x"3593",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27"),
(x"359e",x"3536",x"3710",x"0000",x"0000",x"3c00",x"39f9",x"2a4d",x"3593",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"2f99",x"39db",x"36b4",x"0000",x"0000",x"3c00",x"3a8e",x"3516",x"3004",x"39d4",x"36b4",x"0000",x"0000",x"3c00",x"3a90",x"351d",x"3009",x"39cc",x"36b4",x"0000",x"0000",x"3c00",x"3a92",x"351d"),
(x"2fe5",x"39c1",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"351a",x"2f19",x"39d7",x"36b4",x"0000",x"0000",x"3c00",x"3a8f",x"350d",x"2f99",x"39db",x"36b4",x"0000",x"0000",x"3c00",x"3a8e",x"3516"),
(x"2f10",x"39c0",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"350c",x"2ee6",x"39cd",x"36b4",x"0000",x"0000",x"3c00",x"3a91",x"3509",x"2f19",x"39d7",x"36b4",x"0000",x"0000",x"3c00",x"3a8f",x"350d"),
(x"2fda",x"39bb",x"36b4",x"0000",x"0000",x"3c00",x"3a96",x"3519",x"2f02",x"397e",x"36b4",x"0000",x"0000",x"3c00",x"3aa2",x"3508",x"2f10",x"39c0",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"350c"),
(x"2fda",x"39bb",x"36b4",x"0000",x"0000",x"3c00",x"3a96",x"3519",x"3025",x"397f",x"36b4",x"0000",x"0000",x"3c00",x"3aa3",x"351e",x"2f02",x"397e",x"36b4",x"0000",x"0000",x"3c00",x"3aa2",x"3508"),
(x"2fe5",x"39c1",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"351a",x"2f10",x"39c0",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"350c",x"2f19",x"39d7",x"36b4",x"0000",x"0000",x"3c00",x"3a8f",x"350d"),
(x"2f99",x"39db",x"36b4",x"0000",x"0000",x"3c00",x"3a8e",x"3516",x"3009",x"39cc",x"36b4",x"0000",x"0000",x"3c00",x"3a92",x"351d",x"2fe5",x"39c1",x"36b4",x"0000",x"0000",x"3c00",x"3a94",x"351a"),
(x"358a",x"3c9f",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"2a04",x"359e",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"3593",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"38b7",x"3c68",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38b2",x"3c79",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"38bd",x"3c76",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3107"),
(x"38b7",x"3cae",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38c9",x"3ca1",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a",x"38bd",x"3ca0",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3107"),
(x"3593",x"3c95",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22",x"359e",x"3ca5",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"35f7",x"3c9e",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"358a",x"3c77",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2a0e",x"3587",x"3c7c",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2a04",x"3593",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27"),
(x"3593",x"3c81",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27",x"3592",x"3c83",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20",x"35f7",x"3c78",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"358a",x"35ee",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"2a04",x"359e",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"3593",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"38b7",x"3511",x"3710",x"0000",x"0000",x"3c00",x"39f1",x"30f9",x"38b2",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"30f2",x"38bd",x"3548",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"3107"),
(x"38b7",x"362a",x"3710",x"0000",x"0000",x"3c00",x"3a2d",x"30f9",x"38c9",x"35f7",x"3710",x"0000",x"0000",x"3c00",x"3a22",x"311a",x"38bd",x"35f3",x"3710",x"0000",x"0000",x"3c00",x"3a20",x"3107"),
(x"3593",x"35c7",x"3710",x"0000",x"0000",x"3c00",x"3a18",x"2a22",x"359e",x"3605",x"3710",x"0000",x"0000",x"3c00",x"3a25",x"2a4d",x"35f7",x"35e8",x"3710",x"0000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"358a",x"354d",x"3710",x"0000",x"0000",x"3c00",x"39fd",x"2a0e",x"3587",x"3562",x"3710",x"0000",x"0000",x"3c00",x"3a01",x"2a04",x"3593",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27"),
(x"3593",x"3574",x"3710",x"0000",x"0000",x"3c00",x"3a05",x"2a27",x"3592",x"357c",x"3710",x"0000",x"0000",x"3c00",x"3a08",x"2a20",x"35f7",x"3553",x"3710",x"0000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b936",x"3cc1",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"3a68",x"b936",x"34b8",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"38f3",x"b936",x"3cc1",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"3a68"),
(x"2af5",x"39ca",x"36b2",x"3c00",x"0000",x"0000",x"371d",x"30fe",x"2af5",x"39ca",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30fe",x"2af5",x"3cc1",x"368e",x"3c00",x"0000",x"0000",x"3732",x"345d"),
(x"aaef",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3af7",x"3815",x"aaef",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3af7",x"3810",x"b858",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3a04",x"3815"),
(x"b936",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3a0a",x"b936",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3a0a",x"2af5",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3b6a"),
(x"2af5",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"3ada",x"b936",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"397a",x"2af5",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"3ada"),
(x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"b86b",x"3c28",x"36fb",x"8000",x"0000",x"3c00",x"3aff",x"3bb2",x"b86c",x"376a",x"36fb",x"8000",x"0000",x"3c00",x"3aff",x"3ad6"),
(x"9da8",x"39d4",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3b",x"9e2f",x"39cc",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3a",x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1"),
(x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96",x"b936",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3a96",x"aaef",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3ac4"),
(x"b858",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3bbd",x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"aaef",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3bbd"),
(x"aaef",x"36aa",x"36d0",x"8000",x"0000",x"3c00",x"35d1",x"3ae0",x"b858",x"36aa",x"36d0",x"8000",x"0000",x"3c00",x"346e",x"3ae0",x"aaef",x"3c44",x"36d0",x"8000",x"0000",x"3c00",x"35d1",x"3bfa"),
(x"aaef",x"36aa",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"370d",x"36e5",x"bc00",x"0000",x"0000",x"3ae4",x"3545",x"aaef",x"36e5",x"36fb",x"bc00",x"0000",x"0000",x"3ae5",x"3546"),
(x"b858",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3a05",x"3821",x"b858",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3a05",x"3826",x"aaef",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3af8",x"3821"),
(x"a9a6",x"3c25",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8",x"aaef",x"3c28",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"aa60",x"3c38",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1"),
(x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96",x"aaef",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3ac4",x"aa24",x"3716",x"36fb",x"8000",x"0000",x"3c00",x"3bc4",x"3ace"),
(x"aa60",x"3c38",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1",x"aaef",x"3c37",x"36e4",x"ba1e",x"b322",x"38d5",x"351b",x"38d1",x"aaef",x"3c41",x"36fb",x"b9d6",x"b5ae",x"38ac",x"351f",x"38d6"),
(x"aaef",x"36aa",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"3c44",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"3743",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545"),
(x"aaef",x"3c44",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"3c44",x"36fb",x"bc00",x"0000",x"0000",x"3a7f",x"3557",x"aaef",x"3c41",x"36fb",x"bc00",x"0000",x"0000",x"3a83",x"3557"),
(x"a9ae",x"374d",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3ad3",x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96",x"aa24",x"3716",x"36fb",x"8000",x"0000",x"3c00",x"3bc4",x"3ace"),
(x"a9ae",x"374d",x"36fb",x"b993",x"1c9b",x"39bd",x"3526",x"3740",x"aaef",x"3743",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"a9a6",x"3c25",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8"),
(x"aaef",x"370d",x"36e5",x"b96c",x"347c",x"396f",x"351c",x"3730",x"aaef",x"3743",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"aa24",x"3716",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"aaef",x"36e5",x"36fb",x"b969",x"359e",x"392e",x"351f",x"3725",x"aaef",x"370d",x"36e5",x"b96c",x"347c",x"396f",x"351c",x"3730",x"aa24",x"3716",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"b857",x"3c37",x"36e5",x"3bfe",x"2104",x"a780",x"3b41",x"34eb",x"b857",x"3c42",x"36fb",x"3bfe",x"276c",x"a4f7",x"3b42",x"34ec",x"b858",x"3c44",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9"),
(x"b858",x"36aa",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b858",x"36aa",x"36fb",x"3bff",x"a5e9",x"0000",x"3ad1",x"34ff",x"b857",x"36db",x"36fb",x"3bff",x"a3a0",x"a0dd",x"3ade",x"3501"),
(x"b863",x"3709",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0",x"b857",x"3709",x"36dd",x"3a1a",x"3321",x"38da",x"357e",x"38d0",x"b857",x"36db",x"36fb",x"39d1",x"35ef",x"389e",x"3584",x"38d6"),
(x"b857",x"3c28",x"36d8",x"3bf1",x"15bc",x"afa2",x"3b3f",x"34eb",x"b858",x"3c44",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b857",x"3761",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed"),
(x"b86c",x"376a",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4",x"b857",x"3761",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b863",x"3709",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0"),
(x"b86b",x"3c28",x"36fb",x"3935",x"9d6d",x"3a12",x"3587",x"373c",x"b857",x"3c28",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b86c",x"376a",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4"),
(x"b857",x"3c37",x"36e5",x"397e",x"b36f",x"3983",x"357d",x"372e",x"b857",x"3c28",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b862",x"3c37",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"b857",x"3c42",x"36fb",x"3958",x"b562",x"394e",x"3580",x"3722",x"b857",x"3c37",x"36e5",x"397e",x"b36f",x"3983",x"357d",x"372e",x"b862",x"3c37",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"2163",x"397e",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b2b",x"20f3",x"39c0",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b38",x"2243",x"39cd",x"36fb",x"8000",x"0000",x"3c00",x"3bdc",x"3b3a"),
(x"b936",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3a79",x"30b7",x"2af5",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3b35",x"30b7",x"b936",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3a79",x"290e"),
(x"9ac5",x"39c1",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"9e2f",x"39cc",x"36fb",x"3b8f",x"3538",x"868d",x"3a18",x"3614",x"9ac5",x"39c1",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603"),
(x"2163",x"397e",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a47",x"a0d7",x"397f",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a51",x"2163",x"397e",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a47"),
(x"20b0",x"39d7",x"36fb",x"b727",x"bb27",x"0000",x"3a23",x"3614",x"2243",x"39cd",x"36fb",x"bbcf",x"b2e8",x"8000",x"3a26",x"3614",x"20b0",x"39d7",x"36b4",x"b93c",x"ba0c",x"0000",x"3a23",x"3603"),
(x"9e2f",x"39cc",x"36fb",x"3b8f",x"3538",x"868d",x"3a18",x"3614",x"9da8",x"39d4",x"36fb",x"3aa7",x"b870",x"8000",x"3a1b",x"3614",x"9e2f",x"39cc",x"36b4",x"3bef",x"3011",x"0000",x"3a18",x"3603"),
(x"a0d7",x"397f",x"36fb",x"3bcb",x"b335",x"0000",x"3a04",x"3614",x"995f",x"39bb",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"a0d7",x"397f",x"36b4",x"3bcb",x"b335",x"0000",x"3a04",x"3603"),
(x"2243",x"39cd",x"36fb",x"bbcf",x"b2e8",x"8000",x"3a26",x"3614",x"20f3",x"39c0",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"2243",x"39cd",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603"),
(x"9da8",x"39d4",x"36fb",x"3aa7",x"b870",x"8000",x"3a1b",x"3614",x"1557",x"39db",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"9da8",x"39d4",x"36b4",x"38fa",x"ba42",x"068d",x"3a1b",x"3603"),
(x"995f",x"39bb",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"9ac5",x"39c1",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"995f",x"39bb",x"36b4",x"3be8",x"b0e3",x"868d",x"3a14",x"3603"),
(x"20f3",x"39c0",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"2163",x"397e",x"36fb",x"bbff",x"a6cf",x"0000",x"3a3b",x"3614",x"20f3",x"39c0",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603"),
(x"1557",x"39db",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"20b0",x"39d7",x"36fb",x"b727",x"bb27",x"0000",x"3a23",x"3614",x"1557",x"39db",x"36b4",x"a8d9",x"bbfe",x"0000",x"3a1f",x"3603"),
(x"9ac5",x"39c1",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a18",x"20f3",x"39c0",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a12",x"995f",x"39bb",x"36b4",x"8000",x"0000",x"3c00",x"3b69",x"3a18"),
(x"2af5",x"399f",x"36b2",x"3c00",x"0000",x"0000",x"371d",x"30d2",x"2af5",x"39ca",x"36b2",x"3c00",x"0000",x"0000",x"371d",x"30fe",x"2af5",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"3732",x"2a26"),
(x"2af5",x"34b8",x"36fb",x"3c00",x"0000",x"0000",x"36f3",x"2a26",x"2af5",x"399f",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30d2",x"2af5",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"3732",x"2a26"),
(x"2975",x"399f",x"36b2",x"3c00",x"0000",x"0000",x"3b75",x"396a",x"2975",x"399f",x"36d6",x"3c00",x"0000",x"0000",x"3b75",x"396e",x"2975",x"39ca",x"36b2",x"3c00",x"0000",x"0000",x"3b81",x"396a"),
(x"2af5",x"399f",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a4e",x"2975",x"399f",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a48",x"2af5",x"39ca",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a4e"),
(x"2af5",x"399f",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30d2",x"2af5",x"34b8",x"36fb",x"3c00",x"0000",x"0000",x"36f3",x"2a26",x"2af5",x"39ca",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30fe"),
(x"2af5",x"39ca",x"36b2",x"0000",x"bc00",x"0000",x"3b98",x"396e",x"2975",x"39ca",x"36b2",x"0000",x"bc00",x"0000",x"3b9e",x"396e",x"2af5",x"39ca",x"36d6",x"0000",x"bc00",x"0000",x"3b98",x"396a"),
(x"2af5",x"399f",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"39a5",x"2975",x"399f",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"399f",x"2af5",x"399f",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"39a5"),
(x"2af5",x"39ca",x"36d6",x"0000",x"19f0",x"bc00",x"3b80",x"3a4b",x"2975",x"39ca",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a4b",x"2af5",x"399f",x"36d6",x"0000",x"19f0",x"bc00",x"3b80",x"3a41"),
(x"b936",x"34b8",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"38f3",x"b936",x"34b8",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"38f3",x"b936",x"3cc1",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"3a68"),
(x"2af5",x"39ca",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30fe",x"2af5",x"3cc1",x"36fb",x"3c00",x"0000",x"0000",x"36f3",x"345d",x"2af5",x"3cc1",x"368e",x"3c00",x"0000",x"0000",x"3732",x"345d"),
(x"aaef",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3af7",x"3810",x"b858",x"3c44",x"36d0",x"0000",x"bc00",x"0000",x"3a04",x"3810",x"b858",x"3c44",x"36fb",x"0000",x"bc00",x"0000",x"3a04",x"3815"),
(x"b936",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3a0a",x"2af5",x"34b8",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3b6a",x"2af5",x"34b8",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3b6a"),
(x"b936",x"3cc1",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"397a",x"b936",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"397a",x"2af5",x"3cc1",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"3ada"),
(x"b863",x"3709",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3acd",x"b858",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3ac4",x"b936",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3a96"),
(x"b863",x"3709",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3acd",x"b857",x"36db",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3ac9",x"b858",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3ac4"),
(x"b862",x"3c37",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3bb8",x"b858",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3bbd",x"b857",x"3c42",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3bbc"),
(x"b862",x"3c37",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3bb8",x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"b858",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3bbd"),
(x"b86c",x"376a",x"36fb",x"8000",x"0000",x"3c00",x"3aff",x"3ad6",x"b863",x"3709",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3acd",x"b936",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3a96"),
(x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"b862",x"3c37",x"36fb",x"8000",x"0000",x"3c00",x"3b01",x"3bb8",x"b86b",x"3c28",x"36fb",x"8000",x"0000",x"3c00",x"3aff",x"3bb2"),
(x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"b86c",x"376a",x"36fb",x"8000",x"0000",x"3c00",x"3aff",x"3ad6",x"b936",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3a96"),
(x"aa60",x"3c38",x"36fb",x"8000",x"0000",x"3c00",x"3bc3",x"3bb8",x"aaef",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3bbd",x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb"),
(x"aa60",x"3c38",x"36fb",x"8000",x"0000",x"3c00",x"3bc3",x"3bb8",x"aaef",x"3c41",x"36fb",x"068d",x"0000",x"3c00",x"3bc2",x"3bbb",x"aaef",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3bbd"),
(x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb",x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96",x"2243",x"39cd",x"36fb",x"8000",x"0000",x"3c00",x"3bdc",x"3b3a"),
(x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb",x"2243",x"39cd",x"36fb",x"8000",x"0000",x"3c00",x"3bdc",x"3b3a",x"20b0",x"39d7",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b3c"),
(x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1",x"aa60",x"3c38",x"36fb",x"8000",x"0000",x"3c00",x"3bc3",x"3bb8",x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb"),
(x"a0d7",x"397f",x"36fb",x"8000",x"0000",x"3c00",x"3bd3",x"3b2b",x"a9ae",x"374d",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3ad3",x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1"),
(x"9e2f",x"39cc",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3a",x"995f",x"39bb",x"36fb",x"8000",x"0000",x"3c00",x"3bd6",x"3b37",x"a0d7",x"397f",x"36fb",x"8000",x"0000",x"3c00",x"3bd3",x"3b2b"),
(x"9e2f",x"39cc",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3a",x"9ac5",x"39c1",x"36fb",x"8000",x"0000",x"3c00",x"3bd6",x"3b38",x"995f",x"39bb",x"36fb",x"8000",x"0000",x"3c00",x"3bd6",x"3b37"),
(x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1",x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb",x"20b0",x"39d7",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b3c"),
(x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1",x"20b0",x"39d7",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b3c",x"1557",x"39db",x"36fb",x"8000",x"0000",x"3c00",x"3bd7",x"3b3d"),
(x"9e2f",x"39cc",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3a",x"a0d7",x"397f",x"36fb",x"8000",x"0000",x"3c00",x"3bd3",x"3b2b",x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1"),
(x"a9a6",x"3c25",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3bb1",x"1557",x"39db",x"36fb",x"8000",x"0000",x"3c00",x"3bd7",x"3b3d",x"9da8",x"39d4",x"36fb",x"8000",x"0000",x"3c00",x"3bd5",x"3b3b"),
(x"b936",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3a96",x"b858",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3b03",x"3ac4",x"aaef",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3ac4"),
(x"b936",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3ad9",x"3beb",x"2af5",x"3cc1",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3beb",x"aaef",x"3c44",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3bbd"),
(x"b858",x"36aa",x"36d0",x"8000",x"0000",x"3c00",x"346e",x"3ae0",x"b858",x"3c44",x"36d0",x"8000",x"0000",x"3c00",x"346e",x"3bfa",x"aaef",x"3c44",x"36d0",x"8000",x"0000",x"3c00",x"35d1",x"3bfa"),
(x"aaef",x"36e5",x"36fb",x"bc00",x"0000",x"0000",x"3ae5",x"3546",x"aaef",x"36aa",x"36fb",x"bc00",x"0000",x"0000",x"3ae8",x"3545",x"aaef",x"36aa",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542"),
(x"aaef",x"36aa",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"3743",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545",x"aaef",x"370d",x"36e5",x"bc00",x"0000",x"0000",x"3ae4",x"3545"),
(x"b858",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3a05",x"3826",x"aaef",x"36aa",x"36d0",x"0000",x"3c00",x"0000",x"3af8",x"3826",x"aaef",x"36aa",x"36fb",x"0000",x"3c00",x"0000",x"3af8",x"3821"),
(x"aaef",x"3c28",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"aaef",x"3c37",x"36e4",x"ba1e",x"b322",x"38d5",x"351b",x"38d1",x"aa60",x"3c38",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1"),
(x"aaef",x"36aa",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3ac4",x"aaef",x"36e5",x"36fb",x"8000",x"0000",x"3c00",x"3bc2",x"3aca",x"aa24",x"3716",x"36fb",x"8000",x"0000",x"3c00",x"3bc4",x"3ace"),
(x"aaef",x"3c44",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"3c28",x"36d7",x"bc00",x"0000",x"0000",x"3a9d",x"3546",x"aaef",x"3743",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545"),
(x"aaef",x"3c37",x"36e4",x"bc00",x"0000",x"0000",x"3a8d",x"354c",x"aaef",x"3c28",x"36d7",x"bc00",x"0000",x"0000",x"3a9d",x"3546",x"aaef",x"3c44",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542"),
(x"aaef",x"3c44",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"3c41",x"36fb",x"bc00",x"0000",x"0000",x"3a83",x"3557",x"aaef",x"3c37",x"36e4",x"bc00",x"0000",x"0000",x"3a8d",x"354c"),
(x"aaef",x"3743",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"aaef",x"3c28",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"a9a6",x"3c25",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8"),
(x"aaef",x"3743",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"a9ae",x"374d",x"36fb",x"b993",x"1c9b",x"39bd",x"3526",x"3740",x"aa24",x"3716",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"b858",x"3c44",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b857",x"3c28",x"36d8",x"3bf1",x"15bc",x"afa2",x"3b3f",x"34eb",x"b857",x"3c37",x"36e5",x"3bfe",x"2104",x"a780",x"3b41",x"34eb"),
(x"b857",x"3c42",x"36fb",x"3bfe",x"276c",x"a4f7",x"3b42",x"34ec",x"b858",x"3c44",x"36fb",x"3bf4",x"2eb8",x"0000",x"3b42",x"34eb",x"b858",x"3c44",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9"),
(x"b857",x"3709",x"36dd",x"3bff",x"a074",x"a611",x"3aec",x"34f3",x"b857",x"3761",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed",x"b858",x"36aa",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9"),
(x"b858",x"36aa",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b857",x"36db",x"36fb",x"3bff",x"a3a0",x"a0dd",x"3ade",x"3501",x"b857",x"3709",x"36dd",x"3bff",x"a074",x"a611",x"3aec",x"34f3"),
(x"b858",x"3c44",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b858",x"36aa",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b857",x"3761",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed"),
(x"b857",x"3761",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b857",x"3709",x"36dd",x"3a1a",x"3321",x"38da",x"357e",x"38d0",x"b863",x"3709",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0"),
(x"b857",x"3c28",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b857",x"3761",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b86c",x"376a",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4"),
(x"b857",x"3c28",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b86b",x"3c28",x"36fb",x"3935",x"9d6d",x"3a12",x"3587",x"373c",x"b862",x"3c37",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"2163",x"397e",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b2b",x"a9ae",x"374d",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3ad3",x"a0d7",x"397f",x"36fb",x"8000",x"0000",x"3c00",x"3bd3",x"3b2b"),
(x"2163",x"397e",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b2b",x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96",x"a9ae",x"374d",x"36fb",x"8000",x"0000",x"3c00",x"3bc6",x"3ad3"),
(x"2163",x"397e",x"36fb",x"8000",x"0000",x"3c00",x"3bdb",x"3b2b",x"2243",x"39cd",x"36fb",x"8000",x"0000",x"3c00",x"3bdc",x"3b3a",x"2af5",x"34b8",x"36fb",x"8000",x"0000",x"3c00",x"3bec",x"3a96"),
(x"2af5",x"34b8",x"368e",x"0000",x"8000",x"bc00",x"3b35",x"30b7",x"2af5",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3b35",x"290e",x"b936",x"3cc1",x"368e",x"0000",x"8000",x"bc00",x"3a79",x"290e"),
(x"9e2f",x"39cc",x"36fb",x"3b8f",x"3538",x"868d",x"3a18",x"3614",x"9e2f",x"39cc",x"36b4",x"3bef",x"3011",x"0000",x"3a18",x"3603",x"9ac5",x"39c1",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603"),
(x"a0d7",x"397f",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a51",x"a0d7",x"397f",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a51",x"2163",x"397e",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a47"),
(x"2243",x"39cd",x"36fb",x"bbcf",x"b2e8",x"8000",x"3a26",x"3614",x"2243",x"39cd",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603",x"20b0",x"39d7",x"36b4",x"b93c",x"ba0c",x"0000",x"3a23",x"3603"),
(x"9da8",x"39d4",x"36fb",x"3aa7",x"b870",x"8000",x"3a1b",x"3614",x"9da8",x"39d4",x"36b4",x"38fa",x"ba42",x"068d",x"3a1b",x"3603",x"9e2f",x"39cc",x"36b4",x"3bef",x"3011",x"0000",x"3a18",x"3603"),
(x"995f",x"39bb",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"995f",x"39bb",x"36b4",x"3be8",x"b0e3",x"868d",x"3a14",x"3603",x"a0d7",x"397f",x"36b4",x"3bcb",x"b335",x"0000",x"3a04",x"3603"),
(x"20f3",x"39c0",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"20f3",x"39c0",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603",x"2243",x"39cd",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603"),
(x"1557",x"39db",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"1557",x"39db",x"36b4",x"a8d9",x"bbfe",x"0000",x"3a1f",x"3603",x"9da8",x"39d4",x"36b4",x"38fa",x"ba42",x"068d",x"3a1b",x"3603"),
(x"9ac5",x"39c1",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"9ac5",x"39c1",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603",x"995f",x"39bb",x"36b4",x"3be8",x"b0e3",x"868d",x"3a14",x"3603"),
(x"2163",x"397e",x"36fb",x"bbff",x"a6cf",x"0000",x"3a3b",x"3614",x"2163",x"397e",x"36b4",x"bbff",x"a6cf",x"0000",x"3a3b",x"3603",x"20f3",x"39c0",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603"),
(x"20b0",x"39d7",x"36fb",x"b727",x"bb27",x"0000",x"3a23",x"3614",x"20b0",x"39d7",x"36b4",x"b93c",x"ba0c",x"0000",x"3a23",x"3603",x"1557",x"39db",x"36b4",x"a8d9",x"bbfe",x"0000",x"3a1f",x"3603"),
(x"9da8",x"39d4",x"36b4",x"8000",x"0000",x"3c00",x"3b63",x"3a1a",x"1557",x"39db",x"36b4",x"8000",x"0000",x"3c00",x"3b61",x"3a16",x"9e2f",x"39cc",x"36b4",x"8000",x"0000",x"3c00",x"3b65",x"3a1a"),
(x"20b0",x"39d7",x"36b4",x"8000",x"0000",x"3c00",x"3b62",x"3a12",x"9ac5",x"39c1",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a18",x"1557",x"39db",x"36b4",x"8000",x"0000",x"3c00",x"3b61",x"3a16"),
(x"2243",x"39cd",x"36b4",x"8000",x"0000",x"3c00",x"3b65",x"3a11",x"20f3",x"39c0",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a12",x"20b0",x"39d7",x"36b4",x"8000",x"0000",x"3c00",x"3b62",x"3a12"),
(x"2163",x"397e",x"36b4",x"8000",x"0000",x"3c00",x"3b79",x"3a11",x"995f",x"39bb",x"36b4",x"8000",x"0000",x"3c00",x"3b69",x"3a18",x"20f3",x"39c0",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a12"),
(x"a0d7",x"397f",x"36b4",x"8000",x"0000",x"3c00",x"3b79",x"3a1b",x"995f",x"39bb",x"36b4",x"8000",x"0000",x"3c00",x"3b69",x"3a18",x"2163",x"397e",x"36b4",x"8000",x"0000",x"3c00",x"3b79",x"3a11"),
(x"20f3",x"39c0",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a12",x"9ac5",x"39c1",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a18",x"20b0",x"39d7",x"36b4",x"8000",x"0000",x"3c00",x"3b62",x"3a12"),
(x"9e2f",x"39cc",x"36b4",x"8000",x"0000",x"3c00",x"3b65",x"3a1a",x"1557",x"39db",x"36b4",x"8000",x"0000",x"3c00",x"3b61",x"3a16",x"9ac5",x"39c1",x"36b4",x"8000",x"0000",x"3c00",x"3b68",x"3a18"),
(x"2af5",x"39ca",x"36b2",x"3c00",x"0000",x"0000",x"371d",x"30fe",x"2af5",x"3cc1",x"368e",x"3c00",x"0000",x"0000",x"3732",x"345d",x"2af5",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"3732",x"2a26"),
(x"2af5",x"399f",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30d2",x"2af5",x"399f",x"36b2",x"3c00",x"0000",x"0000",x"371d",x"30d2",x"2af5",x"34b8",x"368e",x"3c00",x"0000",x"0000",x"3732",x"2a26"),
(x"2975",x"399f",x"36d6",x"3c00",x"0000",x"0000",x"3b75",x"396e",x"2975",x"39ca",x"36d6",x"3c00",x"0000",x"0000",x"3b81",x"396e",x"2975",x"39ca",x"36b2",x"3c00",x"0000",x"0000",x"3b81",x"396a"),
(x"2975",x"399f",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a48",x"2975",x"39ca",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a48",x"2af5",x"39ca",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a4e"),
(x"2af5",x"34b8",x"36fb",x"3c00",x"0000",x"0000",x"36f3",x"2a26",x"2af5",x"3cc1",x"36fb",x"3c00",x"0000",x"0000",x"36f3",x"345d",x"2af5",x"39ca",x"36d6",x"3c00",x"0000",x"0000",x"3709",x"30fe"),
(x"2975",x"39ca",x"36b2",x"0000",x"bc00",x"0000",x"3b9e",x"396e",x"2975",x"39ca",x"36d6",x"0000",x"bc00",x"0000",x"3b9e",x"396a",x"2af5",x"39ca",x"36d6",x"0000",x"bc00",x"0000",x"3b98",x"396a"),
(x"2975",x"399f",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"399f",x"2975",x"399f",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"399f",x"2af5",x"399f",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"39a5"),
(x"2975",x"39ca",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a4b",x"2975",x"399f",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a41",x"2af5",x"399f",x"36d6",x"0000",x"19f0",x"bc00",x"3b80",x"3a41"),
(x"b931",x"3c69",x"3710",x"bbe9",x"26a1",x"309e",x"39f4",x"33ca",x"b930",x"3c7f",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0",x"b92b",x"3c69",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa"),
(x"b92b",x"3c69",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa",x"b92a",x"3c7f",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b924",x"3c69",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392"),
(x"b924",x"3c69",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392",x"b922",x"3c7f",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b91f",x"3c69",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387"),
(x"b91f",x"3c69",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387",x"b91b",x"3c7f",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b918",x"3c69",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b"),
(x"b907",x"3c80",x"3713",x"2f5f",x"3bdb",x"30c1",x"3bc0",x"39a6",x"b913",x"3c7f",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b90e",x"3c81",x"370e",x"3754",x"3ae5",x"32eb",x"3bbd",x"39a7"),
(x"b91b",x"3c81",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b913",x"3c81",x"373a",x"3ae3",x"2b4f",x"380a",x"3bb9",x"399f",x"b91b",x"3c7f",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b"),
(x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b906",x"3c69",x"3710",x"2e12",x"a66c",x"3bf6",x"39f2",x"333e",x"b90c",x"3c68",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352"),
(x"b90f",x"3c96",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7",x"b90d",x"3c96",x"3711",x"3be1",x"a6cf",x"3179",x"3be9",x"39fb",x"b90e",x"3c81",x"370e",x"3bcb",x"a949",x"330f",x"3bf9",x"39fa"),
(x"b91a",x"3c96",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b913",x"3c96",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b91b",x"3c81",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed"),
(x"b922",x"3c96",x"3751",x"a11e",x"aa52",x"3bfd",x"3be8",x"39eb",x"b91a",x"3c96",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b924",x"3c82",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b92b",x"3c81",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6",x"b928",x"3c96",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b924",x"3c82",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b930",x"3c81",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3",x"b92f",x"3c96",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b92b",x"3c81",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6"),
(x"b938",x"3c81",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b935",x"3c96",x"3725",x"bb50",x"a63f",x"3678",x"3be8",x"39de",x"b930",x"3c81",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3"),
(x"b935",x"3c96",x"3725",x"bb50",x"a63f",x"3678",x"3be8",x"39de",x"b938",x"3c81",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b93a",x"3c96",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3be8",x"39da"),
(x"b938",x"3c81",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a",x"b930",x"3c81",x"3738",x"b75a",x"bae5",x"32d3",x"3bb5",x"3992",x"b930",x"3c7f",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c"),
(x"b912",x"3c69",x"373c",x"3aea",x"2832",x"3802",x"39f2",x"336a",x"b918",x"3c69",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b",x"b913",x"3c7f",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369"),
(x"b924",x"3c82",x"374d",x"b1ce",x"b808",x"3ac1",x"3bb5",x"3999",x"b91b",x"3c81",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b922",x"3c7f",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998"),
(x"b924",x"3c82",x"374d",x"b1ce",x"b808",x"3ac1",x"3bb5",x"3999",x"b922",x"3c7f",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998",x"b92b",x"3c81",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b92a",x"3c7f",x"3733",x"b800",x"ba99",x"3436",x"3bb7",x"3993",x"b930",x"3c81",x"3738",x"b75a",x"bae5",x"32d3",x"3bb5",x"3992",x"b92b",x"3c81",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b92a",x"3c97",x"3739",x"b604",x"3b4b",x"3148",x"3b22",x"386b",x"b935",x"3c96",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b931",x"3c97",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b925",x"3c97",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e",x"b92f",x"3c96",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b92a",x"3c97",x"3739",x"b604",x"3b4b",x"3148",x"3b22",x"386b"),
(x"b920",x"3c97",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871",x"b928",x"3c96",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e",x"b925",x"3c97",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e"),
(x"b920",x"3c97",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871",x"b922",x"3c96",x"3751",x"9ac2",x"39ac",x"39a3",x"3b24",x"3871",x"b928",x"3c96",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e"),
(x"b919",x"3c97",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873",x"b91a",x"3c96",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b920",x"3c97",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871"),
(x"b913",x"3c98",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875",x"b913",x"3c96",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b919",x"3c97",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873"),
(x"b90b",x"3c97",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879",x"b90f",x"3c96",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879",x"b913",x"3c98",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875"),
(x"b90b",x"3c97",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879",x"b90d",x"3c96",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"387b",x"b90f",x"3c96",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879"),
(x"b906",x"3c97",x"3713",x"2edc",x"bb7b",x"3565",x"3b16",x"387a",x"b90d",x"3c96",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"387b",x"b90b",x"3c97",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879"),
(x"b90e",x"3c81",x"370e",x"b4eb",x"a6e9",x"3b9c",x"3a06",x"334b",x"b90d",x"3c96",x"3711",x"b36d",x"a40b",x"3bc7",x"3a19",x"3349",x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b931",x"3cae",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9",x"b92f",x"3cae",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b931",x"3c97",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4"),
(x"b92a",x"3c97",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b92f",x"3cae",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b92c",x"3cae",x"373a",x"baa5",x"a5fd",x"3872",x"3a2d",x"33a3"),
(x"b925",x"3c97",x"3746",x"b918",x"a84d",x"3a28",x"3a1a",x"338e",x"b92a",x"3c97",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b925",x"3cae",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b91f",x"3cae",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385",x"b920",x"3c97",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b925",x"3cae",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b918",x"3cad",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a2d",x"3378",x"b919",x"3c97",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b91f",x"3cae",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385"),
(x"b911",x"3cae",x"373c",x"3ac9",x"a6b5",x"383a",x"3a2d",x"3366",x"b913",x"3c98",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b918",x"3cad",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a2d",x"3378"),
(x"b90b",x"3c97",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b913",x"3c98",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b90b",x"3cad",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c"),
(x"b906",x"3c97",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b90b",x"3c97",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b907",x"3cae",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340"),
(x"b135",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b116",x"3c8f",x"3710",x"8000",x"0000",x"3c00",x"3a13",x"2451",x"b135",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"b161",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b135",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b161",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f"),
(x"b1a1",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2643",x"b161",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b1a1",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643"),
(x"b1a1",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2643",x"b1a1",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643",x"b1c1",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"b1fd",x"3c9d",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"278b",x"b1c1",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3",x"b1fd",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b"),
(x"b1fd",x"3c9d",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"278b",x"b1fd",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b",x"b22d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"b261",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b22d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a",x"b261",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878"),
(x"b2aa",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b261",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b2aa",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"b2d6",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b2aa",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b2d6",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949"),
(x"b326",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b2d6",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b326",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"b34f",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20",x"b326",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b34f",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"b451",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2c3f",x"b451",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b50c",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"b441",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b451",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b441",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b441",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b34f",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20",x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b34f",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"b413",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2ba0",x"b40b",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b84",x"b413",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"b413",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0",x"b3f4",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b409",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"b409",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d",x"b3d2",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b407",x"3ca0",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"b3f4",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b40b",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b84",x"b413",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"b3d2",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b3f4",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b409",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"b3a5",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b3d2",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b407",x"3c76",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"b368",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b3a5",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b407",x"3ca0",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76",x"b3a5",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b368",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b340",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"2a04",x"b351",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b526",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2dbb",x"b50c",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d",x"b526",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"b5ce",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2ee7",x"b62a",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b",x"b5ce",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"b5ce",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2ee7",x"b5ce",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7",x"b5bd",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"b5a1",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b5bd",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9",x"b5a1",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"b581",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2e5e",x"b5a1",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b581",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"b581",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2e5e",x"b581",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e",x"b568",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b52b",x"3cb1",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b50d",x"3cb2",x"3710",x"8000",x"0000",x"3c00",x"3a30",x"2d8e",x"b4f5",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"b544",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0",x"b52b",x"3cb1",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b4f2",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b52b",x"3c65",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4",x"b4f5",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b50d",x"3c65",x"3710",x"8000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"b544",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b4f2",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b52b",x"3c65",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"b558",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b568",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2e32",x"b575",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"b544",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b558",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b569",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"b575",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2e49",x"b568",x"3cad",x"3710",x"8000",x"0000",x"3c00",x"3a2c",x"2e32",x"b575",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"b575",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47",x"b558",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b569",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"b4d8",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2d2f",x"b4e1",x"3c9d",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2d40",x"b4da",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"b51a",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4e1",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"2d40",x"b4da",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"b528",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b51a",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4f2",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"b4da",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33",x"b51a",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b4f2",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b4f2",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e",x"b528",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b544",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"b4f2",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b544",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b528",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"b569",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33",x"b528",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b568",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"b52c",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5",x"b528",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b568",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b526",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2dbb",x"b526",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb",x"b52c",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"b568",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30",x"b568",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b52c",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"b63d",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac",x"b63d",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b62a",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"b669",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2ffc",x"b669",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b63d",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"b721",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30a2",x"b669",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b721",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b72d",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b72d",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b721",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b794",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"3109",x"b794",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b7c0",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130"),
(x"b77a",x"3c7d",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b794",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b77a",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"b776",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b77a",x"3c7d",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b776",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b72d",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b776",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b72d",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"b705",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088",x"b6fb",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b6f1",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3076"),
(x"b73e",x"3c67",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc",x"b721",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b705",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088"),
(x"b705",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b6f1",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"3076",x"b6fb",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080"),
(x"b73e",x"3caf",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b705",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b721",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"b783",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b73e",x"3caf",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b72e",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b783",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b72e",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b73e",x"3c67",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"b7a4",x"3c6c",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7c7",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3135",x"b7bd",x"3c73",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d"),
(x"b7c7",x"3ca6",x"3710",x"8000",x"0000",x"3c00",x"3a26",x"3136",x"b7c7",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3135",x"b7bd",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d"),
(x"b7bd",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d",x"b7a4",x"3cab",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b7a8",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a"),
(x"b783",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b7a4",x"3c6c",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7a8",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a"),
(x"b72d",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b72e",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b776",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"b77b",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b72e",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae",x"b776",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b783",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b77b",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b72e",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae"),
(x"b77b",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b783",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b72e",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b801",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b",x"b801",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b7c0",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130"),
(x"b820",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"31a2",x"b820",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b801",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b"),
(x"b83a",x"3cab",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"31d0",x"b820",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b83a",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b84a",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed",x"b84a",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b83a",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b85e",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211",x"b85e",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b84a",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"b865",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d",x"b865",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b85e",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211"),
(x"b867",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"3222",x"b867",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b865",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d"),
(x"b86e",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"322d",x"b867",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b86e",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b87d",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248",x"b87d",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b86e",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b88f",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"3269",x"b88f",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b87d",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248"),
(x"b89e",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3284",x"b88f",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b89e",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b8a3",x"3c6a",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b8a3",x"3cac",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b89e",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b906",x"3c97",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b8a3",x"3cac",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b907",x"3cae",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340",x"b8ff",x"3cae",x"3710",x"2904",x"26d5",x"3bfd",x"3a2d",x"3331",x"b906",x"3c97",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d"),
(x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b8a3",x"3c6a",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b906",x"3c69",x"3710",x"2e12",x"a66c",x"3bf6",x"39f2",x"333e"),
(x"b911",x"3cae",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b918",x"3cad",x"374b",x"270a",x"3bfd",x"2877",x"3bce",x"3a59",x"b925",x"3cae",x"3749",x"257a",x"3bfd",x"28f4",x"3bcf",x"3a5e"),
(x"b90b",x"3cad",x"3722",x"2773",x"3bfe",x"22cf",x"3bd6",x"3a54",x"b911",x"3cae",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b92c",x"3cae",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60"),
(x"b907",x"3cae",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b90b",x"3cad",x"3722",x"2773",x"3bfe",x"22cf",x"3bd6",x"3a54",x"b92f",x"3cae",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62"),
(x"b8ff",x"3cae",x"3710",x"257a",x"3bff",x"1553",x"3bd9",x"3a4f",x"b907",x"3cae",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b931",x"3cae",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63"),
(x"b912",x"3c69",x"373c",x"1818",x"bbff",x"26c2",x"3a8e",x"3a57",x"b924",x"3c69",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b918",x"3c69",x"374b",x"2511",x"bbff",x"224c",x"3a91",x"3a59"),
(x"b90c",x"3c68",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55",x"b92b",x"3c69",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b912",x"3c69",x"373c",x"1818",x"bbff",x"26c2",x"3a8e",x"3a57"),
(x"b906",x"3c69",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53",x"b931",x"3c69",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63",x"b90c",x"3c68",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55"),
(x"b1fd",x"3c7a",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90",x"b1fd",x"3c7a",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b22d",x"3c78",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94"),
(x"b6fb",x"3c78",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08",x"b6fb",x"3c78",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6ef",x"3c74",x"3710",x"3b57",x"3658",x"0000",x"3a95",x"3a0c"),
(x"b63d",x"3c97",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5",x"b63d",x"3c97",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b62a",x"3c97",x"3710",x"2fbb",x"3bf1",x"0000",x"3aa1",x"39f9"),
(x"b1c1",x"3c7e",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89",x"b1c1",x"3c7e",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1fd",x"3c7a",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90"),
(x"b906",x"3c69",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53",x"b906",x"3c69",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b931",x"3c69",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63"),
(x"b721",x"3c7c",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00",x"b721",x"3c7c",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b6fb",x"3c78",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08"),
(x"b575",x"3ca7",x"3710",x"ba67",x"b8cb",x"068d",x"3aa1",x"3a26",x"b575",x"3ca7",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"3ca9",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28"),
(x"b1a1",x"3c7f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86",x"b1a1",x"3c7f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1c1",x"3c7e",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89"),
(x"b72e",x"3c7e",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd",x"b72e",x"3c7e",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b721",x"3c7c",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00"),
(x"b62a",x"3c97",x"3710",x"2fbb",x"3bf1",x"0000",x"3aa1",x"39f9",x"b62a",x"3c97",x"36da",x"303b",x"3bed",x"8000",x"3a97",x"39f9",x"b5ce",x"3c94",x"3710",x"2f26",x"3bf3",x"0000",x"3aa1",x"3a0b"),
(x"b161",x"3c80",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80",x"b161",x"3c80",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b1a1",x"3c7f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86"),
(x"b72d",x"3c80",x"3710",x"3778",x"bb13",x"0000",x"3a95",x"39fb",x"b72d",x"3c80",x"36da",x"3a45",x"b8f8",x"0000",x"3a8a",x"39fb",x"b72e",x"3c7e",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd"),
(x"b5ce",x"3c94",x"3710",x"2f26",x"3bf3",x"0000",x"3aa1",x"3a0b",x"b5ce",x"3c94",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5bd",x"3c95",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e"),
(x"b135",x"3c82",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b",x"b135",x"3c82",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b161",x"3c80",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80"),
(x"b721",x"3c81",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf",x"b721",x"3c81",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b72d",x"3c80",x"3710",x"3778",x"bb13",x"0000",x"3a87",x"3bb2"),
(x"b5bd",x"3c95",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e",x"b5bd",x"3c95",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5a1",x"3c99",x"3710",x"b72c",x"3b26",x"8000",x"3aa1",x"3a14"),
(x"b93a",x"3c96",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"3861",x"b93a",x"3c96",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"385a",x"b931",x"3c97",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b116",x"3c87",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77",x"b116",x"3c87",x"36da",x"3b51",x"b675",x"0000",x"3a6e",x"3b77",x"b135",x"3c82",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b"),
(x"b568",x"3c6a",x"3710",x"b810",x"bae4",x"868d",x"3a87",x"3b4e",x"b568",x"3c6a",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b575",x"3c6d",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52"),
(x"b5a1",x"3c99",x"3710",x"b72c",x"3b26",x"8000",x"3aa1",x"3a14",x"b5a1",x"3c99",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b581",x"3c9c",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a"),
(x"b669",x"3c81",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d",x"b669",x"3c81",x"36da",x"a65f",x"bbff",x"0000",x"3a7c",x"3b8d",x"b721",x"3c81",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf"),
(x"b581",x"3c9c",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a",x"b581",x"3c9c",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b568",x"3ca1",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21"),
(x"b8a3",x"3c6a",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d",x"b8a3",x"3c6a",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b906",x"3c69",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53"),
(x"b63d",x"3c7f",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84",x"b63d",x"3c7f",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b669",x"3c81",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d"),
(x"b568",x"3cad",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b",x"b568",x"3cad",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b558",x"3cae",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f"),
(x"b62a",x"3c7f",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81",x"b62a",x"3c7f",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b63d",x"3c7f",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84"),
(x"b558",x"3cae",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f",x"b558",x"3cae",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b544",x"3cae",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32"),
(x"b575",x"3c6d",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52",x"b575",x"3c6d",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3c70",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54"),
(x"b544",x"3cae",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32",x"b544",x"3cae",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b52b",x"3cb1",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37"),
(x"b5ce",x"3c82",x"3710",x"2ae9",x"bbfc",x"0000",x"3a87",x"3b6f",x"b5ce",x"3c82",x"36da",x"2f26",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b62a",x"3c7f",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81"),
(x"b52b",x"3cb1",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37",x"b52b",x"3cb1",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b50d",x"3cb2",x"3710",x"253f",x"3bff",x"8000",x"3aa1",x"3a3d"),
(x"b5bd",x"3c82",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c",x"b5bd",x"3c82",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5ce",x"3c82",x"3710",x"2ae9",x"bbfc",x"0000",x"3a87",x"3b6f"),
(x"b50d",x"3cb2",x"3710",x"253f",x"3bff",x"8000",x"3aa1",x"3a3d",x"b50d",x"3cb2",x"36da",x"324a",x"3bd8",x"0000",x"3a97",x"3a3d",x"b4f9",x"3caf",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41"),
(x"b5a1",x"3c7e",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66",x"b5a1",x"3c7e",x"36da",x"b72c",x"bb26",x"8000",x"3a7c",x"3b66",x"b5bd",x"3c82",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c"),
(x"b4f9",x"3caf",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41",x"b4f9",x"3caf",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f5",x"3cac",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44"),
(x"b581",x"3c7b",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f",x"b581",x"3c7b",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b5a1",x"3c7e",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66"),
(x"b4f5",x"3cac",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44",x"b4f5",x"3cac",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f2",x"3ca9",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47"),
(x"b931",x"3c97",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4",x"b931",x"3c97",x"36da",x"bbff",x"a4d0",x"0000",x"3a18",x"33f3",x"b931",x"3cae",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9"),
(x"b8ff",x"3cae",x"3710",x"257a",x"3bff",x"15bc",x"3bd9",x"3a4f",x"b8ff",x"3cae",x"36da",x"26a1",x"3bff",x"8000",x"3be3",x"3a4f",x"b8a3",x"3cac",x"3710",x"286d",x"3bfe",x"8000",x"3bd9",x"3a2b"),
(x"b568",x"3c75",x"3710",x"bb03",x"b7b2",x"868d",x"3a87",x"3b59",x"b568",x"3c75",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b581",x"3c7b",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f"),
(x"b4f2",x"3ca9",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47",x"b4f2",x"3ca9",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4da",x"3ca2",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d"),
(x"b8a3",x"3cac",x"3710",x"286d",x"3bfe",x"8000",x"3bd9",x"3a2b",x"b8a3",x"3cac",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b89e",x"3cac",x"3710",x"36f0",x"3b35",x"0000",x"3bd9",x"3a29"),
(x"b558",x"3c68",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b",x"b558",x"3c68",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b568",x"3c6a",x"3710",x"b810",x"bae4",x"868d",x"3a87",x"3b4e"),
(x"b4da",x"3ca2",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d",x"b4da",x"3ca2",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4d8",x"3c9f",x"3710",x"3be5",x"b11d",x"868d",x"3aa1",x"3a50"),
(x"b89e",x"3cac",x"3710",x"36f0",x"3b35",x"0000",x"3bd9",x"3a29",x"b89e",x"3cac",x"36da",x"380f",x"3ae4",x"068d",x"3be3",x"3a29",x"b88f",x"3ca7",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22"),
(x"b544",x"3c68",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47",x"b544",x"3c68",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b558",x"3c68",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b"),
(x"b4d8",x"3c9f",x"3710",x"3be5",x"b11d",x"868d",x"3aa1",x"3a50",x"b4d8",x"3c9f",x"36da",x"3af9",x"b7d8",x"8000",x"3a97",x"3a50",x"b4e1",x"3c9d",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52"),
(x"b88f",x"3ca7",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22",x"b88f",x"3ca7",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b87d",x"3ca2",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a"),
(x"b52b",x"3c65",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42",x"b52b",x"3c65",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b544",x"3c68",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47"),
(x"b4e1",x"3c9d",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52",x"b4e1",x"3c9d",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b51a",x"3c9a",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d"),
(x"b87d",x"3ca2",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a",x"b87d",x"3ca2",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b86e",x"3ca2",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14"),
(x"b50d",x"3c65",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c",x"b50d",x"3c65",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b52b",x"3c65",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42"),
(x"b51a",x"3c9a",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d",x"b51a",x"3c9a",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b528",x"3c99",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60"),
(x"b86e",x"3ca2",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14",x"b86e",x"3ca2",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b867",x"3ca4",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11"),
(x"b4f9",x"3c67",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38",x"b4f9",x"3c67",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b50d",x"3c65",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c"),
(x"b528",x"3c99",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60",x"b528",x"3c99",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b52c",x"3c98",x"3710",x"3bfc",x"ab6c",x"0000",x"3aa1",x"3a61"),
(x"b867",x"3ca4",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11",x"b867",x"3ca4",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b865",x"3ca7",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e"),
(x"b4f5",x"3c6a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35",x"b4f5",x"3c6a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f9",x"3c67",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38"),
(x"b52c",x"3c98",x"3710",x"3bfc",x"ab6c",x"0000",x"3a5f",x"39ec",x"b52c",x"3c98",x"36da",x"3b0d",x"378c",x"0000",x"3a54",x"39ec",x"b526",x"3c96",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee"),
(x"b865",x"3ca7",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e",x"b865",x"3ca7",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b85e",x"3cac",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09"),
(x"b4f2",x"3c6d",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33",x"b4f2",x"3c6d",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f5",x"3c6a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35"),
(x"b526",x"3c96",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee",x"b526",x"3c96",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b50c",x"3c95",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3"),
(x"b116",x"3c8f",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70",x"b116",x"3c8f",x"36da",x"3bdf",x"31b0",x"868d",x"3a6e",x"3b70",x"b116",x"3c87",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77"),
(x"b85e",x"3cac",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09",x"b85e",x"3cac",x"36da",x"b5f3",x"3b6d",x"8000",x"3be3",x"3a09",x"b84a",x"3cae",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01"),
(x"b4da",x"3c74",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c",x"b4da",x"3c74",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4f2",x"3c6d",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33"),
(x"b451",x"3c95",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16",x"b451",x"3c95",x"36da",x"a987",x"3bfe",x"8000",x"3a54",x"3a16",x"b441",x"3c96",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19"),
(x"b89e",x"3c6b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b",x"b89e",x"3c6b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b8a3",x"3c6a",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d"),
(x"b84a",x"3cae",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01",x"b84a",x"3cae",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b83a",x"3cab",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa"),
(x"b4d8",x"3c77",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a",x"b4d8",x"3c77",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4da",x"3c74",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c"),
(x"b50c",x"3c95",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3",x"b50c",x"3c95",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b451",x"3c95",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16"),
(x"b88f",x"3c6f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25",x"b88f",x"3c6f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b89e",x"3c6b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b"),
(x"b568",x"3ca1",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21",x"b568",x"3ca1",x"36da",x"bb03",x"37b2",x"068d",x"3a97",x"3a21",x"b569",x"3ca4",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23"),
(x"b4e1",x"3c79",x"3710",x"33d2",x"3bc1",x"0000",x"3a87",x"3b28",x"b4e1",x"3c79",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4d8",x"3c77",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a"),
(x"b441",x"3c96",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19",x"b441",x"3c96",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b40d",x"3c9e",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25"),
(x"b87d",x"3c74",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d",x"b87d",x"3c74",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b88f",x"3c6f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25"),
(x"b83a",x"3cab",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa",x"b83a",x"3cab",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b820",x"3c9e",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec"),
(x"b51a",x"3c7c",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d",x"b51a",x"3c7c",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b4e1",x"3c79",x"3710",x"33d2",x"3bc1",x"0000",x"3a87",x"3b28"),
(x"b40d",x"3c9e",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25",x"b40d",x"3c9e",x"36da",x"b8bf",x"3a70",x"8000",x"3a54",x"3a25",x"b407",x"3ca0",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27"),
(x"b86e",x"3c74",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17",x"b86e",x"3c74",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b87d",x"3c74",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d"),
(x"b569",x"3ca4",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23",x"b569",x"3ca4",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b575",x"3ca7",x"3710",x"ba67",x"b8cb",x"068d",x"3aa1",x"3a26"),
(x"b528",x"3c7e",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a",x"b528",x"3c7e",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b51a",x"3c7c",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d"),
(x"b407",x"3ca0",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27",x"b407",x"3ca0",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b409",x"3ca2",x"3710",x"bb1a",x"b75c",x"0000",x"3a5f",x"3a28"),
(x"b867",x"3c72",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14",x"b867",x"3c72",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b86e",x"3c74",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17"),
(x"b820",x"3c9e",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec",x"b820",x"3c9e",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b801",x"3c96",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de"),
(x"b52c",x"3c7f",x"3710",x"3b0d",x"b78c",x"0000",x"3a87",x"3b19",x"b52c",x"3c7f",x"36da",x"3bfc",x"2b6c",x"0000",x"3a7c",x"3b19",x"b528",x"3c7e",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a"),
(x"b409",x"3ca2",x"3710",x"bb1a",x"b75c",x"0000",x"3a5f",x"3a28",x"b409",x"3ca2",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b413",x"3ca5",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b"),
(x"b865",x"3c6f",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12",x"b865",x"3c6f",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b867",x"3c72",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14"),
(x"b801",x"3c96",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de",x"b801",x"3c96",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b7c0",x"3c94",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1"),
(x"b526",x"3c80",x"3710",x"33bc",x"bbc3",x"0000",x"3b06",x"3a0f",x"b526",x"3c80",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b52c",x"3c7f",x"3710",x"3b0d",x"b78c",x"0000",x"3b06",x"3a11"),
(x"b413",x"3ca5",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b",x"b413",x"3ca5",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"3ca7",x"3710",x"bb8c",x"354a",x"068d",x"3a5f",x"3a2d"),
(x"b85e",x"3c6a",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d",x"b85e",x"3c6a",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b865",x"3c6f",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12"),
(x"b7c0",x"3c94",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1",x"b7c0",x"3c94",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b794",x"3c96",x"3710",x"b358",x"3bc9",x"0000",x"3bd9",x"39c8"),
(x"b50c",x"3c81",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a",x"b50c",x"3c81",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b526",x"3c80",x"3710",x"33bc",x"bbc3",x"0000",x"3b06",x"3a0f"),
(x"b413",x"3ca7",x"3710",x"bb8c",x"354a",x"068d",x"3a5f",x"3a2d",x"b413",x"3ca7",x"36da",x"ba12",x"3935",x"8000",x"3a54",x"3a2d",x"b40b",x"3ca8",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e"),
(x"b84a",x"3c68",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05",x"b84a",x"3c68",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b85e",x"3c6a",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d"),
(x"b794",x"3c96",x"3710",x"b358",x"3bc9",x"0000",x"3bd9",x"39c8",x"b794",x"3c96",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b77a",x"3c99",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2"),
(x"b441",x"3c80",x"3710",x"b7a3",x"bb07",x"0000",x"3b06",x"39e4",x"b441",x"3c80",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b451",x"3c81",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7"),
(x"b40b",x"3ca8",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e",x"b40b",x"3ca8",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b3f4",x"3ca8",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32"),
(x"b83a",x"3c6b",x"3710",x"3953",x"b9f7",x"0000",x"3a85",x"39ff",x"b83a",x"3c6b",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b84a",x"3c68",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05"),
(x"b77a",x"3c99",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2",x"b77a",x"3c99",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b776",x"3c9c",x"3710",x"bbee",x"3037",x"0000",x"3bd9",x"39c0"),
(x"b451",x"3c81",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7",x"b451",x"3c81",x"36da",x"a0dd",x"bc00",x"0000",x"3afb",x"39e7",x"b50c",x"3c81",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a"),
(x"b3f4",x"3ca8",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32",x"b3f4",x"3ca8",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3d2",x"3ca7",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35"),
(x"b569",x"3c72",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57",x"b569",x"3c72",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b568",x"3c75",x"3710",x"bb03",x"b7b2",x"868d",x"3a87",x"3b59"),
(x"b776",x"3c9c",x"3710",x"bbee",x"3037",x"0000",x"3bd9",x"39c0",x"b776",x"3c9c",x"36da",x"bbce",x"b2fc",x"0000",x"3be3",x"39c0",x"b77b",x"3c9e",x"3710",x"b937",x"ba10",x"8000",x"3bd9",x"39be"),
(x"b40d",x"3c78",x"3710",x"b8bf",x"ba70",x"868d",x"3b06",x"39d8",x"b40d",x"3c78",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b441",x"3c80",x"3710",x"b7a3",x"bb07",x"0000",x"3b06",x"39e4"),
(x"b3d2",x"3ca7",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35",x"b3d2",x"3ca7",x"36da",x"abf9",x"3bfc",x"0000",x"3a54",x"3a35",x"b3a5",x"3ca8",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39"),
(x"b820",x"3c79",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1",x"b820",x"3c79",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b83a",x"3c6b",x"3710",x"3953",x"b9f7",x"0000",x"3a85",x"39ff"),
(x"b77b",x"3c9e",x"3710",x"b937",x"ba10",x"8000",x"3a87",x"3ac5",x"b77b",x"3c9e",x"36da",x"b853",x"baba",x"0000",x"3a7d",x"3ac5",x"b790",x"3ca0",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9"),
(x"b407",x"3c76",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6",x"b407",x"3c76",x"36da",x"bb61",x"b62a",x"0000",x"3afb",x"39d6",x"b40d",x"3c78",x"3710",x"b8bf",x"ba70",x"868d",x"3b06",x"39d8"),
(x"b3a5",x"3ca8",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39",x"b3a5",x"3ca8",x"36da",x"32b5",x"3bd2",x"068d",x"3a54",x"3a39",x"b368",x"3ca5",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40"),
(x"b575",x"3c70",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54",x"b575",x"3c70",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b569",x"3c72",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57"),
(x"b790",x"3ca0",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9",x"b790",x"3ca0",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b7a8",x"3ca1",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace"),
(x"b409",x"3c75",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5",x"b409",x"3c75",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b407",x"3c76",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6"),
(x"b368",x"3ca5",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40",x"b368",x"3ca5",x"36da",x"3912",x"3a2f",x"068d",x"3a54",x"3a40",x"b340",x"3c9f",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45"),
(x"b801",x"3c80",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4",x"b801",x"3c80",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b820",x"3c79",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1"),
(x"b7a8",x"3ca1",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace",x"b7a8",x"3ca1",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7bd",x"3ca4",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2"),
(x"b413",x"3c71",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2",x"b413",x"3c71",x"36da",x"bb08",x"37a1",x"8000",x"3afb",x"39d2",x"b409",x"3c75",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5"),
(x"b340",x"3c9f",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45",x"b340",x"3c9f",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b33a",x"3c9a",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49"),
(x"b7c0",x"3c82",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7",x"b7c0",x"3c82",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b801",x"3c80",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4"),
(x"b7bd",x"3ca4",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2",x"b7bd",x"3ca4",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7c7",x"3ca6",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5"),
(x"b931",x"3c69",x"3710",x"bbe9",x"26a1",x"309e",x"39f4",x"33ca",x"b931",x"3c69",x"36da",x"bbff",x"26b5",x"0000",x"39f5",x"33fa",x"b930",x"3c7f",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0"),
(x"b413",x"3c6f",x"3710",x"ba12",x"b935",x"0000",x"3b06",x"39d0",x"b413",x"3c6f",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"3c71",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2"),
(x"b33a",x"3c9a",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49",x"b33a",x"3c9a",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b351",x"3c95",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d"),
(x"b794",x"3c80",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf",x"b794",x"3c80",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b7c0",x"3c82",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7"),
(x"b7c7",x"3ca6",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5",x"b7c7",x"3ca6",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"3ca7",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6"),
(x"b40b",x"3c6e",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce",x"b40b",x"3c6e",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b413",x"3c6f",x"3710",x"ba12",x"b935",x"0000",x"3b06",x"39d0"),
(x"b351",x"3c95",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d",x"b351",x"3c95",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b34f",x"3c93",x"3710",x"3913",x"3a2f",x"0000",x"3a5f",x"3a4f"),
(x"b77a",x"3c7d",x"3710",x"b97c",x"b9d2",x"0000",x"3a85",x"39c9",x"b77a",x"3c7d",x"36da",x"b83f",x"bac7",x"0000",x"3a7b",x"39c9",x"b794",x"3c80",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf"),
(x"b7c7",x"3ca7",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6",x"b7c7",x"3ca7",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7a4",x"3cab",x"3710",x"b654",x"3b58",x"0000",x"3a87",x"3add"),
(x"b3f4",x"3c6e",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb",x"b3f4",x"3c6e",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b40b",x"3c6e",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce"),
(x"b34f",x"3c93",x"3710",x"3913",x"3a2f",x"0000",x"3a79",x"3b35",x"b34f",x"3c93",x"36da",x"3448",x"3bb5",x"0000",x"3a6e",x"3b35",x"b326",x"3c93",x"3710",x"a5e9",x"3bff",x"0000",x"3a79",x"3b39"),
(x"b776",x"3c7b",x"3710",x"bbce",x"32fb",x"0000",x"3a95",x"3a4d",x"b776",x"3c7b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b77a",x"3c7d",x"3710",x"b97c",x"b9d2",x"0000",x"3a95",x"3a50"),
(x"b7a4",x"3cab",x"3710",x"b654",x"3b58",x"0000",x"3a87",x"3add",x"b7a4",x"3cab",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b783",x"3cae",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4"),
(x"b3d2",x"3c70",x"3710",x"abf9",x"bbfc",x"0000",x"3b06",x"39c8",x"b3d2",x"3c70",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3f4",x"3c6e",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb"),
(x"b326",x"3c93",x"3710",x"a5e9",x"3bff",x"0000",x"3a79",x"3b39",x"b326",x"3c93",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b2d6",x"3c94",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41"),
(x"b77b",x"3c79",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c",x"b77b",x"3c79",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b776",x"3c7b",x"3710",x"bbce",x"32fb",x"0000",x"3a95",x"3a4d"),
(x"b783",x"3cae",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4",x"b783",x"3cae",x"36da",x"afa0",x"3bf1",x"8000",x"3a7d",x"3ae4",x"b73e",x"3caf",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1"),
(x"b3a5",x"3c6e",x"3710",x"32b5",x"bbd2",x"8000",x"3b06",x"39c3",x"b3a5",x"3c6e",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3d2",x"3c70",x"3710",x"abf9",x"bbfc",x"0000",x"3b06",x"39c8"),
(x"b2d6",x"3c94",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41",x"b2d6",x"3c94",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2aa",x"3c97",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46"),
(x"b790",x"3c76",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47",x"b790",x"3c76",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b77b",x"3c79",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c"),
(x"b73e",x"3caf",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1",x"b73e",x"3caf",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b705",x"3cac",x"3710",x"34b8",x"3ba4",x"0000",x"3a87",x"3afc"),
(x"b368",x"3c71",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd",x"b368",x"3c71",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b3a5",x"3c6e",x"3710",x"32b5",x"bbd2",x"8000",x"3b06",x"39c3"),
(x"b2aa",x"3c97",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46",x"b2aa",x"3c97",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b261",x"3c9c",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e"),
(x"b7a8",x"3c75",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43",x"b7a8",x"3c75",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b790",x"3c76",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47"),
(x"b705",x"3cac",x"3710",x"34b8",x"3ba4",x"0000",x"3a87",x"3afc",x"b705",x"3cac",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b6f1",x"3ca8",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01"),
(x"b340",x"3c77",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7",x"b340",x"3c77",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b368",x"3c71",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd"),
(x"b261",x"3c9c",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e",x"b261",x"3c9c",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b22d",x"3c9e",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53"),
(x"b7bd",x"3c73",x"3710",x"b821",x"3ada",x"0000",x"3a95",x"3a3e",x"b7bd",x"3c73",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7a8",x"3c75",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43"),
(x"b6f1",x"3ca8",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01",x"b6f1",x"3ca8",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6ef",x"3ca2",x"3710",x"3be9",x"b0b7",x"868d",x"3a87",x"3b05"),
(x"b33a",x"3c7c",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3",x"b33a",x"3c7c",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b340",x"3c77",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7"),
(x"b22d",x"3c9e",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53",x"b22d",x"3c9e",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b1fd",x"3c9d",x"3710",x"35da",x"3b72",x"8000",x"3a79",x"3b57"),
(x"b7c7",x"3c71",x"3710",x"bb43",x"36b4",x"0000",x"3a95",x"3a3c",x"b7c7",x"3c71",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7bd",x"3c73",x"3710",x"b821",x"3ada",x"0000",x"3a95",x"3a3e"),
(x"b6ef",x"3ca2",x"3710",x"3be9",x"b0b7",x"868d",x"3a87",x"3b05",x"b6ef",x"3ca2",x"36da",x"3b57",x"b658",x"8000",x"3a7d",x"3b05",x"b6fb",x"3c9f",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08"),
(x"b351",x"3c81",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af",x"b351",x"3c81",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b33a",x"3c7c",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3"),
(x"b1fd",x"3c9d",x"3710",x"35da",x"3b72",x"8000",x"3a79",x"3b57",x"b1fd",x"3c9d",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1c1",x"3c98",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e"),
(x"b7c7",x"3c6f",x"3710",x"b744",x"bb20",x"0000",x"3a95",x"3a3b",x"b7c7",x"3c6f",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"3c71",x"3710",x"bb43",x"36b4",x"0000",x"3a95",x"3a3c"),
(x"b6fb",x"3c9f",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08",x"b6fb",x"3c9f",x"36da",x"37ed",x"baf2",x"068d",x"3a7d",x"3b08",x"b721",x"3c9a",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10"),
(x"b34f",x"3c83",x"3710",x"3448",x"bbb5",x"0000",x"3b06",x"39ae",x"b34f",x"3c83",x"36da",x"3913",x"ba2f",x"8000",x"3afb",x"39ae",x"b351",x"3c81",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af"),
(x"b1c1",x"3c98",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e",x"b1c1",x"3c98",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1a1",x"3c97",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61"),
(x"b7a4",x"3c6c",x"3710",x"b64a",x"bb5a",x"0000",x"3a95",x"3a34",x"b7a4",x"3c6c",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7c7",x"3c6f",x"3710",x"b744",x"bb20",x"0000",x"3a95",x"3a3b"),
(x"b721",x"3c9a",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10",x"b721",x"3c9a",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b72e",x"3c98",x"3710",x"39a7",x"b9a8",x"0000",x"3a87",x"3b13"),
(x"b326",x"3c83",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae",x"b326",x"3c83",x"36da",x"a5e9",x"bbff",x"0000",x"3a6e",x"3bae",x"b34f",x"3c83",x"3710",x"3448",x"bbb5",x"0000",x"3a79",x"3bb2"),
(x"b1a1",x"3c97",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61",x"b1a1",x"3c97",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b161",x"3c96",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67"),
(x"b783",x"3c68",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d",x"b783",x"3c68",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b7a4",x"3c6c",x"3710",x"b64a",x"bb5a",x"0000",x"3a95",x"3a34"),
(x"b72e",x"3c98",x"3710",x"39a7",x"b9a8",x"0000",x"3aa1",x"39c6",x"b72e",x"3c98",x"36da",x"3b4f",x"b67e",x"0000",x"3a97",x"39c6",x"b72d",x"3c96",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8"),
(x"b2d6",x"3c82",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6",x"b2d6",x"3c82",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b326",x"3c83",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae"),
(x"b161",x"3c96",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67",x"b161",x"3c96",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b135",x"3c94",x"3710",x"3822",x"3ad9",x"868d",x"3a79",x"3b6c"),
(x"b73e",x"3c67",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20",x"b73e",x"3c67",x"36da",x"27ae",x"bbff",x"8000",x"3a8a",x"3a20",x"b783",x"3c68",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d"),
(x"b72d",x"3c96",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8",x"b72d",x"3c96",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b721",x"3c95",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca"),
(x"b2aa",x"3c7f",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2",x"b2aa",x"3c7f",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2d6",x"3c82",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6"),
(x"b135",x"3c94",x"3710",x"3822",x"3ad9",x"868d",x"3a79",x"3b6c",x"b135",x"3c94",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b116",x"3c8f",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70"),
(x"b705",x"3c6a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15",x"b705",x"3c6a",x"36da",x"34b8",x"bba4",x"8000",x"3a8a",x"3a15",x"b73e",x"3c67",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20"),
(x"b575",x"3ca9",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28",x"b575",x"3ca9",x"36da",x"bab5",x"385c",x"8a8d",x"3a97",x"3a28",x"b568",x"3cad",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b"),
(x"b938",x"3c81",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b938",x"3c81",x"36da",x"bbfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"b93a",x"3c96",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3be8",x"39da"),
(x"b261",x"3c7a",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a",x"b261",x"3c7a",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b2aa",x"3c7f",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2"),
(x"b931",x"3cae",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63",x"b931",x"3cae",x"36da",x"23ae",x"3bff",x"0000",x"3be3",x"3a63",x"b8ff",x"3cae",x"3710",x"257a",x"3bff",x"1553",x"3bd9",x"3a4f"),
(x"b6f1",x"3c6f",x"3710",x"3b73",x"b5d3",x"8000",x"3a95",x"3a10",x"b6f1",x"3c6f",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b705",x"3c6a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15"),
(x"b721",x"3c95",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca",x"b721",x"3c95",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b669",x"3c96",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed"),
(x"b22d",x"3c78",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94",x"b22d",x"3c78",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b261",x"3c7a",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a"),
(x"b6ef",x"3c74",x"3710",x"3b57",x"3658",x"0000",x"3a95",x"3a0c",x"b6ef",x"3c74",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6f1",x"3c6f",x"3710",x"3b73",x"b5d3",x"8000",x"3a95",x"3a10"),
(x"b669",x"3c96",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed",x"b669",x"3c96",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b63d",x"3c97",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5"),
(x"b930",x"3c7f",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c",x"b930",x"3c7f",x"36da",x"b67a",x"bb50",x"0000",x"3bc0",x"3984",x"b938",x"3c81",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a"),
(x"a165",x"39b8",x"36eb",x"bbf4",x"2d6d",x"ac2d",x"3929",x"3212",x"a379",x"39c2",x"36eb",x"bba3",x"b453",x"2fdf",x"392c",x"31f8",x"a1bd",x"39b8",x"3715",x"bbf4",x"2da3",x"2b3e",x"3920",x"31fe"),
(x"a271",x"39c2",x"3718",x"bbb8",x"b22d",x"31b0",x"3921",x"31e9",x"a379",x"39c2",x"36eb",x"bba3",x"b453",x"2fdf",x"392c",x"31f8",x"a303",x"39d2",x"3715",x"bbda",x"2e4f",x"312f",x"3924",x"31c9"),
(x"a303",x"39d2",x"3715",x"bbda",x"2e4f",x"312f",x"3924",x"31c9",x"a3d0",x"39d2",x"36eb",x"bb7a",x"3531",x"30a8",x"392e",x"31d7",x"a0f3",x"39e1",x"3714",x"ba0a",x"3915",x"3126",x"3926",x"31a6"),
(x"a0f3",x"39e1",x"3714",x"ba0a",x"3915",x"3126",x"3926",x"31a6",x"a133",x"39e5",x"36eb",x"b8c7",x"3a49",x"310c",x"3931",x"31aa",x"96c5",x"39e9",x"3714",x"b236",x"3bc0",x"30e0",x"3927",x"317f"),
(x"96c5",x"39e9",x"3714",x"b236",x"3bc0",x"30e0",x"3927",x"317f",x"9725",x"39ec",x"36eb",x"a3ae",x"3bec",x"3065",x"3932",x"3182",x"21e6",x"39e6",x"3714",x"335f",x"3baf",x"30fd",x"3928",x"3145"),
(x"21e6",x"39e6",x"3714",x"335f",x"3baf",x"30fd",x"3928",x"3145",x"22b9",x"39e9",x"36eb",x"36e0",x"3b1c",x"3118",x"3933",x"3141",x"24a4",x"39db",x"3715",x"3a37",x"38de",x"311d",x"3928",x"311f"),
(x"24a4",x"39db",x"3715",x"3a37",x"38de",x"311d",x"3928",x"311f",x"2505",x"39db",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3932",x"3119",x"252e",x"39cc",x"3715",x"3bf2",x"2495",x"2f43",x"3926",x"30fd"),
(x"256c",x"39cc",x"36eb",x"3bf7",x"2138",x"2dcf",x"3931",x"30f7",x"250e",x"39be",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"3930",x"30d9",x"252e",x"39cc",x"3715",x"3bf2",x"2495",x"2f43",x"3926",x"30fd"),
(x"250e",x"39be",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"3930",x"30d9",x"2470",x"39b4",x"36eb",x"3bfd",x"212b",x"29e6",x"392f",x"30c2",x"24bc",x"39be",x"3715",x"3b87",x"b537",x"2d81",x"3925",x"30e0"),
(x"24de",x"3981",x"3717",x"3be8",x"30a2",x"2973",x"391f",x"305e",x"250d",x"3981",x"36eb",x"3b9b",x"34d2",x"2ca7",x"392a",x"3055",x"25c0",x"397d",x"3714",x"3b74",x"35a7",x"2d5e",x"391f",x"304d"),
(x"20e0",x"39b7",x"3718",x"bbf1",x"95bc",x"2fb4",x"38d7",x"30e3",x"2066",x"39b7",x"36eb",x"bbf7",x"9e8d",x"2dbc",x"38cc",x"30e5",x"20c8",x"39c0",x"3716",x"bbb5",x"33c6",x"2f0a",x"38d7",x"30f8"),
(x"2116",x"397d",x"3718",x"ba6d",x"3838",x"3468",x"38d7",x"3067",x"2029",x"3983",x"36eb",x"ba79",x"3840",x"3401",x"38cb",x"3076",x"20e0",x"39b7",x"3718",x"bbf1",x"95bc",x"2fb4",x"38d7",x"30e3"),
(x"a4d5",x"3969",x"3715",x"b3c8",x"bbc2",x"236c",x"390e",x"32a2",x"a50e",x"3969",x"36eb",x"b409",x"bbbc",x"27db",x"3918",x"32b5",x"a4b5",x"397f",x"3715",x"bbb4",x"33e8",x"2ed7",x"3913",x"3278"),
(x"25ec",x"397f",x"36eb",x"3b76",x"3593",x"2dee",x"3929",x"3046",x"262b",x"3969",x"36eb",x"36d0",x"bb39",x"2ab1",x"3927",x"3019",x"25c0",x"397d",x"3714",x"3b74",x"35a7",x"2d5e",x"391f",x"304d"),
(x"993e",x"39b7",x"3716",x"3bce",x"b2bb",x"2b41",x"38d9",x"31ad",x"9909",x"39bf",x"3715",x"3b88",x"3531",x"2dc2",x"38d8",x"319c",x"9651",x"39b8",x"36eb",x"3bd3",x"b208",x"2da6",x"38ce",x"31ae"),
(x"9db7",x"39ca",x"3717",x"3bd6",x"323b",x"2a8a",x"38d9",x"3181",x"9caa",x"39c8",x"36ee",x"3b20",x"3725",x"2d51",x"38ce",x"3187",x"9909",x"39bf",x"3715",x"3b88",x"3531",x"2dc2",x"38d8",x"319c"),
(x"9cfd",x"39d2",x"3716",x"3aa5",x"b86c",x"2baa",x"38d8",x"316e",x"9cff",x"39d0",x"36ee",x"3b1d",x"b747",x"2911",x"38ce",x"3174",x"9db7",x"39ca",x"3717",x"3bd6",x"323b",x"2a8a",x"38d9",x"3181"),
(x"21f4",x"39d0",x"3714",x"bb20",x"b711",x"2eb1",x"38d7",x"311c",x"216b",x"39cf",x"36ee",x"ba3f",x"b8f6",x"2c87",x"38ce",x"3120",x"1f52",x"39d7",x"3715",x"b67e",x"bb4e",x"2839",x"38d7",x"3137"),
(x"9651",x"39b8",x"36eb",x"3bd3",x"b208",x"2da6",x"38ce",x"31ae",x"9fcf",x"3985",x"36eb",x"3be6",x"2cac",x"3077",x"38d0",x"321f",x"993e",x"39b7",x"3716",x"3bce",x"b2bb",x"2b41",x"38d9",x"31ad"),
(x"25f4",x"396a",x"3714",x"273e",x"ad9b",x"3bf7",x"3976",x"3263",x"24de",x"3981",x"3717",x"2984",x"a0c2",x"3bfd",x"3974",x"327f",x"25c0",x"397d",x"3714",x"33e6",x"2587",x"3bc0",x"3976",x"327a"),
(x"a4b5",x"397f",x"3715",x"b3f3",x"1d38",x"3bbf",x"395e",x"327d",x"a3f1",x"3980",x"3718",x"a6a1",x"97c8",x"3bff",x"3960",x"327e",x"a4d5",x"3969",x"3715",x"a081",x"ad9e",x"3bf8",x"395e",x"3263"),
(x"a271",x"39c2",x"3718",x"28fa",x"a4f7",x"3bfe",x"3962",x"32cc",x"9909",x"39bf",x"3715",x"28d3",x"a80e",x"3bfd",x"3968",x"32c8",x"a1bd",x"39b8",x"3715",x"a1ae",x"23fc",x"3bff",x"3963",x"32c0"),
(x"a303",x"39d2",x"3715",x"9ea7",x"2bd8",x"3bfc",x"3961",x"32de",x"9db7",x"39ca",x"3717",x"250b",x"281b",x"3bfe",x"3966",x"32d5",x"a271",x"39c2",x"3718",x"28fa",x"a4f7",x"3bfe",x"3962",x"32cc"),
(x"a0f3",x"39e1",x"3714",x"263f",x"27c1",x"3bfe",x"3963",x"32f0",x"9cfd",x"39d2",x"3716",x"252b",x"2c98",x"3bfa",x"3966",x"32df",x"a303",x"39d2",x"3715",x"9ea7",x"2bd8",x"3bfc",x"3961",x"32de"),
(x"96c5",x"39e9",x"3714",x"a194",x"a0d0",x"3bff",x"3968",x"32f9",x"94d9",x"39d7",x"3713",x"1818",x"9cd0",x"3c00",x"3968",x"32e4",x"a0f3",x"39e1",x"3714",x"263f",x"27c1",x"3bfe",x"3963",x"32f0"),
(x"21e6",x"39e6",x"3714",x"1dd6",x"247a",x"3bff",x"3970",x"32f6",x"1f52",x"39d7",x"3715",x"9cd0",x"191e",x"3c00",x"396d",x"32e6",x"96c5",x"39e9",x"3714",x"a194",x"a0d0",x"3bff",x"3968",x"32f9"),
(x"24a4",x"39db",x"3715",x"a793",x"184d",x"3bff",x"3973",x"32e9",x"21f4",x"39d0",x"3714",x"9dbc",x"252b",x"3bff",x"3970",x"32dc",x"21e6",x"39e6",x"3714",x"1dd6",x"247a",x"3bff",x"3970",x"32f6"),
(x"2211",x"39c9",x"3716",x"2338",x"267a",x"3bff",x"3970",x"32d4",x"21f4",x"39d0",x"3714",x"9dbc",x"252b",x"3bff",x"3970",x"32dc",x"252e",x"39cc",x"3715",x"9818",x"26bb",x"3bff",x"3975",x"32d7"),
(x"20c8",x"39c0",x"3716",x"24b5",x"2b17",x"3bfc",x"396e",x"32ca",x"2211",x"39c9",x"3716",x"2338",x"267a",x"3bff",x"3970",x"32d4",x"24bc",x"39be",x"3715",x"264c",x"29dc",x"3bfd",x"3974",x"32c7"),
(x"2464",x"39b5",x"3717",x"27d5",x"236c",x"3bfe",x"3973",x"32bc",x"20e0",x"39b7",x"3718",x"2793",x"2439",x"3bfe",x"396e",x"32be",x"24bc",x"39be",x"3715",x"264c",x"29dc",x"3bfd",x"3974",x"32c7"),
(x"2464",x"39b5",x"3717",x"27d5",x"236c",x"3bfe",x"3973",x"32bc",x"24de",x"3981",x"3717",x"2984",x"a0c2",x"3bfd",x"3974",x"327f",x"20e0",x"39b7",x"3718",x"2793",x"2439",x"3bfe",x"396e",x"32be"),
(x"2211",x"39c9",x"3716",x"bb9f",x"34a8",x"2d68",x"38d7",x"310e",x"219d",x"39c9",x"36ee",x"bb83",x"3534",x"2f10",x"38cd",x"3111",x"21f4",x"39d0",x"3714",x"bb20",x"b711",x"2eb1",x"38d7",x"311c"),
(x"a3f1",x"3980",x"3718",x"bba4",x"33dc",x"313d",x"3913",x"326a",x"a46c",x"3981",x"36eb",x"bbaa",x"3475",x"2c25",x"391d",x"327f",x"a1bd",x"39b8",x"3715",x"bbf4",x"2da3",x"2b3e",x"3920",x"31fe"),
(x"a4fc",x"3981",x"36eb",x"bbc6",x"328d",x"2f71",x"391c",x"3288",x"a46c",x"3981",x"36eb",x"bbaa",x"3475",x"2c25",x"391d",x"327f",x"a4b5",x"397f",x"3715",x"bbb4",x"33e8",x"2ed7",x"3913",x"3278"),
(x"25f4",x"396a",x"3714",x"273e",x"ad9b",x"3bf7",x"3976",x"3263",x"2116",x"397d",x"3718",x"23ae",x"ac2f",x"3bfb",x"396f",x"327a",x"24de",x"3981",x"3717",x"2984",x"a0c2",x"3bfd",x"3974",x"327f"),
(x"a069",x"397e",x"3718",x"a24c",x"a379",x"3bff",x"3964",x"327c",x"2116",x"397d",x"3718",x"23ae",x"ac2f",x"3bfb",x"396f",x"327a",x"a4d5",x"3969",x"3715",x"a081",x"ad9e",x"3bf8",x"395e",x"3263"),
(x"a3f1",x"3980",x"3718",x"a6a1",x"97c8",x"3bff",x"3960",x"327e",x"a069",x"397e",x"3718",x"a24c",x"a379",x"3bff",x"3964",x"327c",x"a4d5",x"3969",x"3715",x"a081",x"ad9e",x"3bf8",x"395e",x"3263"),
(x"9cfd",x"39d2",x"3716",x"3aa5",x"b86c",x"2baa",x"38d8",x"316e",x"94d9",x"39d7",x"3713",x"33d9",x"bbc1",x"a386",x"38d7",x"315c",x"9cff",x"39d0",x"36ee",x"3b1d",x"b747",x"2911",x"38ce",x"3174"),
(x"2464",x"39b5",x"3717",x"3bff",x"2481",x"2487",x"3924",x"30cb",x"2470",x"39b4",x"36eb",x"3bfd",x"212b",x"29e6",x"392f",x"30c2",x"24de",x"3981",x"3717",x"3be8",x"30a2",x"2973",x"391f",x"305e"),
(x"1f52",x"39d7",x"3715",x"b67e",x"bb4e",x"2839",x"38d7",x"3137",x"1f13",x"39d8",x"36ee",x"b233",x"bbd8",x"a538",x"38ce",x"3139",x"94d9",x"39d7",x"3713",x"33d9",x"bbc1",x"a386",x"38d7",x"315c"),
(x"9fcf",x"3985",x"36eb",x"3be6",x"2cac",x"3077",x"38d0",x"321f",x"2029",x"3983",x"36eb",x"ba79",x"3840",x"3401",x"38cb",x"3261",x"a069",x"397e",x"3718",x"398b",x"396b",x"33db",x"38db",x"3229"),
(x"262b",x"3969",x"36eb",x"36d0",x"bb39",x"2ab1",x"3927",x"3019",x"a50e",x"3969",x"36eb",x"b409",x"bbbc",x"27db",x"3918",x"2ec7",x"25f4",x"396a",x"3714",x"2f03",x"bbf3",x"23ef",x"391d",x"3024"),
(x"2211",x"39c9",x"3716",x"bb9f",x"34a8",x"2d68",x"38d7",x"310e",x"20c8",x"39c0",x"3716",x"bbb5",x"33c6",x"2f0a",x"38d7",x"30f8",x"219d",x"39c9",x"36ee",x"bb83",x"3534",x"2f10",x"38cd",x"3111"),
(x"9df1",x"3b85",x"3715",x"2d56",x"20d0",x"3bf8",x"3b50",x"3b10",x"91f4",x"3ba1",x"3716",x"30f9",x"a8b2",x"3be5",x"3b4b",x"3b05",x"20f7",x"3b90",x"370e",x"2fd2",x"2717",x"3bef",x"3b44",x"3b0d"),
(x"9df1",x"3b85",x"3715",x"bbc5",x"2b9a",x"3358",x"397d",x"302d",x"a03c",x"3b86",x"36eb",x"bb99",x"3315",x"330d",x"3982",x"302f",x"91f4",x"3ba1",x"3716",x"badd",x"375a",x"334d",x"397d",x"300e"),
(x"9a85",x"3b15",x"3713",x"ada1",x"2f15",x"3beb",x"3b52",x"3b41",x"8010",x"3b06",x"3714",x"ac39",x"29a5",x"3bf9",x"3b50",x"3b47",x"9d28",x"3b16",x"3712",x"aa69",x"287e",x"3bfc",x"3b54",x"3b40"),
(x"a273",x"3b06",x"3712",x"aa73",x"2a97",x"3bfa",x"3b5a",x"3b47",x"a34c",x"3b12",x"3711",x"a481",x"2546",x"3bff",x"3b5b",x"3b42",x"9ff6",x"3b1a",x"3711",x"a994",x"2977",x"3bfc",x"3b56",x"3b3e"),
(x"9ff6",x"3b1a",x"3711",x"a994",x"2977",x"3bfc",x"3b56",x"3b3e",x"9d28",x"3b16",x"3712",x"aa69",x"287e",x"3bfc",x"3b54",x"3b40",x"a273",x"3b06",x"3712",x"aa73",x"2a97",x"3bfa",x"3b5a",x"3b47"),
(x"9e8d",x"3aff",x"3716",x"af15",x"329c",x"3bc7",x"3b55",x"3b4a",x"9c36",x"3afd",x"3718",x"ae36",x"a153",x"3bf6",x"3b53",x"3b4b",x"a17b",x"3afb",x"3711",x"afec",x"ac2c",x"3beb",x"3b59",x"3b4b"),
(x"9c14",x"3ad5",x"370f",x"2b8a",x"30ae",x"3be6",x"3b54",x"3b5c",x"a035",x"3acc",x"3713",x"ae9c",x"3366",x"3bbd",x"3b58",x"3b60",x"9c56",x"3adb",x"370e",x"26d5",x"25c2",x"3bfe",x"3b54",x"3b5a"),
(x"a425",x"3ad8",x"370f",x"acd8",x"a71d",x"3bf9",x"3b5e",x"3b5a",x"9f72",x"3ae4",x"3713",x"a538",x"ac7a",x"3bfa",x"3b57",x"3b56",x"a289",x"3acf",x"370f",x"9df0",x"a631",x"3bff",x"3b5c",x"3b5e"),
(x"a425",x"3ad8",x"370f",x"acd8",x"a71d",x"3bf9",x"3b5e",x"3b5a",x"a407",x"3aeb",x"370f",x"aec5",x"1a24",x"3bf4",x"3b5d",x"3b52",x"9f72",x"3ae4",x"3713",x"a538",x"ac7a",x"3bfa",x"3b57",x"3b56"),
(x"a17b",x"3afb",x"3711",x"afec",x"ac2c",x"3beb",x"3b59",x"3b4b",x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f",x"9d1a",x"3aec",x"3710",x"ac5b",x"b0a5",x"3be5",x"3b55",x"3b52"),
(x"1d4c",x"3a9f",x"3717",x"97c8",x"9f79",x"3c00",x"3b4c",x"3b73",x"1e77",x"3a8d",x"3715",x"a6c2",x"ac65",x"3bfa",x"3b4b",x"3b7b",x"19fe",x"3a9c",x"3717",x"aff2",x"aa7a",x"3bed",x"3b4e",x"3b74"),
(x"a2cb",x"3a9a",x"3714",x"1553",x"ab62",x"3bfc",x"3b5b",x"3b75",x"a38f",x"3aa2",x"3712",x"b163",x"a345",x"3be2",x"3b5c",x"3b72",x"a13d",x"3aae",x"3716",x"acd8",x"a7e2",x"3bf9",x"3b58",x"3b6d"),
(x"a13d",x"3aae",x"3716",x"acd8",x"a7e2",x"3bf9",x"3b58",x"3b6d",x"9e62",x"3aad",x"3716",x"2818",x"ad02",x"3bf8",x"3b55",x"3b6d",x"a2cb",x"3a9a",x"3714",x"1553",x"ab62",x"3bfc",x"3b5b",x"3b75"),
(x"987a",x"3aa6",x"3714",x"a4f7",x"ada9",x"3bf7",x"3b52",x"3b70",x"9d1e",x"3a94",x"3711",x"240b",x"ad5c",x"3bf8",x"3b54",x"3b78",x"9e62",x"3aad",x"3716",x"2818",x"ad02",x"3bf8",x"3b55",x"3b6d"),
(x"0e53",x"3aa0",x"3714",x"b036",x"a73e",x"3bed",x"3b50",x"3b73",x"19fe",x"3a9c",x"3717",x"aff2",x"aa7a",x"3bed",x"3b4e",x"3b74",x"9a71",x"3a91",x"3711",x"b27d",x"175f",x"3bd5",x"3b53",x"3b79"),
(x"a16d",x"3a60",x"3711",x"b115",x"27d5",x"3be4",x"3b59",x"3b8d",x"9ae8",x"3a82",x"3712",x"b146",x"2c91",x"3bde",x"3b53",x"3b7f",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c"),
(x"1e3f",x"3a60",x"3715",x"28bc",x"afda",x"3bef",x"3b4c",x"3b8e",x"1f1f",x"3a6b",x"3718",x"2138",x"ae95",x"3bf4",x"3b4b",x"3b89",x"21e0",x"3a69",x"3719",x"a90e",x"af00",x"3bf2",x"3b47",x"3b8a"),
(x"1e3f",x"3a60",x"3715",x"28bc",x"afda",x"3bef",x"3b4c",x"3b8e",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c",x"1f1f",x"3a6b",x"3718",x"2138",x"ae95",x"3bf4",x"3b4b",x"3b89"),
(x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"1e5a",x"3a6d",x"3718",x"2b4f",x"2525",x"3bfc",x"3b4c",x"3b89",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c"),
(x"20ca",x"3a73",x"3715",x"2d65",x"ac5a",x"3bf3",x"3b49",x"3b86",x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"2288",x"3a7e",x"3718",x"2cf2",x"191e",x"3bf9",x"3b46",x"3b81"),
(x"2257",x"3a89",x"3712",x"3541",x"30b9",x"3b76",x"3b46",x"3b7c",x"22dc",x"3a86",x"3712",x"359c",x"336a",x"3b42",x"3b46",x"3b7e",x"2091",x"3a89",x"3717",x"2d2d",x"2ecb",x"3bed",x"3b49",x"3b7d"),
(x"2091",x"3a89",x"3717",x"2d2d",x"2ecb",x"3bed",x"3b49",x"3b7d",x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"1f4b",x"3a8a",x"3716",x"b009",x"2da6",x"3be7",x"3b4b",x"3b7c"),
(x"1e77",x"3a8d",x"3715",x"a6c2",x"ac65",x"3bfa",x"3b4b",x"3b7b",x"1f4b",x"3a8a",x"3716",x"b009",x"2da6",x"3be7",x"3b4b",x"3b7c",x"990c",x"3a8d",x"3712",x"af67",x"a981",x"3bf0",x"3b52",x"3b7b"),
(x"1f29",x"3a92",x"3714",x"a57a",x"ae8a",x"3bf4",x"3b4b",x"3b79",x"1e77",x"3a8d",x"3715",x"a6c2",x"ac65",x"3bfa",x"3b4b",x"3b7b",x"1d4c",x"3a9f",x"3717",x"97c8",x"9f79",x"3c00",x"3b4c",x"3b73"),
(x"2147",x"3a9a",x"3718",x"ac00",x"2911",x"3bfa",x"3b48",x"3b75",x"20ef",x"3aa9",x"3715",x"a51e",x"2d06",x"3bf9",x"3b49",x"3b6f",x"2442",x"3ab2",x"3714",x"175f",x"2c2c",x"3bfb",x"3b43",x"3b6b"),
(x"2442",x"3ab2",x"3714",x"175f",x"2c2c",x"3bfb",x"3b43",x"3b6b",x"2308",x"3ab8",x"3714",x"2dba",x"2266",x"3bf7",x"3b45",x"3b69",x"24cc",x"3acb",x"3712",x"3106",x"273e",x"3be5",x"3b41",x"3b61"),
(x"24cc",x"3acb",x"3712",x"3106",x"273e",x"3be5",x"3b41",x"3b61",x"2365",x"3ace",x"3715",x"3468",x"247a",x"3bb0",x"3b45",x"3b60",x"243c",x"3ae3",x"3710",x"3550",x"2e33",x"3b81",x"3b43",x"3b57"),
(x"243c",x"3ae3",x"3710",x"3550",x"2e33",x"3b81",x"3b43",x"3b57",x"22bc",x"3adf",x"3717",x"3273",x"2f43",x"3bc8",x"3b46",x"3b59",x"21ba",x"3af2",x"3712",x"2b5c",x"2345",x"3bfc",x"3b47",x"3b50"),
(x"21ba",x"3af2",x"3712",x"2b5c",x"2345",x"3bfc",x"3b47",x"3b50",x"1f35",x"3aed",x"3711",x"ae24",x"2a2e",x"3bf4",x"3b4b",x"3b52",x"1a19",x"3aef",x"3712",x"2dd2",x"b04b",x"3be4",x"3b4e",x"3b51"),
(x"9588",x"3b01",x"3716",x"a553",x"32c7",x"3bd1",x"3b51",x"3b49",x"08f2",x"3afe",x"3716",x"2f4d",x"aa5f",x"3bf0",x"3b50",x"3b4b",x"9c36",x"3afd",x"3718",x"ae36",x"a153",x"3bf6",x"3b53",x"3b4b"),
(x"9588",x"3b01",x"3716",x"a553",x"32c7",x"3bd1",x"3b51",x"3b49",x"9c36",x"3afd",x"3718",x"ae36",x"a153",x"3bf6",x"3b53",x"3b4b",x"9e8d",x"3aff",x"3716",x"af15",x"329c",x"3bc7",x"3b55",x"3b4a"),
(x"8010",x"3b06",x"3714",x"ac39",x"29a5",x"3bf9",x"3b50",x"3b47",x"9a85",x"3b15",x"3713",x"ada1",x"2f15",x"3beb",x"3b52",x"3b41",x"1f40",x"3b15",x"3717",x"b0e7",x"3057",x"3bd4",x"3b4a",x"3b41"),
(x"1f40",x"3b15",x"3717",x"b0e7",x"3057",x"3bd4",x"3b4a",x"3b41",x"1820",x"3b1f",x"370f",x"aedc",x"2cd0",x"3bee",x"3b4e",x"3b3d",x"221f",x"3b30",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3b45",x"3b36"),
(x"221f",x"3b30",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3b45",x"3b36",x"1d56",x"3b33",x"3716",x"aadf",x"a6b5",x"3bfc",x"3b4b",x"3b34",x"2273",x"3b4b",x"3717",x"abf6",x"25ae",x"3bfb",x"3b44",x"3b2a"),
(x"2273",x"3b4b",x"3717",x"abf6",x"25ae",x"3bfb",x"3b44",x"3b2a",x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c",x"2386",x"3b62",x"370f",x"36c9",x"2fac",x"3b2e",x"3b41",x"3b21"),
(x"2243",x"3b6c",x"3713",x"2f9d",x"b907",x"3a25",x"3b43",x"3b1c",x"2312",x"3b69",x"370d",x"3809",x"2e09",x"3add",x"3b41",x"3b1e",x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c"),
(x"20f7",x"3b90",x"370e",x"2fd2",x"2717",x"3bef",x"3b44",x"3b0d",x"21a5",x"3b7a",x"3712",x"29f0",x"2b1d",x"3bfa",x"3b43",x"3b16",x"9df1",x"3b85",x"3715",x"2d56",x"20d0",x"3bf8",x"3b50",x"3b10"),
(x"9cbb",x"3b6c",x"3715",x"bb81",x"b440",x"330f",x"397c",x"3048",x"1882",x"3b48",x"370e",x"bb5f",x"b5f1",x"2f4d",x"397b",x"306f",x"9f02",x"3b6a",x"36eb",x"bb89",x"b473",x"31fc",x"3981",x"304c"),
(x"a122",x"3a3e",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3bd9",x"396c",x"a167",x"3a20",x"36eb",x"3bf5",x"2e59",x"2467",x"3bd2",x"396c",x"a175",x"3a2c",x"3710",x"3bfd",x"a997",x"a0a8",x"3bd5",x"3971"),
(x"8dee",x"3a63",x"36eb",x"b46a",x"bb91",x"316a",x"3be4",x"396c",x"a122",x"3a3e",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3bd9",x"396c",x"9c3a",x"3a58",x"3714",x"3b1c",x"b754",x"223f",x"3be1",x"3971"),
(x"a167",x"3a20",x"36eb",x"3bf5",x"2e59",x"2467",x"3bd2",x"396c",x"a051",x"3a11",x"36eb",x"3ab1",x"3862",x"21e3",x"3bcd",x"396c",x"a099",x"3a14",x"3712",x"3b76",x"35c5",x"204d",x"3bce",x"3971"),
(x"a051",x"3a11",x"36eb",x"3ab1",x"3862",x"21e3",x"3bcd",x"396c",x"9b3f",x"3a09",x"36eb",x"37e1",x"3af5",x"269a",x"3bca",x"396c",x"9ecc",x"3a0d",x"3714",x"395a",x"39f1",x"2025",x"3bcc",x"3971"),
(x"9b3f",x"3a09",x"36eb",x"37e1",x"3af5",x"269a",x"3bca",x"396c",x"197e",x"3a06",x"36eb",x"303c",x"3beb",x"299b",x"3bc7",x"396c",x"9aa8",x"3a08",x"3714",x"35bf",x"3b76",x"27db",x"3bca",x"3971"),
(x"197e",x"3a06",x"36eb",x"303c",x"3beb",x"299b",x"3bc7",x"396c",x"20a0",x"3a08",x"36eb",x"b868",x"3aab",x"296a",x"3bc3",x"396c",x"1a1e",x"3a04",x"3715",x"a836",x"3bfd",x"294f",x"3bc6",x"3972"),
(x"20b2",x"3a07",x"3716",x"b86f",x"3aa7",x"2604",x"3bc3",x"3972",x"20a0",x"3a08",x"36eb",x"b868",x"3aab",x"296a",x"3bc3",x"396c",x"2335",x"3a14",x"3714",x"bb01",x"37b5",x"2839",x"3bbf",x"3971"),
(x"2300",x"3a14",x"36eb",x"baf3",x"37df",x"2b38",x"3bbf",x"396c",x"23d0",x"3a1e",x"36eb",x"bbf9",x"2d11",x"2511",x"3bbc",x"396c",x"2335",x"3a14",x"3714",x"bb01",x"37b5",x"2839",x"3bbf",x"3971"),
(x"23d0",x"3a1e",x"36eb",x"bbf9",x"2d11",x"2511",x"3bbc",x"396c",x"2300",x"3a28",x"36eb",x"b90c",x"ba34",x"2532",x"3bba",x"396c",x"23d3",x"3a1f",x"3714",x"bbe6",x"b10f",x"9bfc",x"3bbc",x"3971"),
(x"22d3",x"3a28",x"3715",x"b928",x"ba1d",x"1553",x"3b62",x"39e9",x"2300",x"3a28",x"36eb",x"b90c",x"ba34",x"2532",x"3b61",x"39ee",x"20d5",x"3a29",x"3714",x"2fe4",x"bbee",x"28fd",x"3b64",x"39e9"),
(x"20d5",x"3a29",x"3714",x"2fe4",x"bbee",x"28fd",x"3b64",x"39e9",x"20b2",x"3a28",x"36eb",x"35dd",x"bb6d",x"2be9",x"3b64",x"39ee",x"1e4f",x"3a25",x"3711",x"364f",x"bb52",x"2d1b",x"3b66",x"39ea"),
(x"865b",x"3a3e",x"36eb",x"b9db",x"396c",x"2c1a",x"3b71",x"39ef",x"13e1",x"3a42",x"36eb",x"bbf6",x"2a70",x"2d61",x"3b72",x"39ef",x"3d81",x"3a3e",x"3711",x"ba7a",x"38b0",x"283c",x"3b70",x"39ea"),
(x"1e4f",x"3a25",x"3711",x"364f",x"bb52",x"2d1b",x"3b66",x"39ea",x"1ead",x"3a23",x"36eb",x"32b1",x"bbc8",x"2e54",x"3b66",x"39ef",x"14bb",x"3a24",x"3710",x"b416",x"bbad",x"2f8d",x"3b68",x"39eb"),
(x"998f",x"3ad4",x"36eb",x"3b7d",x"b521",x"3095",x"3966",x"312c",x"9f83",x"3ac9",x"36eb",x"35e4",x"bb4d",x"31a2",x"396a",x"3125",x"9c14",x"3ad5",x"370f",x"3a9c",x"b854",x"30fa",x"3965",x"311a"),
(x"9cbb",x"3b6c",x"3715",x"bb81",x"b440",x"330f",x"397c",x"3048",x"9f02",x"3b6a",x"36eb",x"bb89",x"b473",x"31fc",x"3981",x"304c",x"9df1",x"3b85",x"3715",x"bbc5",x"2b9a",x"3358",x"397d",x"302d"),
(x"2375",x"3a3d",x"3711",x"a8d9",x"a52b",x"3bfe",x"3b45",x"3b9e",x"983c",x"3a38",x"3710",x"a856",x"a9ab",x"3bfc",x"3b53",x"3b9f",x"1f0f",x"3a43",x"3718",x"ab65",x"b528",x"3b8e",x"3b4b",x"3b9a"),
(x"210e",x"3b6e",x"36eb",x"3be3",x"2ce8",x"30c3",x"397a",x"2f8e",x"20f8",x"3b6d",x"3716",x"38de",x"3a57",x"297d",x"3976",x"2fa6",x"20d5",x"3b70",x"3715",x"3bd7",x"b1f9",x"2c2a",x"3977",x"2fab"),
(x"21ba",x"3af2",x"3712",x"384e",x"3ab0",x"2ec7",x"3965",x"2e4d",x"2267",x"3af4",x"36eb",x"3958",x"39de",x"2fdf",x"396a",x"2e4c",x"243c",x"3ae3",x"3710",x"3b6a",x"35bb",x"2efe",x"3965",x"2e26"),
(x"0f13",x"3a23",x"36eb",x"b37e",x"bbba",x"2ef6",x"3b69",x"39ef",x"9889",x"3a27",x"36eb",x"baa4",x"b859",x"2fe5",x"3b6b",x"39ef",x"14bb",x"3a24",x"3710",x"b416",x"bbad",x"2f8d",x"3b68",x"39eb"),
(x"1e18",x"3a5b",x"36eb",x"3bfa",x"a0b5",x"2cb4",x"38fe",x"29d0",x"1e52",x"3a48",x"36eb",x"3be6",x"308e",x"2c41",x"3900",x"2982",x"1d4f",x"3a5b",x"3715",x"3bfa",x"a70a",x"2c48",x"38f9",x"29b5"),
(x"951c",x"3a29",x"3711",x"ba7f",x"b887",x"3089",x"3b6a",x"39eb",x"9889",x"3a27",x"36eb",x"baa4",x"b859",x"2fe5",x"3b6b",x"39ef",x"99ac",x"3a30",x"3710",x"bbcc",x"b227",x"2f2e",x"3b6c",x"39eb"),
(x"9aca",x"3ada",x"36eb",x"3b19",x"3744",x"2cf7",x"3965",x"312d",x"998f",x"3ad4",x"36eb",x"3b7d",x"b521",x"3095",x"3966",x"312c",x"9c56",x"3adb",x"370e",x"3b25",x"370d",x"2d68",x"3963",x"311c"),
(x"9c70",x"3a93",x"36eb",x"b7d8",x"baf6",x"2a35",x"398c",x"2af2",x"a30f",x"3a97",x"36eb",x"b6fe",x"bb25",x"2ea6",x"398d",x"2aa4",x"9d1e",x"3a94",x"3711",x"b4dc",x"bb97",x"2d61",x"3987",x"2ad2"),
(x"9a2a",x"3a3a",x"36eb",x"bb02",x"3776",x"2fc8",x"3b6f",x"39ef",x"865b",x"3a3e",x"36eb",x"b9db",x"396c",x"2c1a",x"3b71",x"39ef",x"983c",x"3a38",x"3710",x"bb2f",x"36d9",x"2e52",x"3b6e",x"39eb"),
(x"08f2",x"3afe",x"3716",x"37e9",x"3af1",x"2aa7",x"3963",x"2e82",x"8d14",x"3b00",x"36eb",x"3776",x"3b0b",x"2d41",x"3969",x"2e88",x"21ba",x"3af2",x"3712",x"384e",x"3ab0",x"2ec7",x"3965",x"2e4d"),
(x"1e3f",x"3a60",x"3715",x"395d",x"b9e3",x"2de3",x"38f9",x"29c9",x"1e6c",x"3a5e",x"36eb",x"39df",x"b964",x"2d28",x"38fe",x"29db",x"1d4f",x"3a5b",x"3715",x"3bfa",x"a70a",x"2c48",x"38f9",x"29b5"),
(x"9f72",x"3ae4",x"3713",x"3b5b",x"3634",x"2c03",x"3961",x"311c",x"9f02",x"3ae5",x"36eb",x"3ad3",x"3822",x"2c4d",x"3962",x"3131",x"9c56",x"3adb",x"370e",x"3b25",x"370d",x"2d68",x"3963",x"311c"),
(x"1d56",x"3b33",x"3716",x"bbff",x"20c2",x"2138",x"3978",x"3084",x"1d3a",x"3b33",x"36eb",x"bbfe",x"1ea7",x"2828",x"397e",x"308a",x"1882",x"3b48",x"370e",x"bb5f",x"b5f1",x"2f4d",x"397b",x"306f"),
(x"9427",x"3b01",x"36eb",x"3b23",x"b71c",x"2cde",x"3969",x"2e8c",x"8d14",x"3b00",x"36eb",x"3776",x"3b0b",x"2d41",x"3969",x"2e88",x"9588",x"3b01",x"3716",x"3bde",x"31b5",x"2825",x"3963",x"2e8b"),
(x"21e0",x"3a69",x"3719",x"39a6",x"b994",x"2fc6",x"38f8",x"2a02",x"22d4",x"3a69",x"36eb",x"39ed",x"b94b",x"2f45",x"38fd",x"2a25",x"1e3f",x"3a60",x"3715",x"395d",x"b9e3",x"2de3",x"38f9",x"29c9"),
(x"9acb",x"3a8c",x"36eb",x"bbf8",x"a379",x"2d44",x"38fb",x"1f47",x"9c70",x"3a93",x"36eb",x"b7d8",x"baf6",x"2a35",x"38fb",x"1e54",x"9a71",x"3a91",x"3711",x"bb12",x"b763",x"2ca3",x"38f6",x"1f45"),
(x"9f87",x"3ae7",x"3713",x"3b09",x"b791",x"2ab8",x"3960",x"311d",x"9f11",x"3ae7",x"36eb",x"39e9",x"b955",x"2e31",x"3961",x"3132",x"9f72",x"3ae4",x"3713",x"3b5b",x"3634",x"2c03",x"3961",x"311c"),
(x"173f",x"3b20",x"36eb",x"bab4",x"3859",x"2a66",x"397c",x"309f",x"1d3a",x"3b33",x"36eb",x"bbfe",x"1ea7",x"2828",x"397e",x"308a",x"1820",x"3b1f",x"370f",x"bad7",x"3821",x"29e6",x"3978",x"309b"),
(x"141e",x"3b05",x"36eb",x"397a",x"b9b6",x"309a",x"3964",x"2ee0",x"9427",x"3b01",x"36eb",x"3b23",x"b71c",x"2cde",x"3963",x"2eda",x"8010",x"3b06",x"3714",x"39e8",x"b951",x"2f27",x"3961",x"2f04"),
(x"2283",x"3a6d",x"36eb",x"32cb",x"3bc1",x"2fc5",x"38fc",x"2a36",x"22d4",x"3a69",x"36eb",x"39ed",x"b94b",x"2f45",x"38fd",x"2a25",x"21d8",x"3a6b",x"3719",x"3250",x"3bca",x"2f22",x"38f7",x"2a09"),
(x"9bea",x"3a84",x"36eb",x"bb57",x"3625",x"2e99",x"38fc",x"2028",x"9acb",x"3a8c",x"36eb",x"bbf8",x"a379",x"2d44",x"38fb",x"1f47",x"9ae8",x"3a82",x"3712",x"bb92",x"3509",x"2cb0",x"38f7",x"2098"),
(x"9096",x"3aef",x"36eb",x"3046",x"bbe8",x"2cb7",x"398d",x"27a9",x"9f11",x"3ae7",x"36eb",x"39e9",x"b955",x"2e31",x"398e",x"2729",x"9d1a",x"3aec",x"3710",x"3833",x"bac7",x"2d1d",x"3989",x"274a"),
(x"9a85",x"3b15",x"3713",x"b7c2",x"3af3",x"2e28",x"3977",x"30a9",x"9bdf",x"3b17",x"36eb",x"b73f",x"3b1a",x"2d3c",x"397c",x"30ae",x"1820",x"3b1f",x"370f",x"bad7",x"3821",x"29e6",x"3978",x"309b"),
(x"2078",x"3b14",x"36eb",x"3aff",x"b73c",x"3197",x"3968",x"2efa",x"141e",x"3b05",x"36eb",x"397a",x"b9b6",x"309a",x"3964",x"2ee0",x"1f40",x"3b15",x"3717",x"3a77",x"b889",x"310e",x"3965",x"2f1f"),
(x"1f1f",x"3a6b",x"3718",x"30c6",x"3be6",x"2ad9",x"38f6",x"2a29",x"1e72",x"3a6c",x"36eb",x"3b01",x"3745",x"3141",x"38fa",x"2a64",x"21d8",x"3a6b",x"3719",x"3250",x"3bca",x"2f22",x"38f7",x"2a09"),
(x"a25f",x"3a5e",x"36eb",x"bb99",x"345f",x"30d6",x"38ff",x"22bb",x"9bea",x"3a84",x"36eb",x"bb57",x"3625",x"2e99",x"38fc",x"2028",x"a16d",x"3a60",x"3711",x"bb70",x"3585",x"3014",x"38fa",x"22e8"),
(x"1ecc",x"3aeb",x"36eb",x"b74a",x"bb15",x"2de4",x"398d",x"2814",x"9096",x"3aef",x"36eb",x"3046",x"bbe8",x"2cb7",x"398d",x"27a9",x"1a19",x"3aef",x"3712",x"b2e8",x"bbcb",x"2c10",x"3988",x"27d6"),
(x"9d97",x"3b18",x"36eb",x"38ae",x"3a73",x"2d49",x"397c",x"30b1",x"9bdf",x"3b17",x"36eb",x"b73f",x"3b1a",x"2d3c",x"397c",x"30ae",x"9d28",x"3b16",x"3712",x"3721",x"3b24",x"2bf9",x"3977",x"30ae"),
(x"231e",x"3b30",x"36eb",x"3bbf",x"b113",x"322d",x"396e",x"2f22",x"2078",x"3b14",x"36eb",x"3aff",x"b73c",x"3197",x"3968",x"2efa",x"221f",x"3b30",x"3713",x"3bc6",x"b1be",x"30de",x"396b",x"2f42"),
(x"a397",x"3a41",x"36eb",x"bbe6",x"2c77",x"308c",x"3901",x"2450",x"a25f",x"3a5e",x"36eb",x"bb99",x"345f",x"30d6",x"38ff",x"22bb",x"a2e9",x"3a41",x"3711",x"bbe4",x"2d1d",x"308c",x"38fc",x"2478"),
(x"22bc",x"3adf",x"3717",x"bb6f",x"b5e4",x"261e",x"3987",x"285d",x"2284",x"3adf",x"36eb",x"baaf",x"b860",x"2a70",x"398d",x"285d",x"1f35",x"3aed",x"3711",x"b934",x"ba0d",x"2c16",x"3988",x"280f"),
(x"9f8c",x"3b1c",x"36eb",x"2e28",x"3be6",x"3005",x"397c",x"30b7",x"9d97",x"3b18",x"36eb",x"38ae",x"3a73",x"2d49",x"397c",x"30b1",x"9ff6",x"3b1a",x"3711",x"35dd",x"3b65",x"2eae",x"3977",x"30b5"),
(x"2273",x"3b4b",x"3717",x"3bf0",x"af0f",x"2aec",x"396f",x"2f6c",x"22be",x"3b4b",x"36eb",x"3bea",x"ae0a",x"2f10",x"3973",x"2f49",x"221f",x"3b30",x"3713",x"3bc6",x"b1be",x"30de",x"396b",x"2f42"),
(x"1e72",x"3a6c",x"36eb",x"3b01",x"3745",x"3141",x"3969",x"2cf7",x"1f1f",x"3a6b",x"3718",x"30c6",x"3be6",x"2ad9",x"3963",x"2cfe",x"1e5a",x"3a6d",x"3718",x"3af5",x"b7e1",x"2460",x"3963",x"2d03"),
(x"a2ee",x"3a1f",x"3714",x"bbec",x"ad02",x"2f4a",x"38fe",x"258f",x"a382",x"3a1e",x"36eb",x"bbe8",x"ad68",x"3010",x"3903",x"256b",x"a2e9",x"3a41",x"3711",x"bbe4",x"2d1d",x"308c",x"38fc",x"2478"),
(x"2365",x"3ace",x"3715",x"bbfe",x"2412",x"2867",x"3988",x"28a3",x"234c",x"3acf",x"36eb",x"bbfa",x"ac62",x"2617",x"398d",x"28a0",x"22bc",x"3adf",x"3717",x"bb6f",x"b5e4",x"261e",x"3987",x"285d"),
(x"a2ba",x"3b1c",x"36eb",x"b913",x"3a0d",x"310f",x"397b",x"30c4",x"9f8c",x"3b1c",x"36eb",x"2e28",x"3be6",x"3005",x"397c",x"30b7",x"a20d",x"3b19",x"3712",x"b5a6",x"3b63",x"30cc",x"3977",x"30bd"),
(x"2414",x"3b61",x"36eb",x"3be4",x"aadf",x"30ee",x"3977",x"2f68",x"22be",x"3b4b",x"36eb",x"3bea",x"ae0a",x"2f10",x"3973",x"2f49",x"2386",x"3b62",x"370f",x"3bdd",x"b0de",x"2e6c",x"3974",x"2f86"),
(x"2349",x"3a7d",x"36eb",x"3bbf",x"b333",x"2ed2",x"396a",x"2d27",x"21d1",x"3a75",x"36eb",x"3a0e",x"b929",x"2e76",x"3969",x"2d12",x"2288",x"3a7e",x"3718",x"3b13",x"b732",x"2fec",x"3964",x"2d2f"),
(x"a269",x"3a0c",x"36eb",x"bab2",x"b834",x"30cb",x"3904",x"2600",x"a382",x"3a1e",x"36eb",x"bbe8",x"ad68",x"3010",x"3903",x"256b",x"a1ea",x"3a0f",x"3712",x"bb45",x"b640",x"30a6",x"38ff",x"2610"),
(x"99ac",x"3a30",x"3710",x"bbcc",x"b227",x"2f2e",x"3b6c",x"39eb",x"9b9c",x"3a30",x"36eb",x"bbf4",x"9ef6",x"2ebb",x"3b6d",x"39ef",x"983c",x"3a38",x"3710",x"bb2f",x"36d9",x"2e52",x"3b6e",x"39eb"),
(x"2308",x"3ab8",x"3714",x"bb81",x"3558",x"2da6",x"3988",x"2900",x"22be",x"3aba",x"36eb",x"bbcf",x"32aa",x"2bc5",x"398d",x"28f8",x"2365",x"3ace",x"3715",x"bbfe",x"2412",x"2867",x"3988",x"28a3"),
(x"a3f7",x"3b12",x"36eb",x"bbe5",x"adbc",x"3036",x"397a",x"30ce",x"a2ba",x"3b1c",x"36eb",x"b913",x"3a0d",x"310f",x"397b",x"30c4",x"a34c",x"3b12",x"3711",x"bbb2",x"332f",x"30f4",x"3976",x"30c7"),
(x"23bf",x"3b6c",x"36eb",x"3af6",x"3714",x"32f0",x"3979",x"2f79",x"2414",x"3b61",x"36eb",x"3be4",x"aadf",x"30ee",x"3977",x"2f68",x"2312",x"3b69",x"370d",x"3b0d",x"370c",x"3169",x"3976",x"2f8f"),
(x"2324",x"3a89",x"36eb",x"3bbf",x"3370",x"2dad",x"396a",x"2d3f",x"2349",x"3a7d",x"36eb",x"3bbf",x"b333",x"2ed2",x"396a",x"2d27",x"22dc",x"3a86",x"3712",x"3bf0",x"2c20",x"2e95",x"3965",x"2d3f"),
(x"9dfd",x"39fc",x"36eb",x"b7cb",x"bae6",x"3068",x"3904",x"26ad",x"a269",x"3a0c",x"36eb",x"bab2",x"b834",x"30cb",x"3904",x"2600",x"9d7f",x"3a00",x"3715",x"b93c",x"b9e9",x"3110",x"38ff",x"26b7"),
(x"20ef",x"3aa9",x"3715",x"ba65",x"38c1",x"2d9c",x"3988",x"2949",x"207d",x"3aaa",x"36eb",x"bac2",x"3833",x"2e8a",x"398d",x"2945",x"2308",x"3ab8",x"3714",x"bb81",x"3558",x"2da6",x"3988",x"2900"),
(x"a2c3",x"3b03",x"36eb",x"b902",x"ba23",x"306a",x"3979",x"30dd",x"a3f7",x"3b12",x"36eb",x"bbe5",x"adbc",x"3036",x"397a",x"30ce",x"a273",x"3b06",x"3712",x"bae4",x"b7c3",x"30c9",x"3975",x"30d1"),
(x"2243",x"3b6c",x"3713",x"3451",x"3bac",x"2d81",x"3976",x"2f9b",x"226e",x"3b6e",x"36eb",x"3571",x"3b6d",x"30cc",x"397a",x"2f84",x"2312",x"3b69",x"370d",x"3b0d",x"370c",x"3169",x"3976",x"2f8f"),
(x"22c6",x"3a8b",x"36eb",x"2eda",x"3bea",x"2e47",x"396a",x"2d45",x"2324",x"3a89",x"36eb",x"3bbf",x"3370",x"2dad",x"396a",x"2d3f",x"2257",x"3a89",x"3712",x"3298",x"3bcc",x"2d84",x"3965",x"2d48"),
(x"17aa",x"39f8",x"36eb",x"96f6",x"bbf5",x"2e99",x"3905",x"2736",x"9dfd",x"39fc",x"36eb",x"b7cb",x"bae6",x"3068",x"3904",x"26ad",x"17a2",x"39fb",x"3715",x"9ef6",x"bbee",x"302a",x"38ff",x"273a"),
(x"1d4c",x"3a9f",x"3717",x"b939",x"3a0b",x"29e0",x"3988",x"2980",x"1ce6",x"3aa0",x"36eb",x"b9cd",x"3979",x"2caa",x"398d",x"297b",x"20ef",x"3aa9",x"3715",x"ba65",x"38c1",x"2d9c",x"3988",x"2949"),
(x"9ff8",x"3b01",x"36eb",x"b3f1",x"bbbc",x"2b5c",x"3977",x"30e7",x"a2c3",x"3b03",x"36eb",x"b902",x"ba23",x"306a",x"3979",x"30dd",x"a040",x"3b03",x"3713",x"b607",x"bb5e",x"2e4f",x"3973",x"30d9"),
(x"20f8",x"3b6d",x"3716",x"38de",x"3a57",x"297d",x"3976",x"2fa6",x"210e",x"3b6e",x"36eb",x"3be3",x"2ce8",x"30c3",x"397a",x"2f8e",x"2243",x"3b6c",x"3713",x"3451",x"3bac",x"2d81",x"3976",x"2f9b"),
(x"2091",x"3a89",x"3717",x"2a0a",x"3bfc",x"284d",x"3964",x"2d56",x"2058",x"3a8a",x"36eb",x"2c58",x"3bf7",x"2bc5",x"396a",x"2d59",x"2257",x"3a89",x"3712",x"3298",x"3bcc",x"2d84",x"3965",x"2d48"),
(x"210b",x"3a00",x"3713",x"382e",x"baba",x"306c",x"3900",x"27ca",x"20e4",x"39fc",x"36eb",x"366a",x"bb44",x"2f81",x"3905",x"27be",x"17a2",x"39fb",x"3715",x"9ef6",x"bbee",x"302a",x"38ff",x"273a"),
(x"19fe",x"3a9c",x"3717",x"2c95",x"3bf9",x"2918",x"3988",x"2997",x"1a1b",x"3a9d",x"36eb",x"35a5",x"3b74",x"2d53",x"398d",x"298f",x"1d4c",x"3a9f",x"3717",x"b939",x"3a0b",x"29e0",x"3988",x"2980"),
(x"9e8d",x"3aff",x"3716",x"bac7",x"383c",x"283f",x"3972",x"30dd",x"9efd",x"3aff",x"36eb",x"b94d",x"39f2",x"2dc5",x"3977",x"30e9",x"a040",x"3b03",x"3713",x"b607",x"bb5e",x"2e4f",x"3973",x"30d9"),
(x"1882",x"3b48",x"370e",x"b004",x"a71d",x"3bef",x"3b4d",x"3b2b",x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c",x"2273",x"3b4b",x"3717",x"abf6",x"25ae",x"3bfb",x"3b44",x"3b2a"),
(x"1f7b",x"3a8c",x"36eb",x"3b71",x"b58a",x"2fc3",x"396a",x"2d60",x"2058",x"3a8a",x"36eb",x"2c58",x"3bf7",x"2bc5",x"396a",x"2d59",x"1f4b",x"3a8a",x"3716",x"38f4",x"3a42",x"2c09",x"3964",x"2d5e"),
(x"2466",x"3a0c",x"3715",x"3ae0",x"b7cf",x"30d4",x"38ff",x"2836",x"24bd",x"3a0a",x"36eb",x"39f2",x"b938",x"30b5",x"3904",x"283d",x"210b",x"3a00",x"3713",x"382e",x"baba",x"306c",x"3900",x"27ca"),
(x"98cf",x"3aa9",x"36eb",x"3976",x"39cc",x"2dcc",x"398e",x"29d2",x"1a1b",x"3a9d",x"36eb",x"35a5",x"3b74",x"2d53",x"398d",x"298f",x"0e53",x"3aa0",x"3714",x"39a7",x"399e",x"2d1e",x"3988",x"29b0"),
(x"a282",x"3afc",x"36eb",x"b9ec",x"392b",x"31e4",x"3975",x"30f4",x"9efd",x"3aff",x"36eb",x"b94d",x"39f2",x"2dc5",x"3977",x"30e9",x"a17b",x"3afb",x"3711",x"b8c8",x"3a4e",x"30a8",x"3971",x"30e7"),
(x"1f7b",x"3a8c",x"36eb",x"3b71",x"b58a",x"2fc3",x"396a",x"2d60",x"1f4b",x"3a8a",x"3716",x"38f4",x"3a42",x"2c09",x"3964",x"2d5e",x"1e77",x"3a8d",x"3715",x"3ac1",x"b812",x"3146",x"3964",x"2d67"),
(x"253f",x"3a1e",x"3715",x"3bec",x"abe2",x"2fce",x"38ff",x"2887",x"2585",x"3a1d",x"36eb",x"3bc4",x"b27a",x"3012",x"3904",x"2891",x"2466",x"3a0c",x"3715",x"3ae0",x"b7cf",x"30d4",x"38ff",x"2836"),
(x"9e13",x"3aae",x"36eb",x"353f",x"3b87",x"2d28",x"398e",x"29f7",x"98cf",x"3aa9",x"36eb",x"3976",x"39cc",x"2dcc",x"398e",x"29d2",x"9e62",x"3aad",x"3716",x"37d5",x"3af0",x"2d8e",x"3989",x"29ff"),
(x"a471",x"3aeb",x"36eb",x"bbbc",x"3212",x"3175",x"3972",x"3105",x"a282",x"3afc",x"36eb",x"b9ec",x"392b",x"31e4",x"3975",x"30f4",x"a407",x"3aeb",x"370f",x"bb4b",x"35cc",x"3223",x"396f",x"30f8"),
(x"21ae",x"3b92",x"36eb",x"3ade",x"37ab",x"31d3",x"397f",x"2fd1",x"229f",x"3b7b",x"36eb",x"3bdb",x"1c67",x"320a",x"397c",x"2fa6",x"20f7",x"3b90",x"370e",x"3b7b",x"34a9",x"3270",x"397b",x"2fe0"),
(x"22bc",x"3a9c",x"36eb",x"3adb",x"b7e7",x"30ac",x"396a",x"2d88",x"1e77",x"3a8d",x"3715",x"3ac1",x"b812",x"3146",x"3964",x"2d67",x"2147",x"3a9a",x"3718",x"3ac6",x"b7dc",x"3286",x"3964",x"2d86"),
(x"24fc",x"3a2f",x"3717",x"3b55",x"35fd",x"307e",x"38fd",x"28cc",x"255d",x"3a30",x"36eb",x"3b6e",x"3575",x"309f",x"3903",x"28e0",x"253f",x"3a1e",x"3715",x"3bec",x"abe2",x"2fce",x"38ff",x"2887"),
(x"a16d",x"3a60",x"3711",x"b115",x"27d5",x"3be4",x"3b59",x"3b8d",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c",x"9c3a",x"3a58",x"3714",x"b05e",x"2194",x"3bec",x"3b54",x"3b91"),
(x"a172",x"3ab0",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"398e",x"2a20",x"9e13",x"3aae",x"36eb",x"353f",x"3b87",x"2d28",x"398e",x"29f7",x"a13d",x"3aae",x"3716",x"a345",x"3bf7",x"2dcc",x"3989",x"2a21"),
(x"a482",x"3ad7",x"36eb",x"bb61",x"b5a0",x"3119",x"396f",x"3114",x"a471",x"3aeb",x"36eb",x"bbbc",x"3212",x"3175",x"3972",x"3105",x"a425",x"3ad8",x"370f",x"bbd3",x"af46",x"3182",x"396c",x"3106"),
(x"2496",x"3ab2",x"36eb",x"3bba",x"b376",x"2f14",x"396a",x"2dbb",x"22bc",x"3a9c",x"36eb",x"3adb",x"b7e7",x"30ac",x"396a",x"2d88",x"2442",x"3ab2",x"3714",x"3b6b",x"b587",x"3095",x"3965",x"2dbe"),
(x"2409",x"3a40",x"36eb",x"3884",x"3a69",x"3249",x"3902",x"292c",x"255d",x"3a30",x"36eb",x"3b6e",x"3575",x"309f",x"3903",x"28e0",x"2375",x"3a3d",x"3711",x"38a4",x"3a69",x"309a",x"38fd",x"2913"),
(x"a38b",x"3aac",x"36eb",x"bacb",x"3812",x"3064",x"398e",x"2a48",x"a172",x"3ab0",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"398e",x"2a20",x"a2d9",x"3aab",x"3714",x"b976",x"39c0",x"3023",x"3989",x"2a41"),
(x"a2ad",x"3acb",x"36eb",x"b86e",x"ba87",x"313e",x"396c",x"311e",x"a482",x"3ad7",x"36eb",x"bb61",x"b5a0",x"3119",x"396f",x"3114",x"a289",x"3acf",x"370f",x"b891",x"ba73",x"30f5",x"396a",x"310e"),
(x"1a0c",x"3ba6",x"36eb",x"38a6",x"3a54",x"3207",x"3982",x"3001",x"21ae",x"3b92",x"36eb",x"3ade",x"37ab",x"31d3",x"397f",x"2fd1",x"1aac",x"3ba1",x"3712",x"38b5",x"3a3e",x"32bd",x"397d",x"3005"),
(x"250f",x"3acc",x"36eb",x"3bef",x"2d09",x"2e69",x"396a",x"2df2",x"2496",x"3ab2",x"36eb",x"3bba",x"b376",x"2f14",x"396a",x"2dbb",x"24cc",x"3acb",x"3712",x"3bf0",x"aa00",x"2f46",x"3965",x"2df3"),
(x"1f0f",x"3a43",x"3718",x"38ae",x"3a78",x"2b7c",x"38fb",x"294e",x"1fad",x"3a43",x"36eb",x"360d",x"3b5a",x"2ef3",x"3900",x"296f",x"2375",x"3a3d",x"3711",x"38a4",x"3a69",x"309a",x"38fd",x"2913"),
(x"a422",x"3aa1",x"36eb",x"bbcf",x"b174",x"303e",x"398e",x"2a77",x"a38b",x"3aac",x"36eb",x"bacb",x"3812",x"3064",x"398e",x"2a48",x"a38f",x"3aa2",x"3712",x"bbe0",x"2e5e",x"30a3",x"3989",x"2a66"),
(x"a035",x"3acc",x"3713",x"3583",x"bb63",x"3153",x"3967",x"3112",x"9f83",x"3ac9",x"36eb",x"35e4",x"bb4d",x"31a2",x"396a",x"3125",x"a289",x"3acf",x"370f",x"b891",x"ba73",x"30f5",x"396a",x"310e"),
(x"91f4",x"3ba1",x"3716",x"badd",x"375a",x"334d",x"397d",x"300e",x"980d",x"3ba6",x"36eb",x"b996",x"395f",x"33ec",x"3983",x"300b",x"1aac",x"3ba1",x"3712",x"38b5",x"3a3e",x"32bd",x"397d",x"3005"),
(x"2469",x"3ae4",x"36eb",x"3b75",x"35a2",x"2d46",x"396a",x"2e25",x"250f",x"3acc",x"36eb",x"3bef",x"2d09",x"2e69",x"396a",x"2df2",x"243c",x"3ae3",x"3710",x"3b6a",x"35bb",x"2efe",x"3965",x"2e26"),
(x"1d9c",x"3a48",x"3718",x"3be6",x"309f",x"2baa",x"38fa",x"2966",x"1e52",x"3a48",x"36eb",x"3be6",x"308e",x"2c41",x"3900",x"2982",x"1f0f",x"3a43",x"3718",x"38ae",x"3a78",x"2b7c",x"38fb",x"294e"),
(x"a30f",x"3a97",x"36eb",x"b6fe",x"bb25",x"2ea6",x"398d",x"2aa4",x"a422",x"3aa1",x"36eb",x"bbcf",x"b174",x"303e",x"398e",x"2a77",x"a2cb",x"3a9a",x"3714",x"b972",x"b9bb",x"30de",x"3988",x"2a88"),
(x"a175",x"3a2c",x"3710",x"2828",x"260a",x"3bfe",x"3b5a",x"3ba3",x"a140",x"3a1c",x"3714",x"2946",x"1ffc",x"3bfe",x"3b5a",x"3baa",x"a2ee",x"3a1f",x"3714",x"2eb0",x"28fa",x"3bf3",x"3b5c",x"3ba9"),
(x"a099",x"3a14",x"3712",x"2953",x"27b4",x"3bfd",x"3b59",x"3bae",x"9ecc",x"3a0d",x"3714",x"a8bf",x"2c22",x"3bfa",x"3b57",x"3bb0",x"a1ea",x"3a0f",x"3712",x"a587",x"209b",x"3bff",x"3b5b",x"3baf"),
(x"9aa8",x"3a08",x"3714",x"231d",x"2b5f",x"3bfc",x"3b55",x"3bb3",x"9d7f",x"3a00",x"3715",x"a0ea",x"2afd",x"3bfc",x"3b57",x"3bb6",x"9ecc",x"3a0d",x"3714",x"a8bf",x"2c22",x"3bfa",x"3b57",x"3bb0"),
(x"1a1e",x"3a04",x"3715",x"270a",x"a779",x"3bfe",x"3b50",x"3bb5",x"17a2",x"39fb",x"3715",x"27e2",x"29b2",x"3bfc",x"3b51",x"3bb9",x"9aa8",x"3a08",x"3714",x"231d",x"2b5f",x"3bfc",x"3b55",x"3bb3"),
(x"20b2",x"3a07",x"3716",x"24bc",x"aceb",x"3bf9",x"3b4b",x"3bb4",x"210b",x"3a00",x"3713",x"2b1d",x"aee4",x"3bf0",x"3b4a",x"3bb7",x"1a1e",x"3a04",x"3715",x"270a",x"a779",x"3bfe",x"3b50",x"3bb5"),
(x"2335",x"3a14",x"3714",x"a8e0",x"299e",x"3bfc",x"3b47",x"3baf",x"2466",x"3a0c",x"3715",x"a266",x"9d87",x"3bff",x"3b44",x"3bb2",x"20b2",x"3a07",x"3716",x"24bc",x"aceb",x"3bf9",x"3b4b",x"3bb4"),
(x"23d3",x"3a1f",x"3714",x"a538",x"a9ab",x"3bfd",x"3b45",x"3baa",x"253f",x"3a1e",x"3715",x"a891",x"a7ce",x"3bfd",x"3b41",x"3bab",x"2335",x"3a14",x"3714",x"a8e0",x"299e",x"3bfc",x"3b47",x"3baf"),
(x"23d3",x"3a1f",x"3714",x"a538",x"a9ab",x"3bfd",x"3b45",x"3baa",x"22d3",x"3a28",x"3715",x"ac67",x"28a5",x"3bf9",x"3b47",x"3ba6",x"253f",x"3a1e",x"3715",x"a891",x"a7ce",x"3bfd",x"3b41",x"3bab"),
(x"20d5",x"3a29",x"3714",x"aa45",x"2b10",x"3bfa",x"3b4a",x"3ba6",x"2375",x"3a3d",x"3711",x"a8d9",x"a52b",x"3bfe",x"3b45",x"3b9e",x"22d3",x"3a28",x"3715",x"ac67",x"28a5",x"3bf9",x"3b47",x"3ba6"),
(x"14bb",x"3a24",x"3710",x"a352",x"ae80",x"3bf5",x"3b51",x"3ba7",x"951c",x"3a29",x"3711",x"abef",x"a8a8",x"3bfa",x"3b52",x"3ba5",x"1e4f",x"3a25",x"3711",x"aa66",x"b31a",x"3bca",x"3b4d",x"3ba7"),
(x"1d9c",x"3a48",x"3718",x"b420",x"1418",x"3bba",x"3b4c",x"3b98",x"1f0f",x"3a43",x"3718",x"ab65",x"b528",x"3b8e",x"3b4b",x"3b9a",x"15a0",x"3a42",x"3713",x"b41f",x"ac3a",x"3bb6",x"3b50",x"3b9b"),
(x"16c6",x"3a4b",x"3714",x"ade0",x"a4c2",x"3bf6",x"3b50",x"3b97",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c",x"1d4f",x"3a5b",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3b4d",x"3b90"),
(x"951c",x"3a29",x"3711",x"abef",x"a8a8",x"3bfa",x"3b52",x"3ba5",x"983c",x"3a38",x"3710",x"a856",x"a9ab",x"3bfc",x"3b53",x"3b9f",x"20d5",x"3a29",x"3714",x"aa45",x"2b10",x"3bfa",x"3b4a",x"3ba6"),
(x"a3f1",x"3980",x"3718",x"a6a1",x"97c8",x"3bff",x"3960",x"327e",x"a1bd",x"39b8",x"3715",x"a1ae",x"23fc",x"3bff",x"3963",x"32c0",x"a069",x"397e",x"3718",x"a24c",x"a379",x"3bff",x"3964",x"327c"),
(x"1e3f",x"3a60",x"3715",x"28bc",x"afda",x"3bef",x"3b4c",x"3b8e",x"1d4f",x"3a5b",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3b4d",x"3b90",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c"),
(x"13e1",x"3a42",x"36eb",x"bbf6",x"2a70",x"2d61",x"3b72",x"39ef",x"8dee",x"3a63",x"36eb",x"b46a",x"bb91",x"316a",x"3b7b",x"39ee",x"16c6",x"3a4b",x"3714",x"bbf3",x"ae23",x"2b27",x"3b73",x"39ea"),
(x"20de",x"3798",x"3715",x"ad56",x"a0d0",x"3bf8",x"391b",x"38a5",x"1c89",x"3761",x"3716",x"b0f9",x"28b2",x"3be5",x"3914",x"3896",x"9e24",x"3783",x"370e",x"afd2",x"a717",x"3bef",x"390a",x"38a1"),
(x"20de",x"3798",x"3715",x"3bc5",x"ab9a",x"3358",x"3957",x"300b",x"2222",x"3797",x"36eb",x"3b99",x"b315",x"330d",x"395c",x"300e",x"1c89",x"3761",x"3716",x"3add",x"b75a",x"334d",x"3958",x"2fd9"),
(x"1f0d",x"383c",x"3713",x"2da1",x"af14",x"3beb",x"391e",x"38e5",x"1ba5",x"384b",x"3714",x"2c39",x"a9a5",x"3bf9",x"391a",x"38ee",x"2079",x"383b",x"3712",x"2a69",x"a87e",x"3bfc",x"3920",x"38e4"),
(x"242c",x"384b",x"3712",x"2a73",x"aa97",x"3bfa",x"3928",x"38ed",x"2498",x"383f",x"3711",x"2481",x"a54c",x"3bff",x"392a",x"38e7",x"21e0",x"3837",x"3711",x"2994",x"a977",x"3bfc",x"3922",x"38e2"),
(x"21e0",x"3837",x"3711",x"2994",x"a977",x"3bfc",x"3922",x"38e2",x"2079",x"383b",x"3712",x"2a69",x"a87e",x"3bfc",x"3920",x"38e4",x"242c",x"384b",x"3712",x"2a73",x"aa97",x"3bfa",x"3928",x"38ed"),
(x"212c",x"3852",x"3716",x"2f15",x"b29c",x"3bc7",x"3921",x"38f1",x"2000",x"3854",x"3718",x"2e36",x"2153",x"3bf6",x"391f",x"38f3",x"2360",x"3856",x"3711",x"2fec",x"2c2c",x"3beb",x"3926",x"38f4"),
(x"1fdf",x"387c",x"370f",x"ab8a",x"b0ae",x"3be6",x"3921",x"390a",x"221a",x"3885",x"3713",x"2e9c",x"b367",x"3bbd",x"3926",x"390f",x"2010",x"3876",x"370e",x"a6dc",x"a5c2",x"3bfe",x"3921",x"3907"),
(x"2517",x"3879",x"370f",x"2cd8",x"271d",x"3bf9",x"392e",x"3907",x"219e",x"386d",x"3713",x"2538",x"2c79",x"3bfa",x"3924",x"3901",x"2437",x"3883",x"370f",x"1df0",x"2631",x"3bff",x"392a",x"390d"),
(x"2517",x"3879",x"370f",x"2cd8",x"271d",x"3bf9",x"392e",x"3907",x"24fa",x"3866",x"370f",x"2ec5",x"9a24",x"3bf4",x"392d",x"38fd",x"219e",x"386d",x"3713",x"2538",x"2c79",x"3bfa",x"3924",x"3901"),
(x"2360",x"3856",x"3711",x"2fec",x"2c2c",x"3beb",x"3926",x"38f4",x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8",x"2072",x"3865",x"3710",x"2c5b",x"30a5",x"3be5",x"3921",x"38fd"),
(x"9607",x"38b2",x"3717",x"17c8",x"1f79",x"3c00",x"3915",x"3929",x"9959",x"38c4",x"3715",x"26c2",x"2c65",x"3bfa",x"3914",x"3933",x"125b",x"38b5",x"3717",x"2ff2",x"2a7a",x"3bed",x"3918",x"392b"),
(x"2458",x"38b7",x"3714",x"9553",x"2b62",x"3bfc",x"3929",x"392b",x"24ba",x"38af",x"3712",x"3163",x"2345",x"3be2",x"392b",x"3927",x"2323",x"38a3",x"3716",x"2cd8",x"27e2",x"3bf9",x"3926",x"3920"),
(x"2323",x"38a3",x"3716",x"2cd8",x"27e2",x"3bf9",x"3926",x"3920",x"2116",x"38a4",x"3716",x"a818",x"2d02",x"3bf8",x"3922",x"3921",x"2458",x"38b7",x"3714",x"9553",x"2b62",x"3bfc",x"3929",x"392b"),
(x"1e07",x"38ab",x"3714",x"24fd",x"2da9",x"3bf7",x"391d",x"3925",x"2074",x"38bd",x"3711",x"a412",x"2d5c",x"3bf8",x"3920",x"392f",x"2116",x"38a4",x"3716",x"a818",x"2d02",x"3bf8",x"3922",x"3921"),
(x"1acb",x"38b1",x"3714",x"3036",x"273e",x"3bed",x"391b",x"3928",x"125b",x"38b5",x"3717",x"2ff2",x"2a7a",x"3bed",x"3918",x"392b",x"1f03",x"38c0",x"3711",x"327d",x"975f",x"3bd5",x"391f",x"3931"),
(x"2353",x"38f1",x"3711",x"3115",x"a7d5",x"3be4",x"3927",x"394c",x"1f3f",x"38cf",x"3712",x"3146",x"ac91",x"3bde",x"391f",x"3939",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b"),
(x"98e9",x"38f1",x"3715",x"a8bf",x"2fda",x"3bef",x"3915",x"394d",x"9aa8",x"38e6",x"3718",x"a138",x"2e94",x"3bf4",x"3914",x"3947",x"9ff6",x"38e8",x"3719",x"290e",x"2efe",x"3bf2",x"390f",x"3948"),
(x"98e9",x"38f1",x"3715",x"a8bf",x"2fda",x"3bef",x"3915",x"394d",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b",x"9aa8",x"38e6",x"3718",x"a138",x"2e94",x"3bf4",x"3914",x"3947"),
(x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"9920",x"38e4",x"3718",x"ab4f",x"a52b",x"3bfc",x"3915",x"3946",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b"),
(x"9dca",x"38de",x"3715",x"ad65",x"2c5a",x"3bf3",x"3911",x"3942",x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"a0a3",x"38d3",x"3718",x"acf2",x"991e",x"3bf9",x"390d",x"393c"),
(x"a072",x"38c8",x"3712",x"b541",x"b0b9",x"3b76",x"390e",x"3935",x"a0f6",x"38cb",x"3712",x"b59c",x"b36a",x"3b42",x"390d",x"3937",x"9d58",x"38c8",x"3717",x"ad2f",x"aecb",x"3bed",x"3912",x"3935"),
(x"9d58",x"38c8",x"3717",x"ad2f",x"aecb",x"3bed",x"3912",x"3935",x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"9b02",x"38c7",x"3716",x"3009",x"ada6",x"3be7",x"3914",x"3935"),
(x"9959",x"38c4",x"3715",x"26c2",x"2c65",x"3bfa",x"3914",x"3933",x"9b02",x"38c7",x"3716",x"3009",x"ada6",x"3be7",x"3914",x"3935",x"1e50",x"38c4",x"3712",x"2f67",x"2981",x"3bf0",x"391e",x"3933"),
(x"9abe",x"38bf",x"3714",x"2581",x"2e8a",x"3bf4",x"3913",x"3930",x"9959",x"38c4",x"3715",x"26c2",x"2c65",x"3bfa",x"3914",x"3933",x"9607",x"38b2",x"3717",x"17c8",x"1f79",x"3c00",x"3915",x"3929"),
(x"9ec5",x"38b7",x"3718",x"2c00",x"a90e",x"3bfa",x"3910",x"392c",x"9e13",x"38a8",x"3715",x"251e",x"ad06",x"3bf9",x"3911",x"3924",x"a29f",x"389f",x"3714",x"975f",x"ac2c",x"3bfb",x"3909",x"391e"),
(x"a29f",x"389f",x"3714",x"975f",x"ac2c",x"3bfb",x"3909",x"391e",x"a123",x"3899",x"3714",x"adba",x"a266",x"3bf7",x"390c",x"391b",x"a3b3",x"3886",x"3712",x"b106",x"a738",x"3be5",x"3907",x"3910"),
(x"a3b3",x"3886",x"3712",x"b106",x"a738",x"3be5",x"3907",x"3910",x"a180",x"3883",x"3715",x"b468",x"a47a",x"3bb0",x"390c",x"390f",x"a294",x"386e",x"3710",x"b550",x"ae33",x"3b81",x"3909",x"3903"),
(x"a294",x"386e",x"3710",x"b550",x"ae33",x"3b81",x"3909",x"3903",x"a0d7",x"3872",x"3717",x"b273",x"af43",x"3bc8",x"390d",x"3905",x"9faa",x"385f",x"3712",x"ab5f",x"a345",x"3bfc",x"390f",x"38fa"),
(x"9faa",x"385f",x"3712",x"ab5f",x"a345",x"3bfc",x"390f",x"38fa",x"9ad5",x"3864",x"3711",x"2e23",x"aa31",x"3bf4",x"3914",x"38fd",x"11f0",x"3862",x"3712",x"add2",x"304b",x"3be4",x"3918",x"38fc"),
(x"1d2c",x"3850",x"3716",x"2553",x"b2c7",x"3bd1",x"391c",x"38f1",x"1b46",x"3853",x"3716",x"af4d",x"2a5f",x"3bf0",x"391a",x"38f3",x"2000",x"3854",x"3718",x"2e36",x"2153",x"3bf6",x"391f",x"38f3"),
(x"1d2c",x"3850",x"3716",x"2553",x"b2c7",x"3bd1",x"391c",x"38f1",x"2000",x"3854",x"3718",x"2e36",x"2153",x"3bf6",x"391f",x"38f3",x"212c",x"3852",x"3716",x"2f15",x"b29c",x"3bc7",x"3921",x"38f1"),
(x"1ba5",x"384b",x"3714",x"2c39",x"a9a5",x"3bf9",x"391a",x"38ee",x"1f0d",x"383c",x"3713",x"2da1",x"af14",x"3beb",x"391e",x"38e5",x"9aec",x"383c",x"3717",x"30e7",x"b058",x"3bd4",x"3912",x"38e6"),
(x"9aec",x"383c",x"3717",x"30e7",x"b058",x"3bd4",x"3912",x"38e6",x"16e7",x"3832",x"370f",x"2edc",x"acd0",x"3bee",x"3918",x"38e0",x"a039",x"3821",x"3713",x"29b8",x"26e9",x"3bfd",x"390c",x"38d7"),
(x"a039",x"3821",x"3713",x"29b8",x"26e9",x"3bfd",x"390c",x"38d7",x"9631",x"381e",x"3716",x"2adf",x"26b5",x"3bfc",x"3914",x"38d4",x"a08e",x"3806",x"3717",x"2bf6",x"a5ae",x"3bfb",x"390b",x"38c7"),
(x"a08e",x"3806",x"3717",x"2bf6",x"a5ae",x"3bfb",x"390b",x"38c7",x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4",x"a1a0",x"37df",x"370f",x"b6ca",x"afac",x"3b2e",x"3907",x"38bb"),
(x"a05e",x"37cb",x"3713",x"af9f",x"3907",x"3a26",x"3909",x"38b5",x"a12d",x"37d1",x"370d",x"b809",x"ae09",x"3add",x"3907",x"38b7",x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4"),
(x"9e24",x"3783",x"370e",x"afd2",x"a717",x"3bef",x"390a",x"38a1",x"9f80",x"37ae",x"3712",x"a9f0",x"ab1d",x"3bfa",x"390a",x"38ad",x"20de",x"3798",x"3715",x"ad56",x"a0d0",x"3bf8",x"391b",x"38a5"),
(x"2043",x"37cb",x"3715",x"3b81",x"3440",x"330f",x"3956",x"3026",x"1624",x"3809",x"370e",x"3b5f",x"35f1",x"2f4d",x"3955",x"304d",x"2166",x"37ce",x"36eb",x"3b89",x"3473",x"31fc",x"395b",x"302b"),
(x"2307",x"3913",x"36eb",x"bba1",x"34cc",x"1f45",x"395a",x"291b",x"234d",x"3931",x"36eb",x"bbf5",x"ae59",x"2467",x"395a",x"289e",x"235a",x"3925",x"3710",x"bbfd",x"2997",x"a0a8",x"3956",x"28cc"),
(x"1c29",x"38ee",x"36eb",x"346a",x"3b91",x"316a",x"395a",x"29cb",x"2307",x"3913",x"36eb",x"bba1",x"34cc",x"1f45",x"395a",x"291b",x"2002",x"38f9",x"3714",x"bb1c",x"3754",x"223f",x"3955",x"298e"),
(x"234d",x"3931",x"36eb",x"bbf5",x"ae59",x"2467",x"395a",x"289e",x"2237",x"3940",x"36eb",x"bab1",x"b862",x"21f0",x"395b",x"285c",x"227e",x"393d",x"3712",x"bb76",x"b5c5",x"204d",x"3956",x"2866"),
(x"2237",x"3940",x"36eb",x"bab1",x"b862",x"21f0",x"395b",x"285c",x"1f6a",x"3948",x"36eb",x"b7e1",x"baf5",x"269a",x"395b",x"2826",x"214b",x"3944",x"3714",x"b95a",x"b9f1",x"2025",x"3956",x"2845"),
(x"1f6a",x"3948",x"36eb",x"b7e1",x"baf5",x"269a",x"395b",x"2826",x"142d",x"394c",x"36eb",x"b03c",x"bbeb",x"299b",x"395b",x"27de",x"1f1f",x"3949",x"3714",x"b5bf",x"bb76",x"27db",x"3956",x"2820"),
(x"142d",x"394c",x"36eb",x"b03c",x"bbeb",x"299b",x"395b",x"27de",x"9d76",x"3949",x"36eb",x"3868",x"baab",x"296a",x"395b",x"2770",x"11db",x"394d",x"3715",x"2836",x"bbfd",x"294f",x"3956",x"27d1"),
(x"9d99",x"394a",x"3716",x"386f",x"baa7",x"2604",x"3956",x"2765",x"9d76",x"3949",x"36eb",x"3868",x"baab",x"296a",x"395b",x"2770",x"a14f",x"393d",x"3714",x"3b01",x"b7b5",x"2839",x"3956",x"26e0"),
(x"a11a",x"393d",x"36eb",x"3af3",x"b7df",x"2b38",x"395b",x"26eb",x"a1ea",x"3933",x"36eb",x"3bf9",x"ad11",x"2511",x"395b",x"2695",x"a14f",x"393d",x"3714",x"3b01",x"b7b5",x"2839",x"3956",x"26e0"),
(x"a1ea",x"3933",x"36eb",x"3bf9",x"ad11",x"2511",x"395b",x"2695",x"a11a",x"3929",x"36eb",x"390c",x"3a34",x"2532",x"395c",x"2642",x"a1ee",x"3932",x"3714",x"3be6",x"310f",x"9bfc",x"3956",x"267f"),
(x"a0ed",x"3929",x"3715",x"3928",x"3a1d",x"1553",x"3956",x"262a",x"a11a",x"3929",x"36eb",x"390c",x"3a34",x"2532",x"395c",x"2642",x"9ddf",x"3928",x"3714",x"afe4",x"3bee",x"28fd",x"3957",x"25e8"),
(x"9ddf",x"3928",x"3714",x"afe4",x"3bee",x"28fd",x"3957",x"25e8",x"9d99",x"3929",x"36eb",x"b5dd",x"3b6d",x"2be9",x"395c",x"25f5",x"9908",x"392c",x"3711",x"b64f",x"3b52",x"2d1b",x"3958",x"25a8"),
(x"1bc8",x"3913",x"36eb",x"39db",x"b96c",x"2c1a",x"395b",x"2439",x"199d",x"390f",x"36eb",x"3bf6",x"aa70",x"2d61",x"395b",x"2417",x"1b8a",x"3913",x"3711",x"3a7a",x"b8b0",x"283c",x"3957",x"245d"),
(x"9908",x"392c",x"3711",x"b64f",x"3b52",x"2d1b",x"3958",x"25a8",x"99c6",x"392e",x"36eb",x"b2b1",x"3bc8",x"2e54",x"395c",x"25b8",x"1937",x"392d",x"3710",x"3416",x"3bad",x"2f8d",x"3958",x"2552"),
(x"1e92",x"387d",x"36eb",x"bb7d",x"3521",x"3096",x"3b21",x"3a52",x"21a6",x"3888",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b24",x"3a53",x"1fdf",x"387c",x"370f",x"ba9b",x"3854",x"30fa",x"3b23",x"3a4e"),
(x"2043",x"37cb",x"3715",x"3b81",x"3440",x"330f",x"3956",x"3026",x"2166",x"37ce",x"36eb",x"3b89",x"3473",x"31fc",x"395b",x"302b",x"20de",x"3798",x"3715",x"3bc5",x"ab9a",x"3358",x"3957",x"300b"),
(x"a18f",x"3914",x"3711",x"28d9",x"252b",x"3bfe",x"390c",x"3962",x"1de8",x"3919",x"3710",x"2856",x"29ab",x"3bfc",x"391e",x"3963",x"9a89",x"390e",x"3718",x"2b65",x"3528",x"3b8f",x"3914",x"395d"),
(x"9e52",x"37c7",x"36eb",x"bbe3",x"ace8",x"30c3",x"3955",x"2f4a",x"9e25",x"37c9",x"3716",x"b8de",x"ba57",x"297d",x"3951",x"2f61",x"9de0",x"37c2",x"3715",x"bbd7",x"31f9",x"2c2a",x"3951",x"2f66"),
(x"9faa",x"385f",x"3712",x"b84e",x"bab0",x"2ec8",x"3972",x"28c9",x"a081",x"385d",x"36eb",x"b958",x"b9de",x"2fdf",x"3977",x"28c9",x"a294",x"386e",x"3710",x"bb6b",x"b5ba",x"2efe",x"3972",x"287b"),
(x"1ab2",x"392e",x"36eb",x"337e",x"3bba",x"2ef6",x"395c",x"2550",x"1e0f",x"392a",x"36eb",x"3aa4",x"3859",x"2fe5",x"395c",x"2513",x"1937",x"392d",x"3710",x"3416",x"3bad",x"2f8d",x"3958",x"2552"),
(x"989a",x"38f6",x"36eb",x"bbfa",x"20b5",x"2cb4",x"398c",x"2c6a",x"990f",x"3909",x"36eb",x"bbe6",x"b08e",x"2c41",x"398e",x"2c46",x"9613",x"38f6",x"3715",x"bbfa",x"2710",x"2c48",x"3988",x"2c55"),
(x"1d11",x"3928",x"3711",x"3a7e",x"3887",x"3089",x"3958",x"2517",x"1e0f",x"392a",x"36eb",x"3aa4",x"3859",x"2fe5",x"395c",x"2513",x"1ea1",x"3921",x"3710",x"3bcc",x"3227",x"2f2f",x"3958",x"24db"),
(x"1f2f",x"3877",x"36eb",x"bb19",x"b744",x"2cf7",x"3b1f",x"3a51",x"1e92",x"387d",x"36eb",x"bb7d",x"3521",x"3096",x"3b21",x"3a52",x"2010",x"3876",x"370e",x"bb25",x"b70d",x"2d6a",x"3b22",x"3a4d"),
(x"201d",x"38be",x"36eb",x"37d8",x"3af6",x"2a35",x"3997",x"27b6",x"247a",x"38ba",x"36eb",x"36fe",x"3b25",x"2ea4",x"3997",x"2711",x"2074",x"38bd",x"3711",x"34dc",x"3b97",x"2d60",x"3993",x"27ac"),
(x"1edf",x"3917",x"36eb",x"3b02",x"b777",x"2fc8",x"395c",x"2477",x"1bc8",x"3913",x"36eb",x"39db",x"b96c",x"2c1a",x"395b",x"2439",x"1de8",x"3919",x"3710",x"3b2f",x"b6d9",x"2e52",x"3957",x"2492"),
(x"1b46",x"3853",x"3716",x"b7e9",x"baf1",x"2aa7",x"3972",x"2932",x"1c1b",x"3851",x"36eb",x"b776",x"bb0b",x"2d41",x"3977",x"2941",x"9faa",x"385f",x"3712",x"b84e",x"bab0",x"2ec8",x"3972",x"28c9"),
(x"98e9",x"38f1",x"3715",x"b95d",x"39e3",x"2de3",x"3987",x"2c5d",x"9943",x"38f3",x"36eb",x"b9df",x"3964",x"2d28",x"398c",x"2c6f",x"9613",x"38f6",x"3715",x"bbfa",x"2710",x"2c48",x"3988",x"2c55"),
(x"219e",x"386d",x"3713",x"bb5b",x"b634",x"2c03",x"3b20",x"3a4b",x"2166",x"386c",x"36eb",x"bad3",x"b822",x"2c4d",x"3b1c",x"3a4f",x"2010",x"3876",x"370e",x"bb25",x"b70d",x"2d6a",x"3b22",x"3a4d"),
(x"9631",x"381e",x"3716",x"3bff",x"a0b5",x"2138",x"3952",x"3062",x"95be",x"381e",x"36eb",x"3bfe",x"9e8d",x"2828",x"3958",x"3068",x"1624",x"3809",x"370e",x"3b5f",x"35f1",x"2f4d",x"3955",x"304d"),
(x"1cd4",x"3850",x"36eb",x"bb24",x"371c",x"2cde",x"3977",x"294a",x"1c1b",x"3851",x"36eb",x"b776",x"bb0b",x"2d41",x"3977",x"2941",x"1d2c",x"3850",x"3716",x"bbde",x"b1b6",x"2825",x"3971",x"2944"),
(x"9ff6",x"38e8",x"3719",x"b9a6",x"3994",x"2fc6",x"3985",x"2c77",x"a0ef",x"38e8",x"36eb",x"b9ed",x"394b",x"2f45",x"398a",x"2c92",x"98e9",x"38f1",x"3715",x"b95d",x"39e3",x"2de3",x"3987",x"2c5d"),
(x"1f30",x"38c5",x"36eb",x"3bf8",x"2379",x"2d44",x"3997",x"27f5",x"201d",x"38be",x"36eb",x"37d8",x"3af6",x"2a35",x"3997",x"27b6",x"1f03",x"38c0",x"3711",x"3b12",x"3763",x"2ca3",x"3993",x"27d5"),
(x"21a8",x"386a",x"3713",x"bb09",x"3791",x"2ab8",x"3983",x"1da7",x"216e",x"386a",x"36eb",x"b9e9",x"3955",x"2e31",x"3988",x"1d1f",x"219e",x"386d",x"3713",x"bb5b",x"b634",x"2c03",x"3983",x"1d26"),
(x"17ea",x"3831",x"36eb",x"3ab4",x"b859",x"2a66",x"3956",x"307d",x"95be",x"381e",x"36eb",x"3bfe",x"9e8d",x"2828",x"3958",x"3068",x"16e7",x"3832",x"370f",x"3ad7",x"b821",x"29e6",x"3952",x"3079"),
(x"1986",x"384c",x"36eb",x"b97a",x"39b6",x"3099",x"3977",x"2960",x"1cd4",x"3850",x"36eb",x"bb24",x"371c",x"2cde",x"3977",x"294a",x"1ba5",x"384b",x"3714",x"b9e8",x"3951",x"2f27",x"3972",x"295e"),
(x"a09e",x"38e4",x"36eb",x"b2cb",x"bbc1",x"2fc5",x"3989",x"2c99",x"a0ef",x"38e8",x"36eb",x"b9ed",x"394b",x"2f45",x"398a",x"2c92",x"9fe7",x"38e6",x"3719",x"b250",x"bbca",x"2f22",x"3985",x"2c7b"),
(x"1fbf",x"38cd",x"36eb",x"3b57",x"b625",x"2e99",x"3997",x"281d",x"1f30",x"38c5",x"36eb",x"3bf8",x"2379",x"2d44",x"3997",x"27f5",x"1f3f",x"38cf",x"3712",x"3b92",x"b509",x"2cb0",x"3993",x"2829"),
(x"1c5d",x"3862",x"36eb",x"b046",x"3be8",x"2cb7",x"3989",x"1f14",x"216e",x"386a",x"36eb",x"b9e9",x"3955",x"2e31",x"3988",x"1d1f",x"2072",x"3865",x"3710",x"b833",x"3ac7",x"2d1d",x"3984",x"1e78"),
(x"1f0d",x"383c",x"3713",x"37c2",x"baf3",x"2e28",x"3951",x"3087",x"1fba",x"383a",x"36eb",x"373f",x"bb1a",x"2d3c",x"3956",x"308c",x"16e7",x"3832",x"370f",x"3ad7",x"b821",x"29e6",x"3952",x"3079"),
(x"9d26",x"383d",x"36eb",x"baff",x"373c",x"3197",x"3977",x"29bc",x"1986",x"384c",x"36eb",x"b97a",x"39b6",x"3099",x"3977",x"2960",x"9aec",x"383c",x"3717",x"ba77",x"3889",x"310e",x"3972",x"29b5"),
(x"9aa8",x"38e6",x"3718",x"b0c5",x"bbe6",x"2ad9",x"3983",x"2c88",x"9950",x"38e5",x"36eb",x"bb01",x"b745",x"3141",x"3987",x"2cac",x"9fe7",x"38e6",x"3719",x"b250",x"bbca",x"2f22",x"3985",x"2c7b"),
(x"2422",x"38f3",x"36eb",x"3b99",x"b45f",x"30d6",x"3999",x"28c9",x"1fbf",x"38cd",x"36eb",x"3b57",x"b625",x"2e99",x"3997",x"281d",x"2353",x"38f1",x"3711",x"3b70",x"b585",x"3014",x"3994",x"28c4"),
(x"9a03",x"3866",x"36eb",x"374a",x"3b15",x"2de4",x"398a",x"2082",x"1c5d",x"3862",x"36eb",x"b046",x"3be8",x"2cb7",x"3989",x"1f14",x"11f0",x"3862",x"3712",x"32e8",x"3bcb",x"2c10",x"3985",x"2052"),
(x"20b1",x"3839",x"36eb",x"b8ae",x"ba73",x"2d49",x"3b47",x"3a50",x"1fba",x"383a",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b48",x"3a50",x"2079",x"383b",x"3712",x"b722",x"bb24",x"2bf9",x"3b44",x"3a4c"),
(x"a139",x"3821",x"36eb",x"bbbf",x"3113",x"322d",x"3977",x"2a39",x"9d26",x"383d",x"36eb",x"baff",x"373c",x"3197",x"3977",x"29bc",x"a039",x"3821",x"3713",x"bbc6",x"31be",x"30de",x"3972",x"2a2e"),
(x"24be",x"3910",x"36eb",x"3be6",x"ac77",x"308c",x"3999",x"2946",x"2422",x"38f3",x"36eb",x"3b99",x"b45f",x"30d6",x"3999",x"28c9",x"2467",x"3910",x"3711",x"3be4",x"ad1d",x"308c",x"3995",x"294b"),
(x"a0d7",x"3872",x"3717",x"3b6f",x"35e4",x"261e",x"3986",x"2216",x"a09f",x"3872",x"36eb",x"3aaf",x"3860",x"2a70",x"398b",x"2196",x"9ad5",x"3864",x"3711",x"3934",x"3a0d",x"2c16",x"3986",x"20db"),
(x"21ab",x"3835",x"36eb",x"ae28",x"bbe6",x"3005",x"3b46",x"3a51",x"20b1",x"3839",x"36eb",x"b8ae",x"ba73",x"2d49",x"3b47",x"3a50",x"21e0",x"3837",x"3711",x"b5dd",x"bb65",x"2eae",x"3b43",x"3a4d"),
(x"a08e",x"3806",x"3717",x"bbf0",x"2f0f",x"2aec",x"3970",x"2a9d",x"a0d9",x"3806",x"36eb",x"bbea",x"2e0a",x"2f12",x"3976",x"2aaa",x"a039",x"3821",x"3713",x"bbc6",x"31be",x"30de",x"3972",x"2a2e"),
(x"9950",x"38e5",x"36eb",x"bb01",x"b745",x"3141",x"398c",x"2f51",x"9aa8",x"38e6",x"3718",x"b0c5",x"bbe6",x"2ad9",x"398c",x"2f81",x"9920",x"38e4",x"3718",x"baf6",x"37e0",x"2460",x"398d",x"2f80"),
(x"2469",x"3932",x"3714",x"3bec",x"2d02",x"2f4a",x"3995",x"29d9",x"24b3",x"3933",x"36eb",x"3be8",x"2d66",x"3010",x"399a",x"29d7",x"2467",x"3910",x"3711",x"3be4",x"ad1d",x"308c",x"3995",x"294b"),
(x"a180",x"3883",x"3715",x"3bfe",x"a412",x"2867",x"3988",x"231a",x"a166",x"3882",x"36eb",x"3bfa",x"2c62",x"2617",x"398d",x"2295",x"a0d7",x"3872",x"3717",x"3b6f",x"35e4",x"261e",x"3986",x"2216"),
(x"244f",x"3835",x"36eb",x"3913",x"ba0d",x"310f",x"3b43",x"3a52",x"21ab",x"3835",x"36eb",x"ae28",x"bbe6",x"3005",x"3b46",x"3a51",x"23f2",x"3838",x"3712",x"35a6",x"bb63",x"30cc",x"3b41",x"3a4e"),
(x"a243",x"37e1",x"36eb",x"bbe4",x"2adf",x"30ee",x"3975",x"2b06",x"a0d9",x"3806",x"36eb",x"bbea",x"2e0a",x"2f12",x"3976",x"2aaa",x"a1a0",x"37df",x"370f",x"bbdd",x"30de",x"2e6c",x"3971",x"2afe"),
(x"a164",x"38d4",x"36eb",x"bbbf",x"3333",x"2ed0",x"3992",x"2f4c",x"9fd8",x"38dc",x"36eb",x"ba0e",x"3929",x"2e76",x"3990",x"2f4e",x"a0a3",x"38d3",x"3718",x"bb13",x"3732",x"2fec",x"3992",x"2f7c"),
(x"2427",x"3945",x"36eb",x"3ab2",x"3834",x"30cb",x"399a",x"2a24",x"24b3",x"3933",x"36eb",x"3be8",x"2d66",x"3010",x"399a",x"29d7",x"23cf",x"3942",x"3712",x"3b45",x"3640",x"30a6",x"3995",x"2a1c"),
(x"1ea1",x"3921",x"3710",x"3bcc",x"3227",x"2f2f",x"3958",x"24db",x"1f98",x"3921",x"36eb",x"3bf4",x"1edc",x"2ebb",x"395c",x"24c5",x"1de8",x"3919",x"3710",x"3b2f",x"b6d9",x"2e52",x"3957",x"2492"),
(x"a123",x"3899",x"3714",x"3b81",x"b558",x"2da5",x"398a",x"243a",x"a0d8",x"3897",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"398e",x"23e2",x"a180",x"3883",x"3715",x"3bfe",x"a412",x"2867",x"3988",x"231a"),
(x"24ee",x"383f",x"36eb",x"3be5",x"2dbc",x"3036",x"3b40",x"3a53",x"244f",x"3835",x"36eb",x"3913",x"ba0d",x"310f",x"3b43",x"3a52",x"2498",x"383f",x"3711",x"3bb2",x"b32f",x"30f4",x"3b3f",x"3a4f"),
(x"a1da",x"37ca",x"36eb",x"baf6",x"b714",x"32f0",x"3975",x"2b36",x"a243",x"37e1",x"36eb",x"bbe4",x"2adf",x"30ee",x"3975",x"2b06",x"a12d",x"37d1",x"370d",x"bb0d",x"b70c",x"3169",x"3971",x"2b1d"),
(x"a13e",x"38c8",x"36eb",x"bbbf",x"b371",x"2dad",x"3995",x"2f4c",x"a164",x"38d4",x"36eb",x"bbbf",x"3333",x"2ed0",x"3992",x"2f4c",x"a0f6",x"38cb",x"3712",x"bbf0",x"ac20",x"2e95",x"3994",x"2f75"),
(x"20e4",x"3955",x"36eb",x"37cb",x"3ae6",x"3068",x"3999",x"2a7b",x"2427",x"3945",x"36eb",x"3ab2",x"3834",x"30cb",x"399a",x"2a24",x"20a5",x"3951",x"3715",x"393c",x"39e9",x"3110",x"3994",x"2a6f"),
(x"9e13",x"38a8",x"3715",x"3a65",x"b8c1",x"2d9c",x"398b",x"24c4",x"9d2f",x"38a7",x"36eb",x"3ac2",x"b833",x"2e8a",x"3990",x"2480",x"a123",x"3899",x"3714",x"3b81",x"b558",x"2da5",x"398a",x"243a"),
(x"2454",x"384e",x"36eb",x"3902",x"3a23",x"3069",x"3b3c",x"3a54",x"24ee",x"383f",x"36eb",x"3be5",x"2dbc",x"3036",x"3b40",x"3a53",x"242c",x"384b",x"3712",x"3ae4",x"37c3",x"30c9",x"3b3c",x"3a4f"),
(x"a05e",x"37cb",x"3713",x"b451",x"bbac",x"2d81",x"3970",x"2b2a",x"a088",x"37c6",x"36eb",x"b571",x"bb6d",x"30cc",x"3974",x"2b4c",x"a12d",x"37d1",x"370d",x"bb0d",x"b70c",x"3169",x"3971",x"2b1d"),
(x"a0e1",x"38c6",x"36eb",x"aeda",x"bbea",x"2e47",x"3996",x"2f4c",x"a13e",x"38c8",x"36eb",x"bbbf",x"b371",x"2dad",x"3995",x"2f4c",x"a072",x"38c8",x"3712",x"b297",x"bbcc",x"2d84",x"3995",x"2f76"),
(x"177f",x"3959",x"36eb",x"16f6",x"3bf5",x"2e99",x"3999",x"2abf",x"20e4",x"3955",x"36eb",x"37cb",x"3ae6",x"3068",x"3999",x"2a7b",x"1788",x"3956",x"3715",x"1ef6",x"3bee",x"302a",x"3994",x"2ab0"),
(x"9607",x"38b2",x"3717",x"3939",x"ba0b",x"29e0",x"398c",x"252b",x"9470",x"38b1",x"36eb",x"39cd",x"b979",x"2caa",x"3991",x"24e4",x"9e13",x"38a8",x"3715",x"3a65",x"b8c1",x"2d9c",x"398b",x"24c4"),
(x"21e1",x"3850",x"36eb",x"33f1",x"3bbc",x"2b58",x"3b39",x"3a54",x"2454",x"384e",x"36eb",x"3902",x"3a23",x"3069",x"3b3c",x"3a54",x"2226",x"384e",x"3713",x"3607",x"3b5e",x"2e4d",x"3b39",x"3a4f"),
(x"9e25",x"37c9",x"3716",x"b8de",x"ba57",x"297d",x"396f",x"2b3c",x"9e52",x"37c7",x"36eb",x"bbe3",x"ace8",x"30c3",x"3974",x"2b61",x"a05e",x"37cb",x"3713",x"b451",x"bbac",x"2d81",x"3970",x"2b2a"),
(x"9d58",x"38c8",x"3717",x"aa07",x"bbfc",x"284d",x"3997",x"2f7e",x"9ce6",x"38c7",x"36eb",x"ac58",x"bbf7",x"2bc1",x"3998",x"2f50",x"a072",x"38c8",x"3712",x"b297",x"bbcc",x"2d84",x"3995",x"2f76"),
(x"9e4d",x"3951",x"3713",x"b82e",x"3aba",x"306c",x"3993",x"2af7",x"9dfd",x"3955",x"36eb",x"b66a",x"3b44",x"2f81",x"3998",x"2b02",x"1788",x"3956",x"3715",x"1ef6",x"3bee",x"302a",x"3994",x"2ab0"),
(x"125b",x"38b5",x"3717",x"ac93",x"bbf9",x"2918",x"398d",x"2556",x"11e3",x"38b4",x"36eb",x"b5a5",x"bb74",x"2d53",x"3992",x"2508",x"9607",x"38b2",x"3717",x"3939",x"ba0b",x"29e0",x"398c",x"252b"),
(x"212c",x"3852",x"3716",x"3ac7",x"b83c",x"283f",x"3b38",x"3a4f",x"2164",x"3852",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b39",x"3a54",x"2226",x"384e",x"3713",x"3607",x"3b5e",x"2e4d",x"3b39",x"3a4f"),
(x"1624",x"3809",x"370e",x"3004",x"271d",x"3bef",x"3916",x"38c8",x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4",x"a08e",x"3806",x"3717",x"2bf6",x"a5ae",x"3bfb",x"390b",x"38c7"),
(x"9b62",x"38c5",x"36eb",x"ba75",x"b8ad",x"2ccc",x"3999",x"2f51",x"9ce6",x"38c7",x"36eb",x"ac58",x"bbf7",x"2bc1",x"3998",x"2f50",x"9b02",x"38c7",x"3716",x"b8f4",x"ba42",x"2c09",x"3998",x"2f7d"),
(x"a2e7",x"3945",x"3715",x"bae0",x"37cf",x"30d4",x"3992",x"2b45",x"a395",x"3947",x"36eb",x"b9f2",x"3938",x"30b5",x"3997",x"2b5e",x"9e4d",x"3951",x"3713",x"b82e",x"3aba",x"306c",x"3993",x"2af7"),
(x"1e32",x"38a8",x"36eb",x"b976",x"b9cc",x"2dcc",x"3993",x"2580",x"11e3",x"38b4",x"36eb",x"b5a5",x"bb74",x"2d53",x"3992",x"2508",x"1acb",x"38b1",x"3714",x"b9a7",x"b99e",x"2d1e",x"398e",x"2580"),
(x"2433",x"3855",x"36eb",x"39ec",x"b92b",x"31e4",x"3b35",x"3a55",x"2164",x"3852",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b39",x"3a54",x"2360",x"3856",x"3711",x"38c8",x"ba4e",x"30a8",x"3b35",x"3a50"),
(x"9b62",x"38c5",x"36eb",x"ba75",x"b8ad",x"2ccc",x"3999",x"2f51",x"9b02",x"38c7",x"3716",x"b8f4",x"ba42",x"2c09",x"3998",x"2f7d",x"9959",x"38c4",x"3715",x"bb3f",x"b6b6",x"2b9d",x"3999",x"2f7e"),
(x"a44d",x"3933",x"3715",x"bbec",x"2be2",x"2fce",x"3990",x"2b92",x"a493",x"3934",x"36eb",x"bbc4",x"327a",x"3012",x"3995",x"2bae",x"a2e7",x"3945",x"3715",x"bae0",x"37cf",x"30d4",x"3992",x"2b45"),
(x"20ef",x"38a3",x"36eb",x"b53f",x"bb87",x"2d28",x"3994",x"25c5",x"1e32",x"38a8",x"36eb",x"b976",x"b9cc",x"2dcc",x"3993",x"2580",x"2116",x"38a4",x"3716",x"b7d5",x"baf0",x"2d8e",x"3990",x"260f"),
(x"2563",x"3866",x"36eb",x"3bbc",x"b212",x"3175",x"3b30",x"3a55",x"2433",x"3855",x"36eb",x"39ec",x"b92b",x"31e4",x"3b35",x"3a55",x"24fa",x"3866",x"370f",x"3b4b",x"b5cc",x"3223",x"3b30",x"3a51"),
(x"9f92",x"377e",x"36eb",x"bade",x"b7ab",x"31d3",x"395a",x"2f8e",x"a0ba",x"37ad",x"36eb",x"bbdb",x"9c67",x"320a",x"3957",x"2f62",x"9e24",x"3783",x"370e",x"bb7b",x"b4a9",x"3270",x"3956",x"2f9c"),
(x"a0d7",x"38b5",x"36eb",x"bafe",x"375c",x"30f4",x"3975",x"2683",x"9959",x"38c4",x"3715",x"ba5f",x"3873",x"3388",x"396f",x"25f6",x"9ec5",x"38b7",x"3718",x"bac6",x"37dc",x"3286",x"3970",x"2672"),
(x"a409",x"3922",x"3717",x"bb55",x"b5fd",x"307e",x"398e",x"2bd3",x"a46a",x"3921",x"36eb",x"bb6e",x"b575",x"309f",x"3993",x"2bf8",x"a44d",x"3933",x"3715",x"bbec",x"2be2",x"2fce",x"3990",x"2b92"),
(x"2353",x"38f1",x"3711",x"3115",x"a7d5",x"3be4",x"3927",x"394c",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b",x"2002",x"38f9",x"3714",x"305e",x"a1a1",x"3bec",x"3920",x"3951"),
(x"2357",x"38a1",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3995",x"2610",x"20ef",x"38a3",x"36eb",x"b53f",x"bb87",x"2d28",x"3994",x"25c5",x"2323",x"38a3",x"3716",x"2345",x"bbf7",x"2dcc",x"3990",x"2650"),
(x"2574",x"387a",x"36eb",x"3b61",x"35a0",x"3119",x"3b2b",x"3a55",x"2563",x"3866",x"36eb",x"3bbc",x"b212",x"3175",x"3b30",x"3a55",x"2517",x"3879",x"370f",x"3bd3",x"2f46",x"3182",x"3b2b",x"3a50"),
(x"a348",x"389f",x"36eb",x"bbba",x"3376",x"2f14",x"3976",x"2750",x"a0d7",x"38b5",x"36eb",x"bafe",x"375c",x"30f4",x"3975",x"2683",x"a29f",x"389f",x"3714",x"bb6b",x"3587",x"3096",x"3971",x"2754"),
(x"a22e",x"3911",x"36eb",x"b884",x"ba69",x"3249",x"3991",x"2c1f",x"a46a",x"3921",x"36eb",x"bb6e",x"b575",x"309f",x"3993",x"2bf8",x"a18f",x"3914",x"3711",x"b8a4",x"ba69",x"309a",x"398d",x"2c0c"),
(x"24b8",x"38a5",x"36eb",x"3acc",x"b812",x"3064",x"3996",x"265b",x"2357",x"38a1",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3995",x"2610",x"245f",x"38a6",x"3714",x"3976",x"b9c0",x"3023",x"3991",x"2689"),
(x"2449",x"3886",x"36eb",x"386e",x"3a87",x"313e",x"3b27",x"3a54",x"2574",x"387a",x"36eb",x"3b61",x"35a0",x"3119",x"3b2b",x"3a55",x"2437",x"3883",x"370f",x"3891",x"3a72",x"30f5",x"3b28",x"3a50"),
(x"1222",x"3756",x"36eb",x"b8a6",x"ba54",x"3207",x"395d",x"2fc0",x"9f92",x"377e",x"36eb",x"bade",x"b7ab",x"31d3",x"395a",x"2f8e",x"0f4a",x"3761",x"3712",x"b8b5",x"ba3e",x"32bc",x"3958",x"2fc7"),
(x"a41c",x"3885",x"36eb",x"bbef",x"ad0b",x"2e69",x"3977",x"2816",x"a348",x"389f",x"36eb",x"bbba",x"3376",x"2f14",x"3976",x"2750",x"a3b3",x"3886",x"3712",x"bbf0",x"2a00",x"2f46",x"3972",x"2814"),
(x"9a89",x"390e",x"3718",x"b8ae",x"ba78",x"2b7c",x"398a",x"2c25",x"9bc5",x"390e",x"36eb",x"b60d",x"bb5a",x"2ef3",x"398f",x"2c3d",x"a18f",x"3914",x"3711",x"b8a4",x"ba69",x"309a",x"398d",x"2c0c"),
(x"2515",x"38b0",x"36eb",x"3bcf",x"3174",x"303e",x"3997",x"26b6",x"24b8",x"38a5",x"36eb",x"3acc",x"b812",x"3064",x"3996",x"265b",x"24ba",x"38af",x"3712",x"3be0",x"ae5e",x"30a3",x"3992",x"26ce"),
(x"221a",x"3885",x"3713",x"b583",x"3b63",x"3153",x"3b26",x"3a4f",x"21a6",x"3888",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b24",x"3a53",x"2437",x"3883",x"370f",x"3891",x"3a72",x"30f5",x"3b28",x"3a50"),
(x"1c89",x"3761",x"3716",x"3add",x"b75a",x"334d",x"3958",x"2fd9",x"1dd1",x"3756",x"36eb",x"3996",x"b95f",x"33ec",x"395d",x"2fd5",x"0f4a",x"3761",x"3712",x"b8b5",x"ba3e",x"32bc",x"3958",x"2fc7"),
(x"a2ed",x"386d",x"36eb",x"bb75",x"b5a2",x"2d46",x"3977",x"287b",x"a41c",x"3885",x"36eb",x"bbef",x"ad0b",x"2e69",x"3977",x"2816",x"a294",x"386e",x"3710",x"bb6b",x"b5ba",x"2efe",x"3972",x"287b"),
(x"9747",x"3909",x"3718",x"bbe6",x"b09e",x"2baa",x"398a",x"2c2f",x"990f",x"3909",x"36eb",x"bbe6",x"b08e",x"2c41",x"398e",x"2c46",x"9a89",x"390e",x"3718",x"b8ae",x"ba78",x"2b7c",x"398a",x"2c25"),
(x"247a",x"38ba",x"36eb",x"36fe",x"3b25",x"2ea4",x"3997",x"2711",x"2515",x"38b0",x"36eb",x"3bcf",x"3174",x"303e",x"3997",x"26b6",x"2458",x"38b7",x"3714",x"3972",x"39bb",x"30de",x"3992",x"2716"),
(x"235a",x"3925",x"3710",x"a828",x"a60a",x"3bfe",x"3928",x"396a",x"2325",x"3935",x"3714",x"a946",x"9ffc",x"3bfe",x"3928",x"3972",x"2469",x"3932",x"3714",x"aeb0",x"a8fa",x"3bf3",x"392b",x"3971"),
(x"227e",x"393d",x"3712",x"a953",x"a7ae",x"3bfd",x"3927",x"3977",x"214b",x"3944",x"3714",x"28bf",x"ac20",x"3bfa",x"3924",x"397b",x"23cf",x"3942",x"3712",x"2587",x"a08e",x"3bff",x"3929",x"397a"),
(x"1f1f",x"3949",x"3714",x"a31d",x"ab5f",x"3bfc",x"3921",x"397e",x"20a5",x"3951",x"3715",x"20ea",x"aafd",x"3bfc",x"3923",x"3983",x"214b",x"3944",x"3714",x"28bf",x"ac20",x"3bfa",x"3924",x"397b"),
(x"11db",x"394d",x"3715",x"a70a",x"2779",x"3bfe",x"391a",x"3981",x"1788",x"3956",x"3715",x"a7e2",x"a9b2",x"3bfc",x"391c",x"3986",x"1f1f",x"3949",x"3714",x"a31d",x"ab5f",x"3bfc",x"3921",x"397e"),
(x"9d99",x"394a",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3914",x"397f",x"9e4d",x"3951",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3913",x"3984",x"11db",x"394d",x"3715",x"a70a",x"2779",x"3bfe",x"391a",x"3981"),
(x"a14f",x"393d",x"3714",x"28e0",x"a99e",x"3bfc",x"390e",x"3979",x"a2e7",x"3945",x"3715",x"2266",x"1d87",x"3bff",x"390b",x"397d",x"9d99",x"394a",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3914",x"397f"),
(x"a1ee",x"3932",x"3714",x"2538",x"29ab",x"3bfd",x"390c",x"3972",x"a44d",x"3933",x"3715",x"288e",x"27ce",x"3bfd",x"3907",x"3973",x"a14f",x"393d",x"3714",x"28e0",x"a99e",x"3bfc",x"390e",x"3979"),
(x"a1ee",x"3932",x"3714",x"2538",x"29ab",x"3bfd",x"390c",x"3972",x"a0ed",x"3929",x"3715",x"2c67",x"a8a5",x"3bf9",x"390e",x"396d",x"a44d",x"3933",x"3715",x"288e",x"27ce",x"3bfd",x"3907",x"3973"),
(x"9ddf",x"3928",x"3714",x"2a45",x"ab10",x"3bfa",x"3912",x"396c",x"a18f",x"3914",x"3711",x"28d9",x"252b",x"3bfe",x"390c",x"3962",x"a0ed",x"3929",x"3715",x"2c67",x"a8a5",x"3bf9",x"390e",x"396d"),
(x"1937",x"392d",x"3710",x"2352",x"2e80",x"3bf5",x"391b",x"396f",x"1d11",x"3928",x"3711",x"2bef",x"28a8",x"3bfa",x"391e",x"396c",x"9908",x"392c",x"3711",x"2a66",x"331a",x"3bca",x"3916",x"396f"),
(x"9747",x"3909",x"3718",x"3420",x"9418",x"3bba",x"3916",x"395a",x"9a89",x"390e",x"3718",x"2b65",x"3528",x"3b8f",x"3914",x"395d",x"18c5",x"3910",x"3713",x"341f",x"2c3a",x"3bb6",x"391a",x"395e"),
(x"1832",x"3906",x"3714",x"2de0",x"24c2",x"3bf6",x"391a",x"3958",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b",x"9613",x"38f6",x"3715",x"27ae",x"24ea",x"3bfe",x"3916",x"394f"),
(x"1d11",x"3928",x"3711",x"2bef",x"28a8",x"3bfa",x"391e",x"396c",x"1de8",x"3919",x"3710",x"2856",x"29ab",x"3bfc",x"391e",x"3963",x"9ddf",x"3928",x"3714",x"2a45",x"ab10",x"3bfa",x"3912",x"396c"),
(x"98e9",x"38f1",x"3715",x"a8bf",x"2fda",x"3bef",x"3915",x"394d",x"9613",x"38f6",x"3715",x"27ae",x"24ea",x"3bfe",x"3916",x"394f",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b"),
(x"199d",x"390f",x"36eb",x"3bf6",x"aa70",x"2d61",x"395b",x"2417",x"1c29",x"38ee",x"36eb",x"346a",x"3b91",x"316a",x"395a",x"2202",x"1832",x"3906",x"3714",x"3bf3",x"2e23",x"2b27",x"3956",x"23d5"),
(x"22bc",x"3a9c",x"36eb",x"3adb",x"b7e7",x"30ac",x"396a",x"2d88",x"1f7b",x"3a8c",x"36eb",x"3b71",x"b58a",x"2fc3",x"396a",x"2d60",x"1e77",x"3a8d",x"3715",x"3ac1",x"b812",x"3146",x"3964",x"2d67"),
(x"b930",x"3c7f",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0",x"b92a",x"3c7f",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b92b",x"3c69",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa"),
(x"b92a",x"3c7f",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b922",x"3c7f",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b924",x"3c69",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392"),
(x"b922",x"3c7f",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b91b",x"3c7f",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b91f",x"3c69",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387"),
(x"b91b",x"3c7f",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b913",x"3c7f",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b918",x"3c69",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b"),
(x"b913",x"3c7f",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b913",x"3c81",x"373a",x"3ae3",x"2b4f",x"380a",x"3bb9",x"399f",x"b90e",x"3c81",x"370e",x"3754",x"3ae5",x"32eb",x"3bbd",x"39a7"),
(x"b913",x"3c81",x"373a",x"3ae3",x"2b4f",x"380a",x"3bb9",x"399f",x"b913",x"3c7f",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b91b",x"3c7f",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b"),
(x"b913",x"3c81",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1",x"b913",x"3c96",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b90f",x"3c96",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7"),
(x"b90f",x"3c96",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7",x"b90e",x"3c81",x"370e",x"3bcb",x"a949",x"330f",x"3bf9",x"39fa",x"b913",x"3c81",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1"),
(x"b913",x"3c96",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b913",x"3c81",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1",x"b91b",x"3c81",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed"),
(x"b91a",x"3c96",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b91b",x"3c81",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed",x"b924",x"3c82",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b928",x"3c96",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b922",x"3c96",x"3751",x"a11e",x"aa52",x"3bfd",x"3be8",x"39eb",x"b924",x"3c82",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b92f",x"3c96",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b928",x"3c96",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b92b",x"3c81",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6"),
(x"b935",x"3c96",x"3725",x"bb50",x"a63f",x"3678",x"3be8",x"39de",x"b92f",x"3c96",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b930",x"3c81",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3"),
(x"b930",x"3c81",x"3738",x"b75a",x"bae5",x"32d3",x"3bb5",x"3992",x"b92a",x"3c7f",x"3733",x"b800",x"ba99",x"3436",x"3bb7",x"3993",x"b930",x"3c7f",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c"),
(x"b913",x"3c7f",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b90c",x"3c68",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352",x"b912",x"3c69",x"373c",x"3aea",x"2832",x"3802",x"39f2",x"336a"),
(x"b913",x"3c7f",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b90c",x"3c68",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352"),
(x"b91b",x"3c81",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b91b",x"3c7f",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b",x"b922",x"3c7f",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998"),
(x"b922",x"3c7f",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998",x"b92a",x"3c7f",x"3733",x"b800",x"ba99",x"3436",x"3bb7",x"3993",x"b92b",x"3c81",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b935",x"3c96",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b93a",x"3c96",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"3861",x"b931",x"3c97",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b92f",x"3c96",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b935",x"3c96",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b92a",x"3c97",x"3739",x"b604",x"3b4b",x"3148",x"3b22",x"386b"),
(x"b928",x"3c96",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e",x"b92f",x"3c96",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b925",x"3c97",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e"),
(x"b91a",x"3c96",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b922",x"3c96",x"3751",x"9ac2",x"39ac",x"39a3",x"3b24",x"3871",x"b920",x"3c97",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871"),
(x"b913",x"3c96",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b91a",x"3c96",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b919",x"3c97",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873"),
(x"b90f",x"3c96",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879",x"b913",x"3c96",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b913",x"3c98",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875"),
(x"b90d",x"3c96",x"3711",x"b36d",x"a40b",x"3bc7",x"3a19",x"3349",x"b906",x"3c97",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b92f",x"3cae",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b92a",x"3c97",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b931",x"3c97",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4"),
(x"b92a",x"3c97",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b92c",x"3cae",x"373a",x"baa5",x"a5fd",x"3872",x"3a2d",x"33a3",x"b925",x"3cae",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b920",x"3c97",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b925",x"3c97",x"3746",x"b918",x"a84d",x"3a28",x"3a1a",x"338e",x"b925",x"3cae",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b919",x"3c97",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b920",x"3c97",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b91f",x"3cae",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385"),
(x"b913",x"3c98",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b919",x"3c97",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b918",x"3cad",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a2d",x"3378"),
(x"b913",x"3c98",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b911",x"3cae",x"373c",x"3ac9",x"a6b5",x"383a",x"3a2d",x"3366",x"b90b",x"3cad",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c"),
(x"b90b",x"3c97",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b90b",x"3cad",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c",x"b907",x"3cae",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340"),
(x"b116",x"3c8f",x"3710",x"8000",x"0000",x"3c00",x"3a13",x"2451",x"b116",x"3c87",x"3710",x"8000",x"0000",x"3c00",x"3a0c",x"2451",x"b135",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"b135",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b135",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1",x"b161",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f"),
(x"b161",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b161",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f",x"b1a1",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643"),
(x"b1a1",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643",x"b1c1",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"26b3",x"b1c1",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"b1c1",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3",x"b1c1",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"26b3",x"b1fd",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b"),
(x"b1fd",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b",x"b22d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"281a",x"b22d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"b22d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a",x"b22d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"281a",x"b261",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878"),
(x"b261",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b261",x"3c7a",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878",x"b2aa",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"b2aa",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b2aa",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb",x"b2d6",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949"),
(x"b2d6",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b2d6",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949",x"b326",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"b326",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b326",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7",x"b34f",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"b451",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b50c",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2d8d",x"b50c",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"b451",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b451",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2c3f",x"b441",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"b441",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b441",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b34f",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"b40b",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b84",x"b3f4",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b413",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"b3f4",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b3d2",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b409",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"b3d2",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b3a5",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b407",x"3ca0",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"b40b",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b84",x"b413",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2ba0",x"b413",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"b3f4",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b413",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0",x"b409",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"b3d2",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b409",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d",x"b407",x"3c76",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"b3a5",x"3c6e",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b407",x"3c76",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76",x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b3a5",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b368",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b50c",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d",x"b50c",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2d8d",x"b526",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"b62a",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b",x"b62a",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2f8b",x"b5ce",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"b5ce",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7",x"b5bd",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ec9",x"b5bd",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"b5bd",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9",x"b5bd",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ec9",x"b5a1",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"b5a1",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b5a1",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97",x"b581",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"b581",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e",x"b568",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b568",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b50d",x"3cb2",x"3710",x"8000",x"0000",x"3c00",x"3a30",x"2d8e",x"b4f9",x"3caf",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"2d6a",x"b4f5",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"b52b",x"3cb1",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b4f5",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63",x"b4f2",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b4f5",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b4f9",x"3c67",x"3710",x"8000",x"0000",x"3c00",x"39f0",x"2d6a",x"b50d",x"3c65",x"3710",x"8000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"b4f2",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b4f5",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b52b",x"3c65",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"b568",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2e32",x"b575",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2e49",x"b575",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"b558",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b575",x"3c70",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47",x"b569",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"b568",x"3cad",x"3710",x"8000",x"0000",x"3c00",x"3a2c",x"2e32",x"b558",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b575",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"b558",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b544",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0",x"b569",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"b4e1",x"3c9d",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2d40",x"b51a",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b4da",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"b4e1",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"2d40",x"b4d8",x"3c77",x"3710",x"8000",x"0000",x"3c00",x"39fe",x"2d2f",x"b4da",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"b51a",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4da",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33",x"b4f2",x"3c6d",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"b51a",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b528",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b4f2",x"3ca9",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b528",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b569",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33",x"b544",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"b544",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b569",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33",x"b528",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"b528",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b52c",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5",x"b568",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"b528",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b569",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33",x"b568",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b526",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb",x"b52c",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5",x"b52c",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"b568",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b52c",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5",x"b52c",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"b63d",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b62a",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2f8b",x"b62a",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"b669",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b63d",x"3c97",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b63d",x"3c7f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"b669",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b669",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2ffc",x"b721",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b72d",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b721",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30a2",x"b721",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b794",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b7c0",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130",x"b7c0",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130"),
(x"b794",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b794",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"3109",x"b77a",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"b77a",x"3c7d",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b77a",x"3c99",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1",x"b776",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b776",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b776",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed",x"b72d",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"b6fb",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b6ef",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3075",x"b6f1",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3076"),
(x"b721",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b6fb",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b705",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088"),
(x"b6f1",x"3ca8",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"3076",x"b6ef",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3075",x"b6fb",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080"),
(x"b705",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b6fb",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080",x"b721",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"b73e",x"3caf",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b721",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2",x"b72e",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b72e",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b721",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b73e",x"3c67",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"b7c7",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3135",x"b7c7",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"3136",x"b7bd",x"3c73",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d"),
(x"b7c7",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3135",x"b7a4",x"3cab",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b7bd",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d"),
(x"b7a4",x"3cab",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b783",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b7a8",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a"),
(x"b7a4",x"3c6c",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7bd",x"3c73",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d",x"b7a8",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a"),
(x"b72e",x"3c7e",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b77b",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b776",x"3c7b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"b72e",x"3c98",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae",x"b72d",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b776",x"3c9c",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b77b",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b783",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b790",x"3c76",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3107"),
(x"b801",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b7c0",x"3c94",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130",x"b7c0",x"3c82",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130"),
(x"b820",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b801",x"3c96",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b801",x"3c80",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b"),
(x"b820",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b820",x"3c79",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"31a2",x"b83a",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b84a",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b83a",x"3cab",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"31d0",x"b83a",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b85e",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b84a",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b84a",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"b865",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b85e",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b85e",x"3c6a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211"),
(x"b867",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b865",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b865",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d"),
(x"b867",x"3ca4",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b867",x"3c72",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"3222",x"b86e",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b87d",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b86e",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"322d",x"b86e",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b88f",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b87d",x"3ca2",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b87d",x"3c74",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248"),
(x"b88f",x"3ca7",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b88f",x"3c6f",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"3269",x"b89e",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b8a3",x"3cac",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b89e",x"3cac",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3284",x"b89e",x"3c6b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b8a3",x"3cac",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b8a3",x"3c6a",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b907",x"3c80",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b8ff",x"3cae",x"3710",x"2904",x"26d5",x"3bfd",x"3a2d",x"3331",x"b8a3",x"3cac",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b906",x"3c97",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d"),
(x"b918",x"3cad",x"374b",x"270a",x"3bfd",x"2877",x"3bce",x"3a59",x"b91f",x"3cae",x"374f",x"28f4",x"3bfa",x"ac28",x"3bcd",x"3a5c",x"b925",x"3cae",x"3749",x"257a",x"3bfd",x"28f4",x"3bcf",x"3a5e"),
(x"b911",x"3cae",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b925",x"3cae",x"3749",x"257a",x"3bfd",x"28f4",x"3bcf",x"3a5e",x"b92c",x"3cae",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60"),
(x"b90b",x"3cad",x"3722",x"2773",x"3bfe",x"22cf",x"3bd6",x"3a54",x"b92c",x"3cae",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60",x"b92f",x"3cae",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62"),
(x"b907",x"3cae",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b92f",x"3cae",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62",x"b931",x"3cae",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63"),
(x"b924",x"3c69",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b91f",x"3c69",x"374e",x"281b",x"bbe6",x"b0f4",x"3a92",x"3a5c",x"b918",x"3c69",x"374b",x"2511",x"bbff",x"224c",x"3a91",x"3a59"),
(x"b92b",x"3c69",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b924",x"3c69",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b912",x"3c69",x"373c",x"1818",x"bbff",x"26c2",x"3a8e",x"3a57"),
(x"b931",x"3c69",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63",x"b92b",x"3c69",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b90c",x"3c68",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55"),
(x"b1fd",x"3c7a",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b22d",x"3c78",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b22d",x"3c78",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94"),
(x"b6fb",x"3c78",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6ef",x"3c74",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6ef",x"3c74",x"3710",x"3b57",x"3658",x"0000",x"3a95",x"3a0c"),
(x"b63d",x"3c97",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b62a",x"3c97",x"36da",x"303b",x"3bed",x"8000",x"3a97",x"39f9",x"b62a",x"3c97",x"3710",x"2fbb",x"3bf1",x"0000",x"3aa1",x"39f9"),
(x"b1c1",x"3c7e",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1fd",x"3c7a",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b1fd",x"3c7a",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90"),
(x"b906",x"3c69",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b931",x"3c69",x"36da",x"9e3f",x"bc00",x"0000",x"3a7b",x"3a63",x"b931",x"3c69",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63"),
(x"b721",x"3c7c",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b6fb",x"3c78",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6fb",x"3c78",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08"),
(x"b575",x"3ca7",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"3ca9",x"36da",x"bab5",x"385c",x"8a8d",x"3a97",x"3a28",x"b575",x"3ca9",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28"),
(x"b1a1",x"3c7f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1c1",x"3c7e",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1c1",x"3c7e",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89"),
(x"b72e",x"3c7e",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b721",x"3c7c",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b721",x"3c7c",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00"),
(x"b62a",x"3c97",x"36da",x"303b",x"3bed",x"8000",x"3a97",x"39f9",x"b5ce",x"3c94",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5ce",x"3c94",x"3710",x"2f26",x"3bf3",x"0000",x"3aa1",x"3a0b"),
(x"b161",x"3c80",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b1a1",x"3c7f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1a1",x"3c7f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86"),
(x"b72d",x"3c80",x"36da",x"3a45",x"b8f8",x"0000",x"3a8a",x"39fb",x"b72e",x"3c7e",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b72e",x"3c7e",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd"),
(x"b5ce",x"3c94",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5bd",x"3c95",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5bd",x"3c95",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e"),
(x"b135",x"3c82",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b161",x"3c80",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b161",x"3c80",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80"),
(x"b721",x"3c81",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b72d",x"3c80",x"36da",x"3a45",x"b8f8",x"0000",x"3a7c",x"3bb2",x"b72d",x"3c80",x"3710",x"3778",x"bb13",x"0000",x"3a87",x"3bb2"),
(x"b5bd",x"3c95",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5a1",x"3c99",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b5a1",x"3c99",x"3710",x"b72c",x"3b26",x"8000",x"3aa1",x"3a14"),
(x"b93a",x"3c96",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"385a",x"b931",x"3c97",x"36da",x"b311",x"3bcd",x"0000",x"3b16",x"385d",x"b931",x"3c97",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b116",x"3c87",x"36da",x"3b51",x"b675",x"0000",x"3a6e",x"3b77",x"b135",x"3c82",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b135",x"3c82",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b"),
(x"b568",x"3c6a",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b575",x"3c6d",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3c6d",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52"),
(x"b5a1",x"3c99",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b581",x"3c9c",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b581",x"3c9c",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a"),
(x"b669",x"3c81",x"36da",x"a65f",x"bbff",x"0000",x"3a7c",x"3b8d",x"b721",x"3c81",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b721",x"3c81",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf"),
(x"b581",x"3c9c",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b568",x"3ca1",x"36da",x"bb03",x"37b2",x"068d",x"3a97",x"3a21",x"b568",x"3ca1",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21"),
(x"b8a3",x"3c6a",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b906",x"3c69",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b906",x"3c69",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53"),
(x"b63d",x"3c7f",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b669",x"3c81",x"36da",x"a65f",x"bbff",x"0000",x"3a7c",x"3b8d",x"b669",x"3c81",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d"),
(x"b568",x"3cad",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b558",x"3cae",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b558",x"3cae",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f"),
(x"b62a",x"3c7f",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b63d",x"3c7f",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b63d",x"3c7f",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84"),
(x"b558",x"3cae",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b544",x"3cae",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b544",x"3cae",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32"),
(x"b575",x"3c6d",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3c70",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b575",x"3c70",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54"),
(x"b544",x"3cae",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b52b",x"3cb1",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b52b",x"3cb1",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37"),
(x"b5ce",x"3c82",x"36da",x"2f26",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b62a",x"3c7f",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b62a",x"3c7f",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81"),
(x"b52b",x"3cb1",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b50d",x"3cb2",x"36da",x"324a",x"3bd8",x"0000",x"3a97",x"3a3d",x"b50d",x"3cb2",x"3710",x"253f",x"3bff",x"8000",x"3aa1",x"3a3d"),
(x"b5bd",x"3c82",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5ce",x"3c82",x"36da",x"2f26",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b5ce",x"3c82",x"3710",x"2ae9",x"bbfc",x"0000",x"3a87",x"3b6f"),
(x"b50d",x"3cb2",x"36da",x"324a",x"3bd8",x"0000",x"3a97",x"3a3d",x"b4f9",x"3caf",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f9",x"3caf",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41"),
(x"b5a1",x"3c7e",x"36da",x"b72c",x"bb26",x"8000",x"3a7c",x"3b66",x"b5bd",x"3c82",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5bd",x"3c82",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c"),
(x"b4f9",x"3caf",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f5",x"3cac",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f5",x"3cac",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44"),
(x"b581",x"3c7b",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b5a1",x"3c7e",x"36da",x"b72c",x"bb26",x"8000",x"3a7c",x"3b66",x"b5a1",x"3c7e",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66"),
(x"b4f5",x"3cac",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f2",x"3ca9",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4f2",x"3ca9",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47"),
(x"b931",x"3c97",x"36da",x"bbff",x"a4d0",x"0000",x"3a18",x"33f3",x"b931",x"3cae",x"36da",x"bbff",x"a4d0",x"0000",x"3a2c",x"33f9",x"b931",x"3cae",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9"),
(x"b8ff",x"3cae",x"36da",x"26a1",x"3bff",x"8000",x"3be3",x"3a4f",x"b8a3",x"3cac",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b8a3",x"3cac",x"3710",x"286d",x"3bfe",x"8000",x"3bd9",x"3a2b"),
(x"b568",x"3c75",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b581",x"3c7b",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b581",x"3c7b",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f"),
(x"b4f2",x"3ca9",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4da",x"3ca2",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4da",x"3ca2",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d"),
(x"b8a3",x"3cac",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b89e",x"3cac",x"36da",x"380f",x"3ae4",x"068d",x"3be3",x"3a29",x"b89e",x"3cac",x"3710",x"36f0",x"3b35",x"0000",x"3bd9",x"3a29"),
(x"b558",x"3c68",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b568",x"3c6a",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b568",x"3c6a",x"3710",x"b810",x"bae4",x"868d",x"3a87",x"3b4e"),
(x"b4da",x"3ca2",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4d8",x"3c9f",x"36da",x"3af9",x"b7d8",x"8000",x"3a97",x"3a50",x"b4d8",x"3c9f",x"3710",x"3be5",x"b11d",x"868d",x"3aa1",x"3a50"),
(x"b89e",x"3cac",x"36da",x"380f",x"3ae4",x"068d",x"3be3",x"3a29",x"b88f",x"3ca7",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b88f",x"3ca7",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22"),
(x"b544",x"3c68",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b558",x"3c68",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b558",x"3c68",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b"),
(x"b4d8",x"3c9f",x"36da",x"3af9",x"b7d8",x"8000",x"3a97",x"3a50",x"b4e1",x"3c9d",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b4e1",x"3c9d",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52"),
(x"b88f",x"3ca7",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b87d",x"3ca2",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b87d",x"3ca2",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a"),
(x"b52b",x"3c65",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b544",x"3c68",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b544",x"3c68",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47"),
(x"b4e1",x"3c9d",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b51a",x"3c9a",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b51a",x"3c9a",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d"),
(x"b87d",x"3ca2",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b86e",x"3ca2",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b86e",x"3ca2",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14"),
(x"b50d",x"3c65",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b52b",x"3c65",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b52b",x"3c65",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42"),
(x"b51a",x"3c9a",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b528",x"3c99",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b528",x"3c99",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60"),
(x"b86e",x"3ca2",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b867",x"3ca4",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b867",x"3ca4",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11"),
(x"b4f9",x"3c67",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b50d",x"3c65",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b50d",x"3c65",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c"),
(x"b528",x"3c99",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b52c",x"3c98",x"36da",x"3b0d",x"378c",x"0000",x"3a97",x"3a61",x"b52c",x"3c98",x"3710",x"3bfc",x"ab6c",x"0000",x"3aa1",x"3a61"),
(x"b867",x"3ca4",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b865",x"3ca7",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b865",x"3ca7",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e"),
(x"b4f5",x"3c6a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f9",x"3c67",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b4f9",x"3c67",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38"),
(x"b52c",x"3c98",x"36da",x"3b0d",x"378c",x"0000",x"3a54",x"39ec",x"b526",x"3c96",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b526",x"3c96",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee"),
(x"b865",x"3ca7",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b85e",x"3cac",x"36da",x"b5f3",x"3b6d",x"8000",x"3be3",x"3a09",x"b85e",x"3cac",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09"),
(x"b4f2",x"3c6d",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f5",x"3c6a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f5",x"3c6a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35"),
(x"b526",x"3c96",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b50c",x"3c95",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b50c",x"3c95",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3"),
(x"b116",x"3c8f",x"36da",x"3bdf",x"31b0",x"868d",x"3a6e",x"3b70",x"b116",x"3c87",x"36da",x"3b51",x"b675",x"0000",x"3a6e",x"3b77",x"b116",x"3c87",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77"),
(x"b85e",x"3cac",x"36da",x"b5f3",x"3b6d",x"8000",x"3be3",x"3a09",x"b84a",x"3cae",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b84a",x"3cae",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01"),
(x"b4da",x"3c74",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4f2",x"3c6d",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f2",x"3c6d",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33"),
(x"b451",x"3c95",x"36da",x"a987",x"3bfe",x"8000",x"3a54",x"3a16",x"b441",x"3c96",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b441",x"3c96",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19"),
(x"b89e",x"3c6b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b8a3",x"3c6a",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b8a3",x"3c6a",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d"),
(x"b84a",x"3cae",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b83a",x"3cab",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b83a",x"3cab",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa"),
(x"b4d8",x"3c77",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4da",x"3c74",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4da",x"3c74",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c"),
(x"b50c",x"3c95",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b451",x"3c95",x"36da",x"a987",x"3bfe",x"8000",x"3a54",x"3a16",x"b451",x"3c95",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16"),
(x"b88f",x"3c6f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b89e",x"3c6b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b89e",x"3c6b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b"),
(x"b568",x"3ca1",x"36da",x"bb03",x"37b2",x"068d",x"3a97",x"3a21",x"b569",x"3ca4",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b569",x"3ca4",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23"),
(x"b4e1",x"3c79",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4d8",x"3c77",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4d8",x"3c77",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a"),
(x"b441",x"3c96",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b40d",x"3c9e",x"36da",x"b8bf",x"3a70",x"8000",x"3a54",x"3a25",x"b40d",x"3c9e",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25"),
(x"b87d",x"3c74",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b88f",x"3c6f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b88f",x"3c6f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25"),
(x"b83a",x"3cab",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b820",x"3c9e",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b820",x"3c9e",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec"),
(x"b51a",x"3c7c",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b4e1",x"3c79",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4e1",x"3c79",x"3710",x"33d2",x"3bc1",x"0000",x"3a87",x"3b28"),
(x"b40d",x"3c9e",x"36da",x"b8bf",x"3a70",x"8000",x"3a54",x"3a25",x"b407",x"3ca0",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b407",x"3ca0",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27"),
(x"b86e",x"3c74",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b87d",x"3c74",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b87d",x"3c74",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d"),
(x"b569",x"3ca4",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b575",x"3ca7",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"3ca7",x"3710",x"ba67",x"b8cb",x"068d",x"3aa1",x"3a26"),
(x"b528",x"3c7e",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b51a",x"3c7c",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b51a",x"3c7c",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d"),
(x"b407",x"3ca0",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b409",x"3ca2",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b409",x"3ca2",x"3710",x"bb1a",x"b75c",x"0000",x"3a5f",x"3a28"),
(x"b867",x"3c72",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b86e",x"3c74",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b86e",x"3c74",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17"),
(x"b820",x"3c9e",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b801",x"3c96",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b801",x"3c96",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de"),
(x"b52c",x"3c7f",x"36da",x"3bfc",x"2b6c",x"0000",x"3a7c",x"3b19",x"b528",x"3c7e",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b528",x"3c7e",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a"),
(x"b409",x"3ca2",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b413",x"3ca5",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"3ca5",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b"),
(x"b865",x"3c6f",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b867",x"3c72",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b867",x"3c72",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14"),
(x"b801",x"3c96",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b7c0",x"3c94",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b7c0",x"3c94",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1"),
(x"b526",x"3c80",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b52c",x"3c7f",x"36da",x"3bfc",x"2b6c",x"0000",x"3afb",x"3a11",x"b52c",x"3c7f",x"3710",x"3b0d",x"b78c",x"0000",x"3b06",x"3a11"),
(x"b413",x"3ca5",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"3ca7",x"36da",x"ba12",x"3935",x"8000",x"3a54",x"3a2d",x"b413",x"3ca7",x"3710",x"bb8c",x"354a",x"068d",x"3a5f",x"3a2d"),
(x"b85e",x"3c6a",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b865",x"3c6f",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b865",x"3c6f",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12"),
(x"b7c0",x"3c94",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b794",x"3c96",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b794",x"3c96",x"3710",x"b358",x"3bc9",x"0000",x"3bd9",x"39c8"),
(x"b50c",x"3c81",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b526",x"3c80",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b526",x"3c80",x"3710",x"33bc",x"bbc3",x"0000",x"3b06",x"3a0f"),
(x"b413",x"3ca7",x"36da",x"ba12",x"3935",x"8000",x"3a54",x"3a2d",x"b40b",x"3ca8",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b40b",x"3ca8",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e"),
(x"b84a",x"3c68",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b85e",x"3c6a",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b85e",x"3c6a",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d"),
(x"b794",x"3c96",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b77a",x"3c99",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b77a",x"3c99",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2"),
(x"b441",x"3c80",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b451",x"3c81",x"36da",x"a0dd",x"bc00",x"0000",x"3afb",x"39e7",x"b451",x"3c81",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7"),
(x"b40b",x"3ca8",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b3f4",x"3ca8",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3f4",x"3ca8",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32"),
(x"b83a",x"3c6b",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b84a",x"3c68",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b84a",x"3c68",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05"),
(x"b77a",x"3c99",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b776",x"3c9c",x"36da",x"bbce",x"b2fc",x"0000",x"3be3",x"39c0",x"b776",x"3c9c",x"3710",x"bbee",x"3037",x"0000",x"3bd9",x"39c0"),
(x"b451",x"3c81",x"36da",x"a0dd",x"bc00",x"0000",x"3afb",x"39e7",x"b50c",x"3c81",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b50c",x"3c81",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a"),
(x"b3f4",x"3ca8",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3d2",x"3ca7",x"36da",x"abf9",x"3bfc",x"0000",x"3a54",x"3a35",x"b3d2",x"3ca7",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35"),
(x"b569",x"3c72",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b568",x"3c75",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b568",x"3c75",x"3710",x"bb03",x"b7b2",x"868d",x"3a87",x"3b59"),
(x"b776",x"3c9c",x"36da",x"bbce",x"b2fc",x"0000",x"3be3",x"39c0",x"b77b",x"3c9e",x"36da",x"b853",x"baba",x"0000",x"3be3",x"39be",x"b77b",x"3c9e",x"3710",x"b937",x"ba10",x"8000",x"3bd9",x"39be"),
(x"b40d",x"3c78",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b441",x"3c80",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b441",x"3c80",x"3710",x"b7a3",x"bb07",x"0000",x"3b06",x"39e4"),
(x"b3d2",x"3ca7",x"36da",x"abf9",x"3bfc",x"0000",x"3a54",x"3a35",x"b3a5",x"3ca8",x"36da",x"32b5",x"3bd2",x"068d",x"3a54",x"3a39",x"b3a5",x"3ca8",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39"),
(x"b820",x"3c79",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b83a",x"3c6b",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b83a",x"3c6b",x"3710",x"3953",x"b9f7",x"0000",x"3a85",x"39ff"),
(x"b77b",x"3c9e",x"36da",x"b853",x"baba",x"0000",x"3a7d",x"3ac5",x"b790",x"3ca0",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b790",x"3ca0",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9"),
(x"b407",x"3c76",x"36da",x"bb61",x"b62a",x"0000",x"3afb",x"39d6",x"b40d",x"3c78",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b40d",x"3c78",x"3710",x"b8bf",x"ba70",x"868d",x"3b06",x"39d8"),
(x"b3a5",x"3ca8",x"36da",x"32b5",x"3bd2",x"068d",x"3a54",x"3a39",x"b368",x"3ca5",x"36da",x"3912",x"3a2f",x"068d",x"3a54",x"3a40",x"b368",x"3ca5",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40"),
(x"b575",x"3c70",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b569",x"3c72",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b569",x"3c72",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57"),
(x"b790",x"3ca0",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b7a8",x"3ca1",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7a8",x"3ca1",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace"),
(x"b409",x"3c75",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b407",x"3c76",x"36da",x"bb61",x"b62a",x"0000",x"3afb",x"39d6",x"b407",x"3c76",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6"),
(x"b368",x"3ca5",x"36da",x"3912",x"3a2f",x"068d",x"3a54",x"3a40",x"b340",x"3c9f",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b340",x"3c9f",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45"),
(x"b801",x"3c80",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b820",x"3c79",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b820",x"3c79",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1"),
(x"b7a8",x"3ca1",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7bd",x"3ca4",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7bd",x"3ca4",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2"),
(x"b413",x"3c71",x"36da",x"bb08",x"37a1",x"8000",x"3afb",x"39d2",x"b409",x"3c75",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b409",x"3c75",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5"),
(x"b340",x"3c9f",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b33a",x"3c9a",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b33a",x"3c9a",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49"),
(x"b7c0",x"3c82",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b801",x"3c80",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b801",x"3c80",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4"),
(x"b7bd",x"3ca4",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7c7",x"3ca6",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"3ca6",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5"),
(x"b931",x"3c69",x"36da",x"bbff",x"26b5",x"0000",x"39f5",x"33fa",x"b930",x"3c7f",x"36da",x"bbff",x"26b5",x"0000",x"3a09",x"33f0",x"b930",x"3c7f",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0"),
(x"b413",x"3c6f",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"3c71",x"36da",x"bb08",x"37a1",x"8000",x"3afb",x"39d2",x"b413",x"3c71",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2"),
(x"b33a",x"3c9a",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b351",x"3c95",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b351",x"3c95",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d"),
(x"b794",x"3c80",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b7c0",x"3c82",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b7c0",x"3c82",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7"),
(x"b7c7",x"3ca6",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"3ca7",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7c7",x"3ca7",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6"),
(x"b40b",x"3c6e",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b413",x"3c6f",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"3c6f",x"3710",x"ba12",x"b935",x"0000",x"3b06",x"39d0"),
(x"b351",x"3c95",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b34f",x"3c93",x"36da",x"3448",x"3bb5",x"0000",x"3a54",x"3a4f",x"b34f",x"3c93",x"3710",x"3913",x"3a2f",x"0000",x"3a5f",x"3a4f"),
(x"b77a",x"3c7d",x"36da",x"b83f",x"bac7",x"0000",x"3a7b",x"39c9",x"b794",x"3c80",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b794",x"3c80",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf"),
(x"b7c7",x"3ca7",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7a4",x"3cab",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b7a4",x"3cab",x"3710",x"b654",x"3b58",x"0000",x"3a87",x"3add"),
(x"b3f4",x"3c6e",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b40b",x"3c6e",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b40b",x"3c6e",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce"),
(x"b34f",x"3c93",x"36da",x"3448",x"3bb5",x"0000",x"3a6e",x"3b35",x"b326",x"3c93",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b326",x"3c93",x"3710",x"a5e9",x"3bff",x"0000",x"3a79",x"3b39"),
(x"b776",x"3c7b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b77a",x"3c7d",x"36da",x"b83f",x"bac7",x"0000",x"3a8a",x"3a50",x"b77a",x"3c7d",x"3710",x"b97c",x"b9d2",x"0000",x"3a95",x"3a50"),
(x"b7a4",x"3cab",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b783",x"3cae",x"36da",x"afa0",x"3bf1",x"8000",x"3a7d",x"3ae4",x"b783",x"3cae",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4"),
(x"b3d2",x"3c70",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3f4",x"3c6e",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b3f4",x"3c6e",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb"),
(x"b326",x"3c93",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b2d6",x"3c94",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2d6",x"3c94",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41"),
(x"b77b",x"3c79",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b776",x"3c7b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b776",x"3c7b",x"3710",x"bbce",x"32fb",x"0000",x"3a95",x"3a4d"),
(x"b783",x"3cae",x"36da",x"afa0",x"3bf1",x"8000",x"3a7d",x"3ae4",x"b73e",x"3caf",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b73e",x"3caf",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1"),
(x"b3a5",x"3c6e",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3d2",x"3c70",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3d2",x"3c70",x"3710",x"abf9",x"bbfc",x"0000",x"3b06",x"39c8"),
(x"b2d6",x"3c94",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2aa",x"3c97",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b2aa",x"3c97",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46"),
(x"b790",x"3c76",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b77b",x"3c79",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b77b",x"3c79",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c"),
(x"b73e",x"3caf",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b705",x"3cac",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b705",x"3cac",x"3710",x"34b8",x"3ba4",x"0000",x"3a87",x"3afc"),
(x"b368",x"3c71",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b3a5",x"3c6e",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3a5",x"3c6e",x"3710",x"32b5",x"bbd2",x"8000",x"3b06",x"39c3"),
(x"b2aa",x"3c97",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b261",x"3c9c",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b261",x"3c9c",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e"),
(x"b7a8",x"3c75",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b790",x"3c76",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b790",x"3c76",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47"),
(x"b705",x"3cac",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b6f1",x"3ca8",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6f1",x"3ca8",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01"),
(x"b340",x"3c77",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b368",x"3c71",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b368",x"3c71",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd"),
(x"b261",x"3c9c",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b22d",x"3c9e",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b22d",x"3c9e",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53"),
(x"b7bd",x"3c73",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7a8",x"3c75",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b7a8",x"3c75",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43"),
(x"b6f1",x"3ca8",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6ef",x"3ca2",x"36da",x"3b57",x"b658",x"8000",x"3a7d",x"3b05",x"b6ef",x"3ca2",x"3710",x"3be9",x"b0b7",x"868d",x"3a87",x"3b05"),
(x"b33a",x"3c7c",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b340",x"3c77",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b340",x"3c77",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7"),
(x"b22d",x"3c9e",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b1fd",x"3c9d",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1fd",x"3c9d",x"3710",x"35da",x"3b72",x"8000",x"3a79",x"3b57"),
(x"b7c7",x"3c71",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7bd",x"3c73",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7bd",x"3c73",x"3710",x"b821",x"3ada",x"0000",x"3a95",x"3a3e"),
(x"b6ef",x"3ca2",x"36da",x"3b57",x"b658",x"8000",x"3a7d",x"3b05",x"b6fb",x"3c9f",x"36da",x"37ed",x"baf2",x"068d",x"3a7d",x"3b08",x"b6fb",x"3c9f",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08"),
(x"b351",x"3c81",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b33a",x"3c7c",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b33a",x"3c7c",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3"),
(x"b1fd",x"3c9d",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1c1",x"3c98",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1c1",x"3c98",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e"),
(x"b7c7",x"3c6f",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"3c71",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7c7",x"3c71",x"3710",x"bb43",x"36b4",x"0000",x"3a95",x"3a3c"),
(x"b6fb",x"3c9f",x"36da",x"37ed",x"baf2",x"068d",x"3a7d",x"3b08",x"b721",x"3c9a",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b721",x"3c9a",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10"),
(x"b34f",x"3c83",x"36da",x"3913",x"ba2f",x"8000",x"3afb",x"39ae",x"b351",x"3c81",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b351",x"3c81",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af"),
(x"b1c1",x"3c98",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1a1",x"3c97",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b1a1",x"3c97",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61"),
(x"b7a4",x"3c6c",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7c7",x"3c6f",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"3c6f",x"3710",x"b744",x"bb20",x"0000",x"3a95",x"3a3b"),
(x"b721",x"3c9a",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b72e",x"3c98",x"36da",x"3b4f",x"b67e",x"0000",x"3a7d",x"3b13",x"b72e",x"3c98",x"3710",x"39a7",x"b9a8",x"0000",x"3a87",x"3b13"),
(x"b326",x"3c83",x"36da",x"a5e9",x"bbff",x"0000",x"3a6e",x"3bae",x"b34f",x"3c83",x"36da",x"3913",x"ba2f",x"8000",x"3a6e",x"3bb2",x"b34f",x"3c83",x"3710",x"3448",x"bbb5",x"0000",x"3a79",x"3bb2"),
(x"b1a1",x"3c97",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b161",x"3c96",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b161",x"3c96",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67"),
(x"b783",x"3c68",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b7a4",x"3c6c",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7a4",x"3c6c",x"3710",x"b64a",x"bb5a",x"0000",x"3a95",x"3a34"),
(x"b72e",x"3c98",x"36da",x"3b4f",x"b67e",x"0000",x"3a97",x"39c6",x"b72d",x"3c96",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b72d",x"3c96",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8"),
(x"b2d6",x"3c82",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b326",x"3c83",x"36da",x"a5e9",x"bbff",x"0000",x"3a6e",x"3bae",x"b326",x"3c83",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae"),
(x"b161",x"3c96",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b135",x"3c94",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b135",x"3c94",x"3710",x"3822",x"3ad9",x"868d",x"3a79",x"3b6c"),
(x"b73e",x"3c67",x"36da",x"27ae",x"bbff",x"8000",x"3a8a",x"3a20",x"b783",x"3c68",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b783",x"3c68",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d"),
(x"b72d",x"3c96",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b721",x"3c95",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b721",x"3c95",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca"),
(x"b2aa",x"3c7f",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2d6",x"3c82",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b2d6",x"3c82",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6"),
(x"b135",x"3c94",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b116",x"3c8f",x"36da",x"3bdf",x"31b0",x"868d",x"3a6e",x"3b70",x"b116",x"3c8f",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70"),
(x"b705",x"3c6a",x"36da",x"34b8",x"bba4",x"8000",x"3a8a",x"3a15",x"b73e",x"3c67",x"36da",x"27ae",x"bbff",x"8000",x"3a8a",x"3a20",x"b73e",x"3c67",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20"),
(x"b575",x"3ca9",x"36da",x"bab5",x"385c",x"8a8d",x"3a97",x"3a28",x"b568",x"3cad",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b568",x"3cad",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b"),
(x"b938",x"3c81",x"36da",x"bbfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"b93a",x"3c96",x"36da",x"bbfe",x"a8f0",x"0000",x"3be9",x"39cf",x"b93a",x"3c96",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3be8",x"39da"),
(x"b261",x"3c7a",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b2aa",x"3c7f",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2aa",x"3c7f",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2"),
(x"b931",x"3cae",x"36da",x"23ae",x"3bff",x"0000",x"3be3",x"3a63",x"b8ff",x"3cae",x"36da",x"26a1",x"3bff",x"8000",x"3be3",x"3a4f",x"b8ff",x"3cae",x"3710",x"257a",x"3bff",x"15bc",x"3bd9",x"3a4f"),
(x"b6f1",x"3c6f",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b705",x"3c6a",x"36da",x"34b8",x"bba4",x"8000",x"3a8a",x"3a15",x"b705",x"3c6a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15"),
(x"b721",x"3c95",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b669",x"3c96",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b669",x"3c96",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed"),
(x"b22d",x"3c78",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b261",x"3c7a",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b261",x"3c7a",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a"),
(x"b6ef",x"3c74",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6f1",x"3c6f",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b6f1",x"3c6f",x"3710",x"3b73",x"b5d3",x"8000",x"3a95",x"3a10"),
(x"b669",x"3c96",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b63d",x"3c97",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b63d",x"3c97",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5"),
(x"b930",x"3c7f",x"36da",x"b67a",x"bb50",x"0000",x"3bc0",x"3984",x"b938",x"3c81",x"36da",x"b67a",x"bb50",x"0000",x"3bbd",x"3982",x"b938",x"3c81",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a"),
(x"a379",x"39c2",x"36eb",x"bba3",x"b453",x"2fdf",x"392c",x"31f8",x"a271",x"39c2",x"3718",x"bbb8",x"b22d",x"31b0",x"3921",x"31e9",x"a1bd",x"39b8",x"3715",x"bbf4",x"2da3",x"2b3e",x"3920",x"31fe"),
(x"a379",x"39c2",x"36eb",x"bba3",x"b453",x"2fdf",x"392c",x"31f8",x"a3d0",x"39d2",x"36eb",x"bb7a",x"3531",x"30a8",x"392e",x"31d7",x"a303",x"39d2",x"3715",x"bbda",x"2e4f",x"312f",x"3924",x"31c9"),
(x"a3d0",x"39d2",x"36eb",x"bb7a",x"3531",x"30a8",x"392e",x"31d7",x"a133",x"39e5",x"36eb",x"b8c7",x"3a49",x"310c",x"3931",x"31aa",x"a0f3",x"39e1",x"3714",x"ba0a",x"3915",x"3126",x"3926",x"31a6"),
(x"a133",x"39e5",x"36eb",x"b8c7",x"3a49",x"310c",x"3931",x"31aa",x"9725",x"39ec",x"36eb",x"a3ae",x"3bec",x"3065",x"3932",x"3182",x"96c5",x"39e9",x"3714",x"b236",x"3bc0",x"30e0",x"3927",x"317f"),
(x"9725",x"39ec",x"36eb",x"a3ae",x"3bec",x"3065",x"3932",x"3182",x"22b9",x"39e9",x"36eb",x"36e0",x"3b1c",x"3118",x"3933",x"3141",x"21e6",x"39e6",x"3714",x"335f",x"3baf",x"30fd",x"3928",x"3145"),
(x"22b9",x"39e9",x"36eb",x"36e0",x"3b1c",x"3118",x"3933",x"3141",x"2505",x"39db",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3932",x"3119",x"24a4",x"39db",x"3715",x"3a37",x"38de",x"311d",x"3928",x"311f"),
(x"2505",x"39db",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3932",x"3119",x"256c",x"39cc",x"36eb",x"3bf7",x"2138",x"2dcf",x"3931",x"30f7",x"252e",x"39cc",x"3715",x"3bf2",x"2495",x"2f43",x"3926",x"30fd"),
(x"250e",x"39be",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"3930",x"30d9",x"24bc",x"39be",x"3715",x"3b87",x"b537",x"2d81",x"3925",x"30e0",x"252e",x"39cc",x"3715",x"3bf2",x"2495",x"2f43",x"3926",x"30fd"),
(x"2470",x"39b4",x"36eb",x"3bfd",x"212b",x"29e6",x"392f",x"30c2",x"2464",x"39b5",x"3717",x"3bff",x"2481",x"2487",x"3924",x"30cb",x"24bc",x"39be",x"3715",x"3b87",x"b537",x"2d81",x"3925",x"30e0"),
(x"250d",x"3981",x"36eb",x"3b9b",x"34d2",x"2ca7",x"392a",x"3055",x"25ec",x"397f",x"36eb",x"3b76",x"3593",x"2dee",x"3929",x"3046",x"25c0",x"397d",x"3714",x"3b74",x"35a7",x"2d5e",x"391f",x"304d"),
(x"2066",x"39b7",x"36eb",x"bbf7",x"9e8d",x"2dbc",x"38cc",x"30e5",x"2019",x"39c2",x"36eb",x"bbab",x"33f1",x"3064",x"38cc",x"30fc",x"20c8",x"39c0",x"3716",x"bbb5",x"33c6",x"2f0a",x"38d7",x"30f8"),
(x"2029",x"3983",x"36eb",x"ba79",x"3840",x"3401",x"38cb",x"3076",x"2066",x"39b7",x"36eb",x"bbf7",x"9e8d",x"2dbc",x"38cc",x"30e5",x"20e0",x"39b7",x"3718",x"bbf1",x"95bc",x"2fb4",x"38d7",x"30e3"),
(x"a50e",x"3969",x"36eb",x"b409",x"bbbc",x"27db",x"3918",x"32b5",x"a4fc",x"3981",x"36eb",x"bbc6",x"328d",x"2f71",x"391c",x"3288",x"a4b5",x"397f",x"3715",x"bbb4",x"33e8",x"2ed7",x"3913",x"3278"),
(x"262b",x"3969",x"36eb",x"36d0",x"bb39",x"2ab1",x"3927",x"3019",x"25f4",x"396a",x"3714",x"2f03",x"bbf3",x"23ef",x"391d",x"3024",x"25c0",x"397d",x"3714",x"3b74",x"35a7",x"2d5e",x"391f",x"304d"),
(x"9909",x"39bf",x"3715",x"3b88",x"3531",x"2dc2",x"38d8",x"319c",x"95ed",x"39c0",x"36ee",x"3b70",x"358e",x"2fc0",x"38ce",x"319b",x"9651",x"39b8",x"36eb",x"3bd3",x"b208",x"2da6",x"38ce",x"31ae"),
(x"9caa",x"39c8",x"36ee",x"3b20",x"3725",x"2d51",x"38ce",x"3187",x"95ed",x"39c0",x"36ee",x"3b70",x"358e",x"2fc0",x"38ce",x"319b",x"9909",x"39bf",x"3715",x"3b88",x"3531",x"2dc2",x"38d8",x"319c"),
(x"9cff",x"39d0",x"36ee",x"3b1d",x"b747",x"2911",x"38ce",x"3174",x"9caa",x"39c8",x"36ee",x"3b20",x"3725",x"2d51",x"38ce",x"3187",x"9db7",x"39ca",x"3717",x"3bd6",x"323b",x"2a8a",x"38d9",x"3181"),
(x"216b",x"39cf",x"36ee",x"ba3f",x"b8f6",x"2c87",x"38ce",x"3120",x"1f13",x"39d8",x"36ee",x"b233",x"bbd8",x"a538",x"38ce",x"3139",x"1f52",x"39d7",x"3715",x"b67e",x"bb4e",x"2839",x"38d7",x"3137"),
(x"9fcf",x"3985",x"36eb",x"3be6",x"2cac",x"3077",x"38d0",x"321f",x"a069",x"397e",x"3718",x"398b",x"396b",x"33db",x"38db",x"3229",x"993e",x"39b7",x"3716",x"3bce",x"b2bb",x"2b41",x"38d9",x"31ad"),
(x"9909",x"39bf",x"3715",x"28d3",x"a80e",x"3bfd",x"3968",x"32c8",x"993e",x"39b7",x"3716",x"a82f",x"2808",x"3bfd",x"3967",x"32be",x"a1bd",x"39b8",x"3715",x"a1ae",x"23fc",x"3bff",x"3963",x"32c0"),
(x"9db7",x"39ca",x"3717",x"250b",x"281b",x"3bfe",x"3966",x"32d5",x"9909",x"39bf",x"3715",x"28d3",x"a80e",x"3bfd",x"3968",x"32c8",x"a271",x"39c2",x"3718",x"28fa",x"a4f7",x"3bfe",x"3962",x"32cc"),
(x"9cfd",x"39d2",x"3716",x"252b",x"2c98",x"3bfa",x"3966",x"32df",x"9db7",x"39ca",x"3717",x"250b",x"281b",x"3bfe",x"3966",x"32d5",x"a303",x"39d2",x"3715",x"9ea7",x"2bd8",x"3bfc",x"3961",x"32de"),
(x"94d9",x"39d7",x"3713",x"1818",x"9cd0",x"3c00",x"3968",x"32e4",x"9cfd",x"39d2",x"3716",x"252b",x"2c98",x"3bfa",x"3966",x"32df",x"a0f3",x"39e1",x"3714",x"263f",x"27c1",x"3bfe",x"3963",x"32f0"),
(x"1f52",x"39d7",x"3715",x"9cd0",x"191e",x"3c00",x"396d",x"32e6",x"94d9",x"39d7",x"3713",x"1818",x"9cd0",x"3c00",x"3968",x"32e4",x"96c5",x"39e9",x"3714",x"a194",x"a0d0",x"3bff",x"3968",x"32f9"),
(x"21f4",x"39d0",x"3714",x"9dbc",x"252b",x"3bff",x"3970",x"32dc",x"1f52",x"39d7",x"3715",x"9cd0",x"191e",x"3c00",x"396d",x"32e6",x"21e6",x"39e6",x"3714",x"1dd6",x"247a",x"3bff",x"3970",x"32f6"),
(x"21f4",x"39d0",x"3714",x"9dbc",x"252b",x"3bff",x"3970",x"32dc",x"24a4",x"39db",x"3715",x"a793",x"184d",x"3bff",x"3973",x"32e9",x"252e",x"39cc",x"3715",x"9818",x"26bb",x"3bff",x"3975",x"32d7"),
(x"2211",x"39c9",x"3716",x"2338",x"267a",x"3bff",x"3970",x"32d4",x"252e",x"39cc",x"3715",x"9818",x"26bb",x"3bff",x"3975",x"32d7",x"24bc",x"39be",x"3715",x"264c",x"29dc",x"3bfd",x"3974",x"32c7"),
(x"20e0",x"39b7",x"3718",x"2793",x"2439",x"3bfe",x"396e",x"32be",x"20c8",x"39c0",x"3716",x"24b5",x"2b17",x"3bfc",x"396e",x"32ca",x"24bc",x"39be",x"3715",x"264c",x"29dc",x"3bfd",x"3974",x"32c7"),
(x"24de",x"3981",x"3717",x"2984",x"a0c2",x"3bfd",x"3974",x"327f",x"2116",x"397d",x"3718",x"23ae",x"ac2f",x"3bfb",x"396f",x"327a",x"20e0",x"39b7",x"3718",x"2793",x"2439",x"3bfe",x"396e",x"32be"),
(x"219d",x"39c9",x"36ee",x"bb83",x"3534",x"2f10",x"38cd",x"3111",x"216b",x"39cf",x"36ee",x"ba3f",x"b8f6",x"2c87",x"38ce",x"3120",x"21f4",x"39d0",x"3714",x"bb20",x"b711",x"2eb1",x"38d7",x"311c"),
(x"a46c",x"3981",x"36eb",x"bbaa",x"3475",x"2c25",x"391d",x"327f",x"a165",x"39b8",x"36eb",x"bbf4",x"2d6d",x"ac2d",x"3929",x"3212",x"a1bd",x"39b8",x"3715",x"bbf4",x"2da3",x"2b3e",x"3920",x"31fe"),
(x"a46c",x"3981",x"36eb",x"bbaa",x"3475",x"2c25",x"391d",x"327f",x"a3f1",x"3980",x"3718",x"bba4",x"33dc",x"313d",x"3913",x"326a",x"a4b5",x"397f",x"3715",x"bbb4",x"33e8",x"2ed7",x"3913",x"3278"),
(x"2116",x"397d",x"3718",x"23ae",x"ac2f",x"3bfb",x"396f",x"327a",x"25f4",x"396a",x"3714",x"273e",x"ad9b",x"3bf7",x"3976",x"3263",x"a4d5",x"3969",x"3715",x"a081",x"ad9e",x"3bf8",x"395e",x"3263"),
(x"94d9",x"39d7",x"3713",x"33d9",x"bbc1",x"a386",x"38d7",x"315c",x"9548",x"39d8",x"36ee",x"348f",x"bba6",x"ac10",x"38ce",x"315d",x"9cff",x"39d0",x"36ee",x"3b1d",x"b747",x"2911",x"38ce",x"3174"),
(x"2470",x"39b4",x"36eb",x"3bfd",x"212b",x"29e6",x"392f",x"30c2",x"250d",x"3981",x"36eb",x"3b9b",x"34d2",x"2ca7",x"392a",x"3055",x"24de",x"3981",x"3717",x"3be8",x"30a2",x"2973",x"391f",x"305e"),
(x"1f13",x"39d8",x"36ee",x"b233",x"bbd8",x"a538",x"38ce",x"3139",x"9548",x"39d8",x"36ee",x"348f",x"bba6",x"ac10",x"38ce",x"315d",x"94d9",x"39d7",x"3713",x"33d9",x"bbc1",x"a386",x"38d7",x"315c"),
(x"2029",x"3983",x"36eb",x"ba79",x"3840",x"3401",x"38cb",x"3261",x"2116",x"397d",x"3718",x"ba6d",x"3838",x"3468",x"38d6",x"3278",x"a069",x"397e",x"3718",x"398b",x"396b",x"33db",x"38db",x"3229"),
(x"a50e",x"3969",x"36eb",x"b409",x"bbbc",x"27db",x"3918",x"2ec7",x"a4d5",x"3969",x"3715",x"b3c8",x"bbc2",x"236c",x"390e",x"2eed",x"25f4",x"396a",x"3714",x"2f03",x"bbf3",x"23ef",x"391d",x"3024"),
(x"20c8",x"39c0",x"3716",x"bbb5",x"33c6",x"2f0a",x"38d7",x"30f8",x"2019",x"39c2",x"36eb",x"bbab",x"33f1",x"3064",x"38cc",x"30fc",x"219d",x"39c9",x"36ee",x"bb83",x"3534",x"2f10",x"38cd",x"3111"),
(x"91f4",x"3ba1",x"3716",x"30f9",x"a8b2",x"3be5",x"3b4b",x"3b05",x"1aac",x"3ba1",x"3712",x"342b",x"2e69",x"3bae",x"3b48",x"3b06",x"20f7",x"3b90",x"370e",x"2fd2",x"2717",x"3bef",x"3b44",x"3b0d"),
(x"a03c",x"3b86",x"36eb",x"bb99",x"3315",x"330d",x"3982",x"302f",x"980d",x"3ba6",x"36eb",x"b996",x"395f",x"33ec",x"3983",x"300b",x"91f4",x"3ba1",x"3716",x"badd",x"375a",x"334d",x"397d",x"300e"),
(x"8010",x"3b06",x"3714",x"ac39",x"29a5",x"3bf9",x"3b50",x"3b47",x"a040",x"3b03",x"3713",x"a91b",x"2b55",x"3bfb",x"3b57",x"3b48",x"9d28",x"3b16",x"3712",x"aa69",x"287e",x"3bfc",x"3b54",x"3b40"),
(x"a34c",x"3b12",x"3711",x"a481",x"2546",x"3bff",x"3b5b",x"3b42",x"a20d",x"3b19",x"3712",x"2a38",x"ad35",x"3bf6",x"3b59",x"3b3f",x"9ff6",x"3b1a",x"3711",x"a994",x"2977",x"3bfc",x"3b56",x"3b3e"),
(x"9d28",x"3b16",x"3712",x"aa69",x"287e",x"3bfc",x"3b54",x"3b40",x"a040",x"3b03",x"3713",x"a91b",x"2b55",x"3bfb",x"3b57",x"3b48",x"a273",x"3b06",x"3712",x"aa73",x"2a97",x"3bfa",x"3b5a",x"3b47"),
(x"9c36",x"3afd",x"3718",x"ae36",x"a153",x"3bf6",x"3b53",x"3b4b",x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f",x"a17b",x"3afb",x"3711",x"afec",x"ac2c",x"3beb",x"3b59",x"3b4b"),
(x"a035",x"3acc",x"3713",x"ae9c",x"3366",x"3bbd",x"3b58",x"3b60",x"a289",x"3acf",x"370f",x"9df0",x"a631",x"3bff",x"3b5c",x"3b5e",x"9c56",x"3adb",x"370e",x"26d5",x"25c2",x"3bfe",x"3b54",x"3b5a"),
(x"9f72",x"3ae4",x"3713",x"a538",x"ac7a",x"3bfa",x"3b57",x"3b56",x"9c56",x"3adb",x"370e",x"26d5",x"25c2",x"3bfe",x"3b54",x"3b5a",x"a289",x"3acf",x"370f",x"9df0",x"a631",x"3bff",x"3b5c",x"3b5e"),
(x"a407",x"3aeb",x"370f",x"aec5",x"1a24",x"3bf4",x"3b5d",x"3b52",x"9f87",x"3ae7",x"3713",x"a7e9",x"2846",x"3bfd",x"3b57",x"3b54",x"9f72",x"3ae4",x"3713",x"a538",x"ac7a",x"3bfa",x"3b57",x"3b56"),
(x"9f87",x"3ae7",x"3713",x"a7e9",x"2846",x"3bfd",x"3b57",x"3b54",x"a407",x"3aeb",x"370f",x"aec5",x"1a24",x"3bf4",x"3b5d",x"3b52",x"a17b",x"3afb",x"3711",x"afec",x"ac2c",x"3beb",x"3b59",x"3b4b"),
(x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f",x"9476",x"3aef",x"3713",x"25bc",x"b7de",x"3af6",x"3b51",x"3b51",x"9d1a",x"3aec",x"3710",x"ac5b",x"b0a5",x"3be5",x"3b55",x"3b52"),
(x"9d1a",x"3aec",x"3710",x"ac5b",x"b0a5",x"3be5",x"3b55",x"3b52",x"9f87",x"3ae7",x"3713",x"a7e9",x"2846",x"3bfd",x"3b57",x"3b54",x"a17b",x"3afb",x"3711",x"afec",x"ac2c",x"3beb",x"3b59",x"3b4b"),
(x"1e77",x"3a8d",x"3715",x"a6c2",x"ac65",x"3bfa",x"3b4b",x"3b7b",x"990c",x"3a8d",x"3712",x"af67",x"a981",x"3bf0",x"3b52",x"3b7b",x"19fe",x"3a9c",x"3717",x"aff2",x"aa7a",x"3bed",x"3b4e",x"3b74"),
(x"a38f",x"3aa2",x"3712",x"b163",x"a345",x"3be2",x"3b5c",x"3b72",x"a2d9",x"3aab",x"3714",x"a860",x"af8b",x"3bf0",x"3b5b",x"3b6e",x"a13d",x"3aae",x"3716",x"acd8",x"a7e2",x"3bf9",x"3b58",x"3b6d"),
(x"9e62",x"3aad",x"3716",x"2818",x"ad02",x"3bf8",x"3b55",x"3b6d",x"9d1e",x"3a94",x"3711",x"240b",x"ad5c",x"3bf8",x"3b54",x"3b78",x"a2cb",x"3a9a",x"3714",x"1553",x"ab62",x"3bfc",x"3b5b",x"3b75"),
(x"9d1e",x"3a94",x"3711",x"240b",x"ad5c",x"3bf8",x"3b54",x"3b78",x"987a",x"3aa6",x"3714",x"a4f7",x"ada9",x"3bf7",x"3b52",x"3b70",x"0e53",x"3aa0",x"3714",x"b036",x"a73e",x"3bed",x"3b50",x"3b73"),
(x"19fe",x"3a9c",x"3717",x"aff2",x"aa7a",x"3bed",x"3b4e",x"3b74",x"990c",x"3a8d",x"3712",x"af67",x"a981",x"3bf0",x"3b52",x"3b7b",x"9a71",x"3a91",x"3711",x"b27d",x"175f",x"3bd5",x"3b53",x"3b79"),
(x"9a71",x"3a91",x"3711",x"b27d",x"175f",x"3bd5",x"3b53",x"3b79",x"9d1e",x"3a94",x"3711",x"240b",x"ad5c",x"3bf8",x"3b54",x"3b78",x"0e53",x"3aa0",x"3714",x"b036",x"a73e",x"3bed",x"3b50",x"3b73"),
(x"9ae8",x"3a82",x"3712",x"b146",x"2c91",x"3bde",x"3b53",x"3b7f",x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c"),
(x"1f1f",x"3a6b",x"3718",x"2138",x"ae95",x"3bf4",x"3b4b",x"3b89",x"21d8",x"3a6b",x"3719",x"a3bb",x"27c8",x"3bfe",x"3b47",x"3b89",x"21e0",x"3a69",x"3719",x"a90e",x"af00",x"3bf2",x"3b47",x"3b8a"),
(x"1e5a",x"3a6d",x"3718",x"2b4f",x"2525",x"3bfc",x"3b4c",x"3b89",x"1f1f",x"3a6b",x"3718",x"2138",x"ae95",x"3bf4",x"3b4b",x"3b89",x"8dee",x"3a63",x"3718",x"ae3b",x"1fae",x"3bf6",x"3b51",x"3b8c"),
(x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"20ca",x"3a73",x"3715",x"2d65",x"ac5a",x"3bf3",x"3b49",x"3b86",x"1e5a",x"3a6d",x"3718",x"2b4f",x"2525",x"3bfc",x"3b4c",x"3b89"),
(x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"2091",x"3a89",x"3717",x"2d2d",x"2ecb",x"3bed",x"3b49",x"3b7d",x"2288",x"3a7e",x"3718",x"2cf2",x"191e",x"3bf9",x"3b46",x"3b81"),
(x"22dc",x"3a86",x"3712",x"359c",x"336a",x"3b42",x"3b46",x"3b7e",x"2288",x"3a7e",x"3718",x"2cf2",x"191e",x"3bf9",x"3b46",x"3b81",x"2091",x"3a89",x"3717",x"2d2d",x"2ecb",x"3bed",x"3b49",x"3b7d"),
(x"1b8e",x"3a7c",x"3718",x"abb4",x"28d3",x"3bfa",x"3b4d",x"3b82",x"9ae8",x"3a82",x"3712",x"b146",x"2c91",x"3bde",x"3b53",x"3b7f",x"1f4b",x"3a8a",x"3716",x"b009",x"2da6",x"3be7",x"3b4b",x"3b7c"),
(x"1f4b",x"3a8a",x"3716",x"b009",x"2da6",x"3be7",x"3b4b",x"3b7c",x"9ae8",x"3a82",x"3712",x"b146",x"2c91",x"3bde",x"3b53",x"3b7f",x"990c",x"3a8d",x"3712",x"af67",x"a981",x"3bf0",x"3b52",x"3b7b"),
(x"1d4c",x"3a9f",x"3717",x"97c8",x"9f79",x"3c00",x"3b4c",x"3b73",x"2147",x"3a9a",x"3718",x"ac00",x"2911",x"3bfa",x"3b48",x"3b75",x"1f29",x"3a92",x"3714",x"a57a",x"ae8a",x"3bf4",x"3b4b",x"3b79"),
(x"1d4c",x"3a9f",x"3717",x"97c8",x"9f79",x"3c00",x"3b4c",x"3b73",x"20ef",x"3aa9",x"3715",x"a51e",x"2d06",x"3bf9",x"3b49",x"3b6f",x"2147",x"3a9a",x"3718",x"ac00",x"2911",x"3bfa",x"3b48",x"3b75"),
(x"20ef",x"3aa9",x"3715",x"a51e",x"2d06",x"3bf9",x"3b49",x"3b6f",x"2308",x"3ab8",x"3714",x"2dba",x"2266",x"3bf7",x"3b45",x"3b69",x"2442",x"3ab2",x"3714",x"175f",x"2c2c",x"3bfb",x"3b43",x"3b6b"),
(x"2308",x"3ab8",x"3714",x"2dba",x"2266",x"3bf7",x"3b45",x"3b69",x"2365",x"3ace",x"3715",x"3468",x"247a",x"3bb0",x"3b45",x"3b60",x"24cc",x"3acb",x"3712",x"3106",x"273e",x"3be5",x"3b41",x"3b61"),
(x"2365",x"3ace",x"3715",x"3468",x"247a",x"3bb0",x"3b45",x"3b60",x"22bc",x"3adf",x"3717",x"3273",x"2f43",x"3bc8",x"3b46",x"3b59",x"243c",x"3ae3",x"3710",x"3550",x"2e33",x"3b81",x"3b43",x"3b57"),
(x"22bc",x"3adf",x"3717",x"3273",x"2f43",x"3bc8",x"3b46",x"3b59",x"1f35",x"3aed",x"3711",x"ae24",x"2a2e",x"3bf4",x"3b4b",x"3b52",x"21ba",x"3af2",x"3712",x"2b5c",x"2345",x"3bfc",x"3b47",x"3b50"),
(x"1a19",x"3aef",x"3712",x"2dd2",x"b04b",x"3be4",x"3b4e",x"3b51",x"08f2",x"3afe",x"3716",x"2f4d",x"aa5f",x"3bf0",x"3b50",x"3b4b",x"21ba",x"3af2",x"3712",x"2b5c",x"2345",x"3bfc",x"3b47",x"3b50"),
(x"1a19",x"3aef",x"3712",x"2dd2",x"b04b",x"3be4",x"3b4e",x"3b51",x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f",x"08f2",x"3afe",x"3716",x"2f4d",x"aa5f",x"3bf0",x"3b50",x"3b4b"),
(x"1a19",x"3aef",x"3712",x"2dd2",x"b04b",x"3be4",x"3b4e",x"3b51",x"9476",x"3aef",x"3713",x"25bc",x"b7de",x"3af6",x"3b51",x"3b51",x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f"),
(x"08f2",x"3afe",x"3716",x"2f4d",x"aa5f",x"3bf0",x"3b50",x"3b4b",x"91dd",x"3af4",x"3718",x"ac13",x"b1c5",x"3bda",x"3b51",x"3b4f",x"9c36",x"3afd",x"3718",x"ae36",x"a153",x"3bf6",x"3b53",x"3b4b"),
(x"9e8d",x"3aff",x"3716",x"af15",x"329c",x"3bc7",x"3b55",x"3b4a",x"8010",x"3b06",x"3714",x"ac39",x"29a5",x"3bf9",x"3b50",x"3b47",x"9588",x"3b01",x"3716",x"a553",x"32c7",x"3bd1",x"3b51",x"3b49"),
(x"9e8d",x"3aff",x"3716",x"af15",x"329c",x"3bc7",x"3b55",x"3b4a",x"a040",x"3b03",x"3713",x"a91b",x"2b55",x"3bfb",x"3b57",x"3b48",x"8010",x"3b06",x"3714",x"ac39",x"29a5",x"3bf9",x"3b50",x"3b47"),
(x"9a85",x"3b15",x"3713",x"ada1",x"2f15",x"3beb",x"3b52",x"3b41",x"1820",x"3b1f",x"370f",x"aedc",x"2cd0",x"3bee",x"3b4e",x"3b3d",x"1f40",x"3b15",x"3717",x"b0e7",x"3057",x"3bd4",x"3b4a",x"3b41"),
(x"1820",x"3b1f",x"370f",x"aedc",x"2cd0",x"3bee",x"3b4e",x"3b3d",x"1d56",x"3b33",x"3716",x"aadf",x"a6b5",x"3bfc",x"3b4b",x"3b34",x"221f",x"3b30",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3b45",x"3b36"),
(x"2312",x"3b69",x"370d",x"3809",x"2e09",x"3add",x"3b41",x"3b1e",x"2386",x"3b62",x"370f",x"36c9",x"2fac",x"3b2e",x"3b41",x"3b21",x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c"),
(x"21a5",x"3b7a",x"3712",x"29f0",x"2b1d",x"3bfa",x"3b43",x"3b16",x"9cbb",x"3b6c",x"3715",x"19bc",x"a6cf",x"3bff",x"3b51",x"3b1b",x"9df1",x"3b85",x"3715",x"2d56",x"20d0",x"3bf8",x"3b50",x"3b10"),
(x"1882",x"3b48",x"370e",x"bb5f",x"b5f1",x"2f4d",x"397b",x"306f",x"1737",x"3b47",x"36eb",x"bb4a",x"b677",x"2cf9",x"397f",x"3074",x"9f02",x"3b6a",x"36eb",x"bb89",x"b473",x"31fc",x"3981",x"304c"),
(x"a175",x"3a2c",x"3710",x"3bfd",x"a997",x"a0a8",x"3bd5",x"3971",x"a0d2",x"3a3e",x"3713",x"3ba5",x"b497",x"ac28",x"3bd9",x"3971",x"a122",x"3a3e",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3bd9",x"396c"),
(x"a167",x"3a20",x"36eb",x"3bf5",x"2e59",x"2467",x"3bd2",x"396c",x"a140",x"3a1c",x"3714",x"3beb",x"308b",x"98b5",x"3bd1",x"3971",x"a175",x"3a2c",x"3710",x"3bfd",x"a997",x"a0a8",x"3bd5",x"3971"),
(x"9c3a",x"3a58",x"3714",x"3b1c",x"b754",x"223f",x"3be1",x"3971",x"8dee",x"3a63",x"3718",x"b9e5",x"b968",x"0000",x"3be4",x"3972",x"8dee",x"3a63",x"36eb",x"b46a",x"bb91",x"316a",x"3be4",x"396c"),
(x"a122",x"3a3e",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3bd9",x"396c",x"a0d2",x"3a3e",x"3713",x"3ba5",x"b497",x"ac28",x"3bd9",x"3971",x"9c3a",x"3a58",x"3714",x"3b1c",x"b754",x"223f",x"3be1",x"3971"),
(x"a099",x"3a14",x"3712",x"3b76",x"35c5",x"204d",x"3bce",x"3971",x"a140",x"3a1c",x"3714",x"3beb",x"308b",x"98b5",x"3bd1",x"3971",x"a167",x"3a20",x"36eb",x"3bf5",x"2e59",x"2467",x"3bd2",x"396c"),
(x"a051",x"3a11",x"36eb",x"3ab1",x"3862",x"21e3",x"3bcd",x"396c",x"9ecc",x"3a0d",x"3714",x"395a",x"39f1",x"2025",x"3bcc",x"3971",x"a099",x"3a14",x"3712",x"3b76",x"35c5",x"204d",x"3bce",x"3971"),
(x"9b3f",x"3a09",x"36eb",x"37e1",x"3af5",x"269a",x"3bca",x"396c",x"9aa8",x"3a08",x"3714",x"35bf",x"3b76",x"27db",x"3bca",x"3971",x"9ecc",x"3a0d",x"3714",x"395a",x"39f1",x"2025",x"3bcc",x"3971"),
(x"197e",x"3a06",x"36eb",x"303c",x"3beb",x"299b",x"3bc7",x"396c",x"1a1e",x"3a04",x"3715",x"a836",x"3bfd",x"294f",x"3bc6",x"3972",x"9aa8",x"3a08",x"3714",x"35bf",x"3b76",x"27db",x"3bca",x"3971"),
(x"20a0",x"3a08",x"36eb",x"b868",x"3aab",x"296a",x"3bc3",x"396c",x"20b2",x"3a07",x"3716",x"b86f",x"3aa7",x"2604",x"3bc3",x"3972",x"1a1e",x"3a04",x"3715",x"a836",x"3bfd",x"294f",x"3bc6",x"3972"),
(x"20a0",x"3a08",x"36eb",x"b868",x"3aab",x"296a",x"3bc3",x"396c",x"2300",x"3a14",x"36eb",x"baf3",x"37df",x"2b38",x"3bbf",x"396c",x"2335",x"3a14",x"3714",x"bb01",x"37b5",x"2839",x"3bbf",x"3971"),
(x"23d0",x"3a1e",x"36eb",x"bbf9",x"2d11",x"2511",x"3bbc",x"396c",x"23d3",x"3a1f",x"3714",x"bbe6",x"b10f",x"9bfc",x"3bbc",x"3971",x"2335",x"3a14",x"3714",x"bb01",x"37b5",x"2839",x"3bbf",x"3971"),
(x"2300",x"3a28",x"36eb",x"b90c",x"ba34",x"2532",x"3bba",x"396c",x"22d3",x"3a28",x"3715",x"b928",x"ba1d",x"1553",x"3bb9",x"3971",x"23d3",x"3a1f",x"3714",x"bbe6",x"b10f",x"9bfc",x"3bbc",x"3971"),
(x"2300",x"3a28",x"36eb",x"b90c",x"ba34",x"2532",x"3b61",x"39ee",x"20b2",x"3a28",x"36eb",x"35dd",x"bb6d",x"2be9",x"3b64",x"39ee",x"20d5",x"3a29",x"3714",x"2fe4",x"bbee",x"28fd",x"3b64",x"39e9"),
(x"20b2",x"3a28",x"36eb",x"35dd",x"bb6d",x"2be9",x"3b64",x"39ee",x"1ead",x"3a23",x"36eb",x"32b1",x"bbc8",x"2e54",x"3b66",x"39ef",x"1e4f",x"3a25",x"3711",x"364f",x"bb52",x"2d1b",x"3b66",x"39ea"),
(x"13e1",x"3a42",x"36eb",x"bbf6",x"2a70",x"2d61",x"3b72",x"39ef",x"15a0",x"3a42",x"3713",x"bbc2",x"33a5",x"298a",x"3b71",x"39ea",x"3d81",x"3a3e",x"3711",x"ba7a",x"38b0",x"283c",x"3b70",x"39ea"),
(x"1ead",x"3a23",x"36eb",x"32b1",x"bbc8",x"2e54",x"3b66",x"39ef",x"0f13",x"3a23",x"36eb",x"b37e",x"bbba",x"2ef6",x"3b69",x"39ef",x"14bb",x"3a24",x"3710",x"b416",x"bbad",x"2f8d",x"3b68",x"39eb"),
(x"9f83",x"3ac9",x"36eb",x"35e4",x"bb4d",x"31a2",x"396a",x"3125",x"a035",x"3acc",x"3713",x"3583",x"bb63",x"3153",x"3967",x"3112",x"9c14",x"3ad5",x"370f",x"3a9c",x"b854",x"30fa",x"3965",x"311a"),
(x"9f02",x"3b6a",x"36eb",x"bb89",x"b473",x"31fc",x"3981",x"304c",x"a03c",x"3b86",x"36eb",x"bb99",x"3315",x"330d",x"3982",x"302f",x"9df1",x"3b85",x"3715",x"bbc5",x"2b9a",x"3358",x"397d",x"302d"),
(x"983c",x"3a38",x"3710",x"a856",x"a9ab",x"3bfc",x"3b53",x"3b9f",x"3d81",x"3a3e",x"3711",x"b40c",x"26c2",x"3bbc",x"3b51",x"3b9c",x"1f0f",x"3a43",x"3718",x"ab65",x"b528",x"3b8e",x"3b4b",x"3b9a"),
(x"210e",x"3b6e",x"36eb",x"3be3",x"2ce8",x"30c3",x"397a",x"2f8e",x"21a5",x"3b7a",x"3712",x"3bcf",x"b081",x"3141",x"3978",x"2fbc",x"229f",x"3b7b",x"36eb",x"3bdb",x"1c67",x"320a",x"397c",x"2fa6"),
(x"210e",x"3b6e",x"36eb",x"3be3",x"2ce8",x"30c3",x"397a",x"2f8e",x"20d5",x"3b70",x"3715",x"3bd7",x"b1f9",x"2c2a",x"3977",x"2fab",x"21a5",x"3b7a",x"3712",x"3bcf",x"b081",x"3141",x"3978",x"2fbc"),
(x"2267",x"3af4",x"36eb",x"3958",x"39de",x"2fdf",x"396a",x"2e4c",x"2469",x"3ae4",x"36eb",x"3b75",x"35a2",x"2d46",x"396a",x"2e25",x"243c",x"3ae3",x"3710",x"3b6a",x"35bb",x"2efe",x"3965",x"2e26"),
(x"9889",x"3a27",x"36eb",x"baa4",x"b859",x"2fe5",x"3b6b",x"39ef",x"951c",x"3a29",x"3711",x"ba7f",x"b887",x"3089",x"3b6a",x"39eb",x"14bb",x"3a24",x"3710",x"b416",x"bbad",x"2f8d",x"3b68",x"39eb"),
(x"1e52",x"3a48",x"36eb",x"3be6",x"308e",x"2c41",x"3900",x"2982",x"1d9c",x"3a48",x"3718",x"3be6",x"309f",x"2baa",x"38fa",x"2966",x"1d4f",x"3a5b",x"3715",x"3bfa",x"a70a",x"2c48",x"38f9",x"29b5"),
(x"9889",x"3a27",x"36eb",x"baa4",x"b859",x"2fe5",x"3b6b",x"39ef",x"9b9c",x"3a30",x"36eb",x"bbf4",x"9ef6",x"2ebb",x"3b6d",x"39ef",x"99ac",x"3a30",x"3710",x"bbcc",x"b227",x"2f2e",x"3b6c",x"39eb"),
(x"998f",x"3ad4",x"36eb",x"3b7d",x"b521",x"3095",x"3966",x"312c",x"9c14",x"3ad5",x"370f",x"3a9c",x"b854",x"30fa",x"3965",x"311a",x"9c56",x"3adb",x"370e",x"3b25",x"370d",x"2d68",x"3963",x"311c"),
(x"a30f",x"3a97",x"36eb",x"b6fe",x"bb25",x"2ea6",x"398d",x"2aa4",x"a2cb",x"3a9a",x"3714",x"b972",x"b9bb",x"30de",x"3988",x"2a88",x"9d1e",x"3a94",x"3711",x"b4dc",x"bb97",x"2d61",x"3987",x"2ad2"),
(x"865b",x"3a3e",x"36eb",x"b9db",x"396c",x"2c1a",x"3b71",x"39ef",x"3d81",x"3a3e",x"3711",x"ba7a",x"38b0",x"283c",x"3b70",x"39ea",x"983c",x"3a38",x"3710",x"bb2f",x"36d9",x"2e52",x"3b6e",x"39eb"),
(x"8d14",x"3b00",x"36eb",x"3776",x"3b0b",x"2d41",x"3969",x"2e88",x"2267",x"3af4",x"36eb",x"3958",x"39de",x"2fdf",x"396a",x"2e4c",x"21ba",x"3af2",x"3712",x"384e",x"3ab0",x"2ec7",x"3965",x"2e4d"),
(x"1e6c",x"3a5e",x"36eb",x"39df",x"b964",x"2d28",x"38fe",x"29db",x"1e18",x"3a5b",x"36eb",x"3bfa",x"a0b5",x"2cb4",x"38fe",x"29d0",x"1d4f",x"3a5b",x"3715",x"3bfa",x"a70a",x"2c48",x"38f9",x"29b5"),
(x"9f02",x"3ae5",x"36eb",x"3ad3",x"3822",x"2c4d",x"3962",x"3131",x"9aca",x"3ada",x"36eb",x"3b19",x"3744",x"2cf7",x"3965",x"312d",x"9c56",x"3adb",x"370e",x"3b25",x"370d",x"2d68",x"3963",x"311c"),
(x"1d3a",x"3b33",x"36eb",x"bbfe",x"1ea7",x"2828",x"397e",x"308a",x"1737",x"3b47",x"36eb",x"bb4a",x"b677",x"2cf9",x"397f",x"3074",x"1882",x"3b48",x"370e",x"bb5f",x"b5f1",x"2f4d",x"397b",x"306f"),
(x"8d14",x"3b00",x"36eb",x"3776",x"3b0b",x"2d41",x"3969",x"2e88",x"08f2",x"3afe",x"3716",x"37e9",x"3af1",x"2aa7",x"3963",x"2e82",x"9588",x"3b01",x"3716",x"3bde",x"31b5",x"2825",x"3963",x"2e8b"),
(x"22d4",x"3a69",x"36eb",x"39ed",x"b94b",x"2f45",x"38fd",x"2a25",x"1e6c",x"3a5e",x"36eb",x"39df",x"b964",x"2d28",x"38fe",x"29db",x"1e3f",x"3a60",x"3715",x"395d",x"b9e3",x"2de3",x"38f9",x"29c9"),
(x"9a71",x"3a91",x"3711",x"bb12",x"b763",x"2ca3",x"38f6",x"1f45",x"990c",x"3a8d",x"3712",x"bbf7",x"283f",x"2d8f",x"38f7",x"1fc8",x"9acb",x"3a8c",x"36eb",x"bbf8",x"a379",x"2d44",x"38fb",x"1f47"),
(x"9c70",x"3a93",x"36eb",x"b7d8",x"baf6",x"2a35",x"38fb",x"1e54",x"9d1e",x"3a94",x"3711",x"b4dc",x"bb97",x"2d61",x"38f6",x"1ea7",x"9a71",x"3a91",x"3711",x"bb12",x"b763",x"2ca3",x"38f6",x"1f45"),
(x"9f11",x"3ae7",x"36eb",x"39e9",x"b955",x"2e31",x"3961",x"3132",x"9f02",x"3ae5",x"36eb",x"3ad3",x"3822",x"2c4d",x"3962",x"3131",x"9f72",x"3ae4",x"3713",x"3b5b",x"3634",x"2c03",x"3961",x"311c"),
(x"1d3a",x"3b33",x"36eb",x"bbfe",x"1ea7",x"2828",x"397e",x"308a",x"1d56",x"3b33",x"3716",x"bbff",x"20c2",x"2138",x"3978",x"3084",x"1820",x"3b1f",x"370f",x"bad7",x"3821",x"29e6",x"3978",x"309b"),
(x"9427",x"3b01",x"36eb",x"3b23",x"b71c",x"2cde",x"3963",x"2eda",x"9588",x"3b01",x"3716",x"3bde",x"31b5",x"2825",x"3960",x"2efe",x"8010",x"3b06",x"3714",x"39e8",x"b951",x"2f27",x"3961",x"2f04"),
(x"22d4",x"3a69",x"36eb",x"39ed",x"b94b",x"2f45",x"38fd",x"2a25",x"21e0",x"3a69",x"3719",x"39a6",x"b994",x"2fc6",x"38f8",x"2a02",x"21d8",x"3a6b",x"3719",x"3250",x"3bca",x"2f22",x"38f7",x"2a09"),
(x"9acb",x"3a8c",x"36eb",x"bbf8",x"a379",x"2d44",x"38fb",x"1f47",x"990c",x"3a8d",x"3712",x"bbf7",x"283f",x"2d8f",x"38f7",x"1fc8",x"9ae8",x"3a82",x"3712",x"bb92",x"3509",x"2cb0",x"38f7",x"2098"),
(x"9d1a",x"3aec",x"3710",x"3833",x"bac7",x"2d1d",x"3989",x"274a",x"9476",x"3aef",x"3713",x"30a8",x"bbe9",x"22dc",x"3988",x"2790",x"9096",x"3aef",x"36eb",x"3046",x"bbe8",x"2cb7",x"398d",x"27a9"),
(x"9f11",x"3ae7",x"36eb",x"39e9",x"b955",x"2e31",x"398e",x"2729",x"9f87",x"3ae7",x"3713",x"3b09",x"b791",x"2ab8",x"3989",x"2710",x"9d1a",x"3aec",x"3710",x"3833",x"bac7",x"2d1d",x"3989",x"274a"),
(x"9bdf",x"3b17",x"36eb",x"b73f",x"3b1a",x"2d3c",x"397c",x"30ae",x"173f",x"3b20",x"36eb",x"bab4",x"3859",x"2a66",x"397c",x"309f",x"1820",x"3b1f",x"370f",x"bad7",x"3821",x"29e6",x"3978",x"309b"),
(x"141e",x"3b05",x"36eb",x"397a",x"b9b6",x"309a",x"3964",x"2ee0",x"8010",x"3b06",x"3714",x"39e8",x"b951",x"2f27",x"3961",x"2f04",x"1f40",x"3b15",x"3717",x"3a77",x"b889",x"310e",x"3965",x"2f1f"),
(x"1e72",x"3a6c",x"36eb",x"3b01",x"3745",x"3141",x"38fa",x"2a64",x"2283",x"3a6d",x"36eb",x"32cb",x"3bc1",x"2fc5",x"38fc",x"2a36",x"21d8",x"3a6b",x"3719",x"3250",x"3bca",x"2f22",x"38f7",x"2a09"),
(x"9bea",x"3a84",x"36eb",x"bb57",x"3625",x"2e99",x"38fc",x"2028",x"9ae8",x"3a82",x"3712",x"bb92",x"3509",x"2cb0",x"38f7",x"2098",x"a16d",x"3a60",x"3711",x"bb70",x"3585",x"3014",x"38fa",x"22e8"),
(x"1a19",x"3aef",x"3712",x"b2e8",x"bbcb",x"2c10",x"3988",x"27d6",x"1f35",x"3aed",x"3711",x"b934",x"ba0d",x"2c16",x"3988",x"280f",x"1ecc",x"3aeb",x"36eb",x"b74a",x"bb15",x"2de4",x"398d",x"2814"),
(x"9096",x"3aef",x"36eb",x"3046",x"bbe8",x"2cb7",x"398d",x"27a9",x"9476",x"3aef",x"3713",x"30a8",x"bbe9",x"22dc",x"3988",x"2790",x"1a19",x"3aef",x"3712",x"b2e8",x"bbcb",x"2c10",x"3988",x"27d6"),
(x"9bdf",x"3b17",x"36eb",x"b73f",x"3b1a",x"2d3c",x"397c",x"30ae",x"9a85",x"3b15",x"3713",x"b7c2",x"3af3",x"2e28",x"3977",x"30a9",x"9d28",x"3b16",x"3712",x"3721",x"3b24",x"2bf9",x"3977",x"30ae"),
(x"2078",x"3b14",x"36eb",x"3aff",x"b73c",x"3197",x"3968",x"2efa",x"1f40",x"3b15",x"3717",x"3a77",x"b889",x"310e",x"3965",x"2f1f",x"221f",x"3b30",x"3713",x"3bc6",x"b1be",x"30de",x"396b",x"2f42"),
(x"a25f",x"3a5e",x"36eb",x"bb99",x"345f",x"30d6",x"38ff",x"22bb",x"a16d",x"3a60",x"3711",x"bb70",x"3585",x"3014",x"38fa",x"22e8",x"a2e9",x"3a41",x"3711",x"bbe4",x"2d1d",x"308c",x"38fc",x"2478"),
(x"2284",x"3adf",x"36eb",x"baaf",x"b860",x"2a70",x"398d",x"285d",x"1ecc",x"3aeb",x"36eb",x"b74a",x"bb15",x"2de4",x"398d",x"2814",x"1f35",x"3aed",x"3711",x"b934",x"ba0d",x"2c16",x"3988",x"280f"),
(x"9d97",x"3b18",x"36eb",x"38ae",x"3a73",x"2d49",x"397c",x"30b1",x"9d28",x"3b16",x"3712",x"3721",x"3b24",x"2bf9",x"3977",x"30ae",x"9ff6",x"3b1a",x"3711",x"35dd",x"3b65",x"2eae",x"3977",x"30b5"),
(x"22be",x"3b4b",x"36eb",x"3bea",x"ae0a",x"2f10",x"3973",x"2f49",x"231e",x"3b30",x"36eb",x"3bbf",x"b113",x"322d",x"396e",x"2f22",x"221f",x"3b30",x"3713",x"3bc6",x"b1be",x"30de",x"396b",x"2f42"),
(x"1e72",x"3a6c",x"36eb",x"3b01",x"3745",x"3141",x"3969",x"2cf7",x"20ca",x"3a73",x"3715",x"39d1",x"b974",x"2cc6",x"3964",x"2d15",x"21d1",x"3a75",x"36eb",x"3a0e",x"b929",x"2e76",x"3969",x"2d12"),
(x"1e72",x"3a6c",x"36eb",x"3b01",x"3745",x"3141",x"3969",x"2cf7",x"1e5a",x"3a6d",x"3718",x"3af5",x"b7e1",x"2460",x"3963",x"2d03",x"20ca",x"3a73",x"3715",x"39d1",x"b974",x"2cc6",x"3964",x"2d15"),
(x"a382",x"3a1e",x"36eb",x"bbe8",x"ad68",x"3010",x"3903",x"256b",x"a397",x"3a41",x"36eb",x"bbe6",x"2c77",x"308c",x"3901",x"2450",x"a2e9",x"3a41",x"3711",x"bbe4",x"2d1d",x"308c",x"38fc",x"2478"),
(x"234c",x"3acf",x"36eb",x"bbfa",x"ac62",x"2617",x"398d",x"28a0",x"2284",x"3adf",x"36eb",x"baaf",x"b860",x"2a70",x"398d",x"285d",x"22bc",x"3adf",x"3717",x"bb6f",x"b5e4",x"261e",x"3987",x"285d"),
(x"9f8c",x"3b1c",x"36eb",x"2e28",x"3be6",x"3005",x"397c",x"30b7",x"9ff6",x"3b1a",x"3711",x"35dd",x"3b65",x"2eae",x"3977",x"30b5",x"a20d",x"3b19",x"3712",x"b5a6",x"3b63",x"30cc",x"3977",x"30bd"),
(x"22be",x"3b4b",x"36eb",x"3bea",x"ae0a",x"2f10",x"3973",x"2f49",x"2273",x"3b4b",x"3717",x"3bf0",x"af0f",x"2aec",x"396f",x"2f6c",x"2386",x"3b62",x"370f",x"3bdd",x"b0de",x"2e6c",x"3974",x"2f86"),
(x"21d1",x"3a75",x"36eb",x"3a0e",x"b929",x"2e76",x"3969",x"2d12",x"20ca",x"3a73",x"3715",x"39d1",x"b974",x"2cc6",x"3964",x"2d15",x"2288",x"3a7e",x"3718",x"3b13",x"b732",x"2fec",x"3964",x"2d2f"),
(x"a382",x"3a1e",x"36eb",x"bbe8",x"ad68",x"3010",x"3903",x"256b",x"a2ee",x"3a1f",x"3714",x"bbec",x"ad02",x"2f4a",x"38fe",x"258f",x"a1ea",x"3a0f",x"3712",x"bb45",x"b640",x"30a6",x"38ff",x"2610"),
(x"9b9c",x"3a30",x"36eb",x"bbf4",x"9ef6",x"2ebb",x"3b6d",x"39ef",x"9a2a",x"3a3a",x"36eb",x"bb02",x"3776",x"2fc8",x"3b6f",x"39ef",x"983c",x"3a38",x"3710",x"bb2f",x"36d9",x"2e52",x"3b6e",x"39eb"),
(x"22be",x"3aba",x"36eb",x"bbcf",x"32aa",x"2bc5",x"398d",x"28f8",x"234c",x"3acf",x"36eb",x"bbfa",x"ac62",x"2617",x"398d",x"28a0",x"2365",x"3ace",x"3715",x"bbfe",x"2412",x"2867",x"3988",x"28a3"),
(x"a2ba",x"3b1c",x"36eb",x"b913",x"3a0d",x"310f",x"397b",x"30c4",x"a20d",x"3b19",x"3712",x"b5a6",x"3b63",x"30cc",x"3977",x"30bd",x"a34c",x"3b12",x"3711",x"bbb2",x"332f",x"30f4",x"3976",x"30c7"),
(x"2414",x"3b61",x"36eb",x"3be4",x"aadf",x"30ee",x"3977",x"2f68",x"2386",x"3b62",x"370f",x"3bdd",x"b0de",x"2e6c",x"3974",x"2f86",x"2312",x"3b69",x"370d",x"3b0d",x"370c",x"3169",x"3976",x"2f8f"),
(x"2349",x"3a7d",x"36eb",x"3bbf",x"b333",x"2ed2",x"396a",x"2d27",x"2288",x"3a7e",x"3718",x"3b13",x"b732",x"2fec",x"3964",x"2d2f",x"22dc",x"3a86",x"3712",x"3bf0",x"2c20",x"2e95",x"3965",x"2d3f"),
(x"a269",x"3a0c",x"36eb",x"bab2",x"b834",x"30cb",x"3904",x"2600",x"a1ea",x"3a0f",x"3712",x"bb45",x"b640",x"30a6",x"38ff",x"2610",x"9d7f",x"3a00",x"3715",x"b93c",x"b9e9",x"3110",x"38ff",x"26b7"),
(x"207d",x"3aaa",x"36eb",x"bac2",x"3833",x"2e8a",x"398d",x"2945",x"22be",x"3aba",x"36eb",x"bbcf",x"32aa",x"2bc5",x"398d",x"28f8",x"2308",x"3ab8",x"3714",x"bb81",x"3558",x"2da6",x"3988",x"2900"),
(x"a3f7",x"3b12",x"36eb",x"bbe5",x"adbc",x"3036",x"397a",x"30ce",x"a34c",x"3b12",x"3711",x"bbb2",x"332f",x"30f4",x"3976",x"30c7",x"a273",x"3b06",x"3712",x"bae4",x"b7c3",x"30c9",x"3975",x"30d1"),
(x"226e",x"3b6e",x"36eb",x"3571",x"3b6d",x"30cc",x"397a",x"2f84",x"23bf",x"3b6c",x"36eb",x"3af6",x"3714",x"32f0",x"3979",x"2f79",x"2312",x"3b69",x"370d",x"3b0d",x"370c",x"3169",x"3976",x"2f8f"),
(x"2324",x"3a89",x"36eb",x"3bbf",x"3370",x"2dad",x"396a",x"2d3f",x"22dc",x"3a86",x"3712",x"3bf0",x"2c20",x"2e95",x"3965",x"2d3f",x"2257",x"3a89",x"3712",x"3298",x"3bcc",x"2d84",x"3965",x"2d48"),
(x"9dfd",x"39fc",x"36eb",x"b7cb",x"bae6",x"3068",x"3904",x"26ad",x"9d7f",x"3a00",x"3715",x"b93c",x"b9e9",x"3110",x"38ff",x"26b7",x"17a2",x"39fb",x"3715",x"9ef6",x"bbee",x"302a",x"38ff",x"273a"),
(x"1ce6",x"3aa0",x"36eb",x"b9cd",x"3979",x"2caa",x"398d",x"297b",x"207d",x"3aaa",x"36eb",x"bac2",x"3833",x"2e8a",x"398d",x"2945",x"20ef",x"3aa9",x"3715",x"ba65",x"38c1",x"2d9c",x"3988",x"2949"),
(x"a2c3",x"3b03",x"36eb",x"b902",x"ba23",x"306a",x"3979",x"30dd",x"a273",x"3b06",x"3712",x"bae4",x"b7c3",x"30c9",x"3975",x"30d1",x"a040",x"3b03",x"3713",x"b607",x"bb5e",x"2e4f",x"3973",x"30d9"),
(x"210e",x"3b6e",x"36eb",x"3be3",x"2ce8",x"30c3",x"397a",x"2f8e",x"226e",x"3b6e",x"36eb",x"3571",x"3b6d",x"30cc",x"397a",x"2f84",x"2243",x"3b6c",x"3713",x"3451",x"3bac",x"2d81",x"3976",x"2f9b"),
(x"2058",x"3a8a",x"36eb",x"2c58",x"3bf7",x"2bc5",x"396a",x"2d59",x"22c6",x"3a8b",x"36eb",x"2eda",x"3bea",x"2e47",x"396a",x"2d45",x"2257",x"3a89",x"3712",x"3298",x"3bcc",x"2d84",x"3965",x"2d48"),
(x"20e4",x"39fc",x"36eb",x"366a",x"bb44",x"2f81",x"3905",x"27be",x"17aa",x"39f8",x"36eb",x"96f6",x"bbf5",x"2e99",x"3905",x"2736",x"17a2",x"39fb",x"3715",x"9ef6",x"bbee",x"302a",x"38ff",x"273a"),
(x"1a1b",x"3a9d",x"36eb",x"35a5",x"3b74",x"2d53",x"398d",x"298f",x"1ce6",x"3aa0",x"36eb",x"b9cd",x"3979",x"2caa",x"398d",x"297b",x"1d4c",x"3a9f",x"3717",x"b939",x"3a0b",x"29e0",x"3988",x"2980"),
(x"9efd",x"3aff",x"36eb",x"b94d",x"39f2",x"2dc5",x"3977",x"30e9",x"9ff8",x"3b01",x"36eb",x"b3f1",x"bbbc",x"2b5c",x"3977",x"30e7",x"a040",x"3b03",x"3713",x"b607",x"bb5e",x"2e4f",x"3973",x"30d9"),
(x"20d5",x"3b70",x"3715",x"a587",x"307a",x"3beb",x"3b45",x"3b1b",x"9cbb",x"3b6c",x"3715",x"19bc",x"a6cf",x"3bff",x"3b51",x"3b1b",x"21a5",x"3b7a",x"3712",x"29f0",x"2b1d",x"3bfa",x"3b43",x"3b16"),
(x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c",x"1882",x"3b48",x"370e",x"b004",x"a71d",x"3bef",x"3b4d",x"3b2b",x"9cbb",x"3b6c",x"3715",x"19bc",x"a6cf",x"3bff",x"3b51",x"3b1b"),
(x"20f8",x"3b6d",x"3716",x"a0ea",x"a786",x"3bfe",x"3b45",x"3b1c",x"9cbb",x"3b6c",x"3715",x"19bc",x"a6cf",x"3bff",x"3b51",x"3b1b",x"20d5",x"3b70",x"3715",x"a587",x"307a",x"3beb",x"3b45",x"3b1b"),
(x"2273",x"3b4b",x"3717",x"abf6",x"25ae",x"3bfb",x"3b44",x"3b2a",x"1d56",x"3b33",x"3716",x"aadf",x"a6b5",x"3bfc",x"3b4b",x"3b34",x"1882",x"3b48",x"370e",x"b004",x"a71d",x"3bef",x"3b4d",x"3b2b"),
(x"2058",x"3a8a",x"36eb",x"2c58",x"3bf7",x"2bc5",x"396a",x"2d59",x"2091",x"3a89",x"3717",x"2a0a",x"3bfc",x"284d",x"3964",x"2d56",x"1f4b",x"3a8a",x"3716",x"38f4",x"3a42",x"2c09",x"3964",x"2d5e"),
(x"24bd",x"3a0a",x"36eb",x"39f2",x"b938",x"30b5",x"3904",x"283d",x"20e4",x"39fc",x"36eb",x"366a",x"bb44",x"2f81",x"3905",x"27be",x"210b",x"3a00",x"3713",x"382e",x"baba",x"306c",x"3900",x"27ca"),
(x"0e53",x"3aa0",x"3714",x"39a7",x"399e",x"2d1e",x"3988",x"29b0",x"987a",x"3aa6",x"3714",x"397e",x"39c5",x"2dbf",x"3988",x"29d2",x"98cf",x"3aa9",x"36eb",x"3976",x"39cc",x"2dcc",x"398e",x"29d2"),
(x"1a1b",x"3a9d",x"36eb",x"35a5",x"3b74",x"2d53",x"398d",x"298f",x"19fe",x"3a9c",x"3717",x"2c95",x"3bf9",x"2918",x"3988",x"2997",x"0e53",x"3aa0",x"3714",x"39a7",x"399e",x"2d1e",x"3988",x"29b0"),
(x"9efd",x"3aff",x"36eb",x"b94d",x"39f2",x"2dc5",x"3977",x"30e9",x"9e8d",x"3aff",x"3716",x"bac7",x"383c",x"283f",x"3972",x"30dd",x"a17b",x"3afb",x"3711",x"b8c8",x"3a4e",x"30a8",x"3971",x"30e7"),
(x"2585",x"3a1d",x"36eb",x"3bc4",x"b27a",x"3012",x"3904",x"2891",x"24bd",x"3a0a",x"36eb",x"39f2",x"b938",x"30b5",x"3904",x"283d",x"2466",x"3a0c",x"3715",x"3ae0",x"b7cf",x"30d4",x"38ff",x"2836"),
(x"98cf",x"3aa9",x"36eb",x"3976",x"39cc",x"2dcc",x"398e",x"29d2",x"987a",x"3aa6",x"3714",x"397e",x"39c5",x"2dbf",x"3988",x"29d2",x"9e62",x"3aad",x"3716",x"37d5",x"3af0",x"2d8e",x"3989",x"29ff"),
(x"a282",x"3afc",x"36eb",x"b9ec",x"392b",x"31e4",x"3975",x"30f4",x"a17b",x"3afb",x"3711",x"b8c8",x"3a4e",x"30a8",x"3971",x"30e7",x"a407",x"3aeb",x"370f",x"bb4b",x"35cc",x"3223",x"396f",x"30f8"),
(x"229f",x"3b7b",x"36eb",x"3bdb",x"1c67",x"320a",x"397c",x"2fa6",x"21a5",x"3b7a",x"3712",x"3bcf",x"b081",x"3141",x"3978",x"2fbc",x"20f7",x"3b90",x"370e",x"3b7b",x"34a9",x"3270",x"397b",x"2fe0"),
(x"1e77",x"3a8d",x"3715",x"3ac1",x"b812",x"3146",x"3964",x"2d67",x"1f29",x"3a92",x"3714",x"b879",x"347b",x"3a3d",x"3964",x"2d71",x"2147",x"3a9a",x"3718",x"3ac6",x"b7dc",x"3286",x"3964",x"2d86"),
(x"255d",x"3a30",x"36eb",x"3b6e",x"3575",x"309f",x"3903",x"28e0",x"2585",x"3a1d",x"36eb",x"3bc4",x"b27a",x"3012",x"3904",x"2891",x"253f",x"3a1e",x"3715",x"3bec",x"abe2",x"2fce",x"38ff",x"2887"),
(x"9c3a",x"3a58",x"3714",x"b05e",x"2194",x"3bec",x"3b54",x"3b91",x"a2e9",x"3a41",x"3711",x"acd1",x"2504",x"3bf9",x"3b5c",x"3b9b",x"a16d",x"3a60",x"3711",x"b115",x"27d5",x"3be4",x"3b59",x"3b8d"),
(x"9c3a",x"3a58",x"3714",x"b05e",x"2194",x"3bec",x"3b54",x"3b91",x"a0d2",x"3a3e",x"3713",x"b0f4",x"19bc",x"3be7",x"3b59",x"3b9c",x"a2e9",x"3a41",x"3711",x"acd1",x"2504",x"3bf9",x"3b5c",x"3b9b"),
(x"9e13",x"3aae",x"36eb",x"353f",x"3b87",x"2d28",x"398e",x"29f7",x"9e62",x"3aad",x"3716",x"37d5",x"3af0",x"2d8e",x"3989",x"29ff",x"a13d",x"3aae",x"3716",x"a345",x"3bf7",x"2dcc",x"3989",x"2a21"),
(x"a471",x"3aeb",x"36eb",x"bbbc",x"3212",x"3175",x"3972",x"3105",x"a407",x"3aeb",x"370f",x"bb4b",x"35cc",x"3223",x"396f",x"30f8",x"a425",x"3ad8",x"370f",x"bbd3",x"af46",x"3182",x"396c",x"3106"),
(x"22bc",x"3a9c",x"36eb",x"3adb",x"b7e7",x"30ac",x"396a",x"2d88",x"2147",x"3a9a",x"3718",x"3ac6",x"b7dc",x"3286",x"3964",x"2d86",x"2442",x"3ab2",x"3714",x"3b6b",x"b587",x"3095",x"3965",x"2dbe"),
(x"255d",x"3a30",x"36eb",x"3b6e",x"3575",x"309f",x"3903",x"28e0",x"24fc",x"3a2f",x"3717",x"3b55",x"35fd",x"307e",x"38fd",x"28cc",x"2375",x"3a3d",x"3711",x"38a4",x"3a69",x"309a",x"38fd",x"2913"),
(x"a172",x"3ab0",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"398e",x"2a20",x"a13d",x"3aae",x"3716",x"a345",x"3bf7",x"2dcc",x"3989",x"2a21",x"a2d9",x"3aab",x"3714",x"b976",x"39c0",x"3023",x"3989",x"2a41"),
(x"a482",x"3ad7",x"36eb",x"bb61",x"b5a0",x"3119",x"396f",x"3114",x"a425",x"3ad8",x"370f",x"bbd3",x"af46",x"3182",x"396c",x"3106",x"a289",x"3acf",x"370f",x"b891",x"ba73",x"30f5",x"396a",x"310e"),
(x"21ae",x"3b92",x"36eb",x"3ade",x"37ab",x"31d3",x"397f",x"2fd1",x"20f7",x"3b90",x"370e",x"3b7b",x"34a9",x"3270",x"397b",x"2fe0",x"1aac",x"3ba1",x"3712",x"38b5",x"3a3e",x"32bd",x"397d",x"3005"),
(x"2496",x"3ab2",x"36eb",x"3bba",x"b376",x"2f14",x"396a",x"2dbb",x"2442",x"3ab2",x"3714",x"3b6b",x"b587",x"3095",x"3965",x"2dbe",x"24cc",x"3acb",x"3712",x"3bf0",x"aa00",x"2f46",x"3965",x"2df3"),
(x"1fad",x"3a43",x"36eb",x"360d",x"3b5a",x"2ef3",x"3900",x"296f",x"2409",x"3a40",x"36eb",x"3884",x"3a69",x"3249",x"3902",x"292c",x"2375",x"3a3d",x"3711",x"38a4",x"3a69",x"309a",x"38fd",x"2913"),
(x"a38b",x"3aac",x"36eb",x"bacb",x"3812",x"3064",x"398e",x"2a48",x"a2d9",x"3aab",x"3714",x"b976",x"39c0",x"3023",x"3989",x"2a41",x"a38f",x"3aa2",x"3712",x"bbe0",x"2e5e",x"30a3",x"3989",x"2a66"),
(x"9f83",x"3ac9",x"36eb",x"35e4",x"bb4d",x"31a2",x"396a",x"3125",x"a2ad",x"3acb",x"36eb",x"b86e",x"ba87",x"313e",x"396c",x"311e",x"a289",x"3acf",x"370f",x"b891",x"ba73",x"30f5",x"396a",x"310e"),
(x"980d",x"3ba6",x"36eb",x"b996",x"395f",x"33ec",x"3983",x"300b",x"1a0c",x"3ba6",x"36eb",x"38a6",x"3a54",x"3207",x"3982",x"3001",x"1aac",x"3ba1",x"3712",x"38b5",x"3a3e",x"32bd",x"397d",x"3005"),
(x"250f",x"3acc",x"36eb",x"3bef",x"2d09",x"2e69",x"396a",x"2df2",x"24cc",x"3acb",x"3712",x"3bf0",x"aa00",x"2f46",x"3965",x"2df3",x"243c",x"3ae3",x"3710",x"3b6a",x"35bb",x"2efe",x"3965",x"2e26"),
(x"1e52",x"3a48",x"36eb",x"3be6",x"308e",x"2c41",x"3900",x"2982",x"1fad",x"3a43",x"36eb",x"360d",x"3b5a",x"2ef3",x"3900",x"296f",x"1f0f",x"3a43",x"3718",x"38ae",x"3a78",x"2b7c",x"38fb",x"294e"),
(x"a422",x"3aa1",x"36eb",x"bbcf",x"b174",x"303e",x"398e",x"2a77",x"a38f",x"3aa2",x"3712",x"bbe0",x"2e5e",x"30a3",x"3989",x"2a66",x"a2cb",x"3a9a",x"3714",x"b972",x"b9bb",x"30de",x"3988",x"2a88"),
(x"a2e9",x"3a41",x"3711",x"acd1",x"2504",x"3bf9",x"3b5c",x"3b9b",x"a0d2",x"3a3e",x"3713",x"b0f4",x"19bc",x"3be7",x"3b59",x"3b9c",x"a175",x"3a2c",x"3710",x"2828",x"260a",x"3bfe",x"3b5a",x"3ba3"),
(x"a175",x"3a2c",x"3710",x"2828",x"260a",x"3bfe",x"3b5a",x"3ba3",x"a2ee",x"3a1f",x"3714",x"2eb0",x"28fa",x"3bf3",x"3b5c",x"3ba9",x"a2e9",x"3a41",x"3711",x"acd1",x"2504",x"3bf9",x"3b5c",x"3b9b"),
(x"a1ea",x"3a0f",x"3712",x"a587",x"209b",x"3bff",x"3b5b",x"3baf",x"a140",x"3a1c",x"3714",x"2946",x"1ffc",x"3bfe",x"3b5a",x"3baa",x"a099",x"3a14",x"3712",x"2953",x"27b4",x"3bfd",x"3b59",x"3bae"),
(x"a1ea",x"3a0f",x"3712",x"a587",x"209b",x"3bff",x"3b5b",x"3baf",x"a2ee",x"3a1f",x"3714",x"2eb0",x"28fa",x"3bf3",x"3b5c",x"3ba9",x"a140",x"3a1c",x"3714",x"2946",x"1ffc",x"3bfe",x"3b5a",x"3baa"),
(x"9d7f",x"3a00",x"3715",x"a0ea",x"2afd",x"3bfc",x"3b57",x"3bb6",x"a1ea",x"3a0f",x"3712",x"a587",x"209b",x"3bff",x"3b5b",x"3baf",x"9ecc",x"3a0d",x"3714",x"a8bf",x"2c22",x"3bfa",x"3b57",x"3bb0"),
(x"17a2",x"39fb",x"3715",x"27e2",x"29b2",x"3bfc",x"3b51",x"3bb9",x"9d7f",x"3a00",x"3715",x"a0ea",x"2afd",x"3bfc",x"3b57",x"3bb6",x"9aa8",x"3a08",x"3714",x"231d",x"2b5f",x"3bfc",x"3b55",x"3bb3"),
(x"210b",x"3a00",x"3713",x"2b1d",x"aee4",x"3bf0",x"3b4a",x"3bb7",x"17a2",x"39fb",x"3715",x"27e2",x"29b2",x"3bfc",x"3b51",x"3bb9",x"1a1e",x"3a04",x"3715",x"270a",x"a779",x"3bfe",x"3b50",x"3bb5"),
(x"2466",x"3a0c",x"3715",x"a266",x"9d87",x"3bff",x"3b44",x"3bb2",x"210b",x"3a00",x"3713",x"2b1d",x"aee4",x"3bf0",x"3b4a",x"3bb7",x"20b2",x"3a07",x"3716",x"24bc",x"aceb",x"3bf9",x"3b4b",x"3bb4"),
(x"253f",x"3a1e",x"3715",x"a891",x"a7ce",x"3bfd",x"3b41",x"3bab",x"2466",x"3a0c",x"3715",x"a266",x"9d87",x"3bff",x"3b44",x"3bb2",x"2335",x"3a14",x"3714",x"a8e0",x"299e",x"3bfc",x"3b47",x"3baf"),
(x"22d3",x"3a28",x"3715",x"ac67",x"28a5",x"3bf9",x"3b47",x"3ba6",x"24fc",x"3a2f",x"3717",x"ad06",x"2793",x"3bf8",x"3b42",x"3ba3",x"253f",x"3a1e",x"3715",x"a891",x"a7ce",x"3bfd",x"3b41",x"3bab"),
(x"2375",x"3a3d",x"3711",x"a8d9",x"a52b",x"3bfe",x"3b45",x"3b9e",x"24fc",x"3a2f",x"3717",x"ad06",x"2793",x"3bf8",x"3b42",x"3ba3",x"22d3",x"3a28",x"3715",x"ac67",x"28a5",x"3bf9",x"3b47",x"3ba6"),
(x"951c",x"3a29",x"3711",x"abef",x"a8a8",x"3bfa",x"3b52",x"3ba5",x"20d5",x"3a29",x"3714",x"aa45",x"2b10",x"3bfa",x"3b4a",x"3ba6",x"1e4f",x"3a25",x"3711",x"aa66",x"b31a",x"3bca",x"3b4d",x"3ba7"),
(x"1f0f",x"3a43",x"3718",x"ab65",x"b528",x"3b8e",x"3b4b",x"3b9a",x"3d81",x"3a3e",x"3711",x"b40c",x"26c2",x"3bbc",x"3b51",x"3b9c",x"15a0",x"3a42",x"3713",x"b41f",x"ac3a",x"3bb6",x"3b50",x"3b9b"),
(x"16c6",x"3a4b",x"3714",x"ade0",x"a4c2",x"3bf6",x"3b50",x"3b97",x"1d9c",x"3a48",x"3718",x"b420",x"1418",x"3bba",x"3b4c",x"3b98",x"15a0",x"3a42",x"3713",x"b41f",x"ac3a",x"3bb6",x"3b50",x"3b9b"),
(x"16c6",x"3a4b",x"3714",x"ade0",x"a4c2",x"3bf6",x"3b50",x"3b97",x"1d4f",x"3a5b",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3b4d",x"3b90",x"1d9c",x"3a48",x"3718",x"b420",x"1418",x"3bba",x"3b4c",x"3b98"),
(x"20d5",x"3a29",x"3714",x"aa45",x"2b10",x"3bfa",x"3b4a",x"3ba6",x"983c",x"3a38",x"3710",x"a856",x"a9ab",x"3bfc",x"3b53",x"3b9f",x"2375",x"3a3d",x"3711",x"a8d9",x"a52b",x"3bfe",x"3b45",x"3b9e"),
(x"951c",x"3a29",x"3711",x"abef",x"a8a8",x"3bfa",x"3b52",x"3ba5",x"99ac",x"3a30",x"3710",x"aa8d",x"2973",x"3bfb",x"3b53",x"3ba2",x"983c",x"3a38",x"3710",x"a856",x"a9ab",x"3bfc",x"3b53",x"3b9f"),
(x"a1bd",x"39b8",x"3715",x"a1ae",x"23fc",x"3bff",x"3963",x"32c0",x"993e",x"39b7",x"3716",x"a82f",x"2808",x"3bfd",x"3967",x"32be",x"a069",x"397e",x"3718",x"a24c",x"a379",x"3bff",x"3964",x"327c"),
(x"16c6",x"3a4b",x"3714",x"bbf3",x"ae23",x"2b27",x"3b73",x"39ea",x"15a0",x"3a42",x"3713",x"bbc2",x"33a5",x"298a",x"3b71",x"39ea",x"13e1",x"3a42",x"36eb",x"bbf6",x"2a70",x"2d61",x"3b72",x"39ef"),
(x"8dee",x"3a63",x"36eb",x"b46a",x"bb91",x"316a",x"3b7b",x"39ee",x"8dee",x"3a63",x"3718",x"b9e5",x"b968",x"0000",x"3b7a",x"39e9",x"16c6",x"3a4b",x"3714",x"bbf3",x"ae23",x"2b27",x"3b73",x"39ea"),
(x"1c89",x"3761",x"3716",x"b0f9",x"28b2",x"3be5",x"3914",x"3896",x"0f4a",x"3761",x"3712",x"b42b",x"ae69",x"3bae",x"3910",x"3896",x"9e24",x"3783",x"370e",x"afd2",x"a717",x"3bef",x"390a",x"38a1"),
(x"2222",x"3797",x"36eb",x"3b99",x"b315",x"330d",x"395c",x"300e",x"1dd1",x"3756",x"36eb",x"3996",x"b95f",x"33ec",x"395d",x"2fd5",x"1c89",x"3761",x"3716",x"3add",x"b75a",x"334d",x"3958",x"2fd9"),
(x"1ba5",x"384b",x"3714",x"2c39",x"a9a5",x"3bf9",x"391a",x"38ee",x"2226",x"384e",x"3713",x"291b",x"ab55",x"3bfb",x"3923",x"38ef",x"2079",x"383b",x"3712",x"2a69",x"a87e",x"3bfc",x"3920",x"38e4"),
(x"2498",x"383f",x"3711",x"2481",x"a54c",x"3bff",x"392a",x"38e7",x"23f2",x"3838",x"3712",x"aa38",x"2d35",x"3bf6",x"3927",x"38e2",x"21e0",x"3837",x"3711",x"2994",x"a977",x"3bfc",x"3922",x"38e2"),
(x"2079",x"383b",x"3712",x"2a69",x"a87e",x"3bfc",x"3920",x"38e4",x"2226",x"384e",x"3713",x"291b",x"ab55",x"3bfb",x"3923",x"38ef",x"242c",x"384b",x"3712",x"2a73",x"aa97",x"3bfa",x"3928",x"38ed"),
(x"2000",x"3854",x"3718",x"2e36",x"2153",x"3bf6",x"391f",x"38f3",x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8",x"2360",x"3856",x"3711",x"2fec",x"2c2c",x"3beb",x"3926",x"38f4"),
(x"221a",x"3885",x"3713",x"2e9c",x"b367",x"3bbd",x"3926",x"390f",x"2437",x"3883",x"370f",x"1df0",x"2631",x"3bff",x"392a",x"390d",x"2010",x"3876",x"370e",x"a6dc",x"a5c2",x"3bfe",x"3921",x"3907"),
(x"219e",x"386d",x"3713",x"2538",x"2c79",x"3bfa",x"3924",x"3901",x"2010",x"3876",x"370e",x"a6dc",x"a5c2",x"3bfe",x"3921",x"3907",x"2437",x"3883",x"370f",x"1df0",x"2631",x"3bff",x"392a",x"390d"),
(x"24fa",x"3866",x"370f",x"2ec5",x"9a24",x"3bf4",x"392d",x"38fd",x"21a8",x"386a",x"3713",x"27ef",x"a84d",x"3bfd",x"3923",x"38ff",x"219e",x"386d",x"3713",x"2538",x"2c79",x"3bfa",x"3924",x"3901"),
(x"21a8",x"386a",x"3713",x"27ef",x"a84d",x"3bfd",x"3923",x"38ff",x"24fa",x"3866",x"370f",x"2ec5",x"9a24",x"3bf4",x"392d",x"38fd",x"2360",x"3856",x"3711",x"2fec",x"2c2c",x"3beb",x"3926",x"38f4"),
(x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8",x"1ce8",x"3862",x"3713",x"a5bc",x"37de",x"3af6",x"391c",x"38fb",x"2072",x"3865",x"3710",x"2c5b",x"30a5",x"3be5",x"3921",x"38fd"),
(x"2072",x"3865",x"3710",x"2c5b",x"30a5",x"3be5",x"3921",x"38fd",x"21a8",x"386a",x"3713",x"27ef",x"a84d",x"3bfd",x"3923",x"38ff",x"2360",x"3856",x"3711",x"2fec",x"2c2c",x"3beb",x"3926",x"38f4"),
(x"9959",x"38c4",x"3715",x"26c2",x"2c65",x"3bfa",x"3914",x"3933",x"1e50",x"38c4",x"3712",x"2f67",x"2981",x"3bf0",x"391e",x"3933",x"125b",x"38b5",x"3717",x"2ff2",x"2a7a",x"3bed",x"3918",x"392b"),
(x"24ba",x"38af",x"3712",x"3163",x"2345",x"3be2",x"392b",x"3927",x"245f",x"38a6",x"3714",x"2860",x"2f8b",x"3bf0",x"3929",x"3922",x"2323",x"38a3",x"3716",x"2cd8",x"27e2",x"3bf9",x"3926",x"3920"),
(x"2116",x"38a4",x"3716",x"a818",x"2d02",x"3bf8",x"3922",x"3921",x"2074",x"38bd",x"3711",x"a412",x"2d5c",x"3bf8",x"3920",x"392f",x"2458",x"38b7",x"3714",x"9553",x"2b62",x"3bfc",x"3929",x"392b"),
(x"2074",x"38bd",x"3711",x"a412",x"2d5c",x"3bf8",x"3920",x"392f",x"1e07",x"38ab",x"3714",x"24fd",x"2da9",x"3bf7",x"391d",x"3925",x"1acb",x"38b1",x"3714",x"3036",x"273e",x"3bed",x"391b",x"3928"),
(x"125b",x"38b5",x"3717",x"2ff2",x"2a7a",x"3bed",x"3918",x"392b",x"1e50",x"38c4",x"3712",x"2f67",x"2981",x"3bf0",x"391e",x"3933",x"1f03",x"38c0",x"3711",x"327d",x"975f",x"3bd5",x"391f",x"3931"),
(x"1f03",x"38c0",x"3711",x"327d",x"975f",x"3bd5",x"391f",x"3931",x"2074",x"38bd",x"3711",x"a412",x"2d5c",x"3bf8",x"3920",x"392f",x"1acb",x"38b1",x"3714",x"3036",x"273e",x"3bed",x"391b",x"3928"),
(x"1f3f",x"38cf",x"3712",x"3146",x"ac91",x"3bde",x"391f",x"3939",x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b"),
(x"9aa8",x"38e6",x"3718",x"a138",x"2e94",x"3bf4",x"3914",x"3947",x"9fe7",x"38e6",x"3719",x"23bb",x"a7db",x"3bfe",x"390f",x"3947",x"9ff6",x"38e8",x"3719",x"290e",x"2efe",x"3bf2",x"390f",x"3948"),
(x"9920",x"38e4",x"3718",x"ab4f",x"a52b",x"3bfc",x"3915",x"3946",x"9aa8",x"38e6",x"3718",x"a138",x"2e94",x"3bf4",x"3914",x"3947",x"1c29",x"38ee",x"3718",x"2e3a",x"9fc8",x"3bf6",x"391c",x"394b"),
(x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"9dca",x"38de",x"3715",x"ad65",x"2c5a",x"3bf3",x"3911",x"3942",x"9920",x"38e4",x"3718",x"ab4f",x"a52b",x"3bfc",x"3915",x"3946"),
(x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"9d58",x"38c8",x"3717",x"ad2f",x"aecb",x"3bed",x"3912",x"3935",x"a0a3",x"38d3",x"3718",x"acf2",x"991e",x"3bf9",x"390d",x"393c"),
(x"a0f6",x"38cb",x"3712",x"b59c",x"b36a",x"3b42",x"390d",x"3937",x"a0a3",x"38d3",x"3718",x"acf2",x"991e",x"3bf9",x"390d",x"393c",x"9d58",x"38c8",x"3717",x"ad2f",x"aecb",x"3bed",x"3912",x"3935"),
(x"3b57",x"38d5",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3917",x"393d",x"1f3f",x"38cf",x"3712",x"3146",x"ac91",x"3bde",x"391f",x"3939",x"9b02",x"38c7",x"3716",x"3009",x"ada6",x"3be7",x"3914",x"3935"),
(x"9b02",x"38c7",x"3716",x"3009",x"ada6",x"3be7",x"3914",x"3935",x"1f3f",x"38cf",x"3712",x"3146",x"ac91",x"3bde",x"391f",x"3939",x"1e50",x"38c4",x"3712",x"2f67",x"2981",x"3bf0",x"391e",x"3933"),
(x"9607",x"38b2",x"3717",x"17c8",x"1f79",x"3c00",x"3915",x"3929",x"9ec5",x"38b7",x"3718",x"2c00",x"a90e",x"3bfa",x"3910",x"392c",x"9abe",x"38bf",x"3714",x"2581",x"2e8a",x"3bf4",x"3913",x"3930"),
(x"9607",x"38b2",x"3717",x"17c8",x"1f79",x"3c00",x"3915",x"3929",x"9e13",x"38a8",x"3715",x"251e",x"ad06",x"3bf9",x"3911",x"3924",x"9ec5",x"38b7",x"3718",x"2c00",x"a90e",x"3bfa",x"3910",x"392c"),
(x"9e13",x"38a8",x"3715",x"251e",x"ad06",x"3bf9",x"3911",x"3924",x"a123",x"3899",x"3714",x"adba",x"a266",x"3bf7",x"390c",x"391b",x"a29f",x"389f",x"3714",x"975f",x"ac2c",x"3bfb",x"3909",x"391e"),
(x"a123",x"3899",x"3714",x"adba",x"a266",x"3bf7",x"390c",x"391b",x"a180",x"3883",x"3715",x"b468",x"a47a",x"3bb0",x"390c",x"390f",x"a3b3",x"3886",x"3712",x"b106",x"a738",x"3be5",x"3907",x"3910"),
(x"a180",x"3883",x"3715",x"b468",x"a47a",x"3bb0",x"390c",x"390f",x"a0d7",x"3872",x"3717",x"b273",x"af43",x"3bc8",x"390d",x"3905",x"a294",x"386e",x"3710",x"b550",x"ae33",x"3b81",x"3909",x"3903"),
(x"a0d7",x"3872",x"3717",x"b273",x"af43",x"3bc8",x"390d",x"3905",x"9ad5",x"3864",x"3711",x"2e23",x"aa31",x"3bf4",x"3914",x"38fd",x"9faa",x"385f",x"3712",x"ab5f",x"a345",x"3bfc",x"390f",x"38fa"),
(x"11f0",x"3862",x"3712",x"add2",x"304b",x"3be4",x"3918",x"38fc",x"1b46",x"3853",x"3716",x"af4d",x"2a5f",x"3bf0",x"391a",x"38f3",x"9faa",x"385f",x"3712",x"ab5f",x"a345",x"3bfc",x"390f",x"38fa"),
(x"11f0",x"3862",x"3712",x"add2",x"304b",x"3be4",x"3918",x"38fc",x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8",x"1b46",x"3853",x"3716",x"af4d",x"2a5f",x"3bf0",x"391a",x"38f3"),
(x"11f0",x"3862",x"3712",x"add2",x"304b",x"3be4",x"3918",x"38fc",x"1ce8",x"3862",x"3713",x"a5bc",x"37de",x"3af6",x"391c",x"38fb",x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8"),
(x"1b46",x"3853",x"3716",x"af4d",x"2a5f",x"3bf0",x"391a",x"38f3",x"1c86",x"385d",x"3718",x"2c13",x"31c5",x"3bda",x"391c",x"38f8",x"2000",x"3854",x"3718",x"2e36",x"2153",x"3bf6",x"391f",x"38f3"),
(x"212c",x"3852",x"3716",x"2f15",x"b29c",x"3bc7",x"3921",x"38f1",x"1ba5",x"384b",x"3714",x"2c39",x"a9a5",x"3bf9",x"391a",x"38ee",x"1d2c",x"3850",x"3716",x"2553",x"b2c7",x"3bd1",x"391c",x"38f1"),
(x"212c",x"3852",x"3716",x"2f15",x"b29c",x"3bc7",x"3921",x"38f1",x"2226",x"384e",x"3713",x"291b",x"ab55",x"3bfb",x"3923",x"38ef",x"1ba5",x"384b",x"3714",x"2c39",x"a9a5",x"3bf9",x"391a",x"38ee"),
(x"1f0d",x"383c",x"3713",x"2da1",x"af14",x"3beb",x"391e",x"38e5",x"16e7",x"3832",x"370f",x"2edc",x"acd0",x"3bee",x"3918",x"38e0",x"9aec",x"383c",x"3717",x"30e7",x"b058",x"3bd4",x"3912",x"38e6"),
(x"16e7",x"3832",x"370f",x"2edc",x"acd0",x"3bee",x"3918",x"38e0",x"9631",x"381e",x"3716",x"2adf",x"26b5",x"3bfc",x"3914",x"38d4",x"a039",x"3821",x"3713",x"29b8",x"26e9",x"3bfd",x"390c",x"38d7"),
(x"a12d",x"37d1",x"370d",x"b809",x"ae09",x"3add",x"3907",x"38b7",x"a1a0",x"37df",x"370f",x"b6ca",x"afac",x"3b2e",x"3907",x"38bb",x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4"),
(x"9f80",x"37ae",x"3712",x"a9f0",x"ab1d",x"3bfa",x"390a",x"38ad",x"2043",x"37cb",x"3715",x"99bc",x"26cf",x"3bff",x"391b",x"38b3",x"20de",x"3798",x"3715",x"ad56",x"a0d0",x"3bf8",x"391b",x"38a5"),
(x"1624",x"3809",x"370e",x"3b5f",x"35f1",x"2f4d",x"3955",x"304d",x"17f3",x"380a",x"36eb",x"3b4a",x"3677",x"2cf9",x"3959",x"3053",x"2166",x"37ce",x"36eb",x"3b89",x"3473",x"31fc",x"395b",x"302b"),
(x"235a",x"3925",x"3710",x"bbfd",x"2997",x"a0a8",x"3956",x"28cc",x"22b8",x"3913",x"3713",x"bba5",x"3497",x"ac28",x"3955",x"2918",x"2307",x"3913",x"36eb",x"bba1",x"34cc",x"1f45",x"395a",x"291b"),
(x"234d",x"3931",x"36eb",x"bbf5",x"ae59",x"2467",x"395a",x"289e",x"2325",x"3935",x"3714",x"bbeb",x"b08b",x"98b5",x"3956",x"288b",x"235a",x"3925",x"3710",x"bbfd",x"2997",x"a0a8",x"3956",x"28cc"),
(x"2002",x"38f9",x"3714",x"bb1c",x"3754",x"223f",x"3955",x"298e",x"1c29",x"38ee",x"3718",x"39e5",x"3968",x"0000",x"3954",x"29c8",x"1c29",x"38ee",x"36eb",x"346a",x"3b91",x"316a",x"395a",x"29cb"),
(x"2307",x"3913",x"36eb",x"bba1",x"34cc",x"1f45",x"395a",x"291b",x"22b8",x"3913",x"3713",x"bba5",x"3497",x"ac28",x"3955",x"2918",x"2002",x"38f9",x"3714",x"bb1c",x"3754",x"223f",x"3955",x"298e"),
(x"227e",x"393d",x"3712",x"bb76",x"b5c5",x"204d",x"3956",x"2866",x"2325",x"3935",x"3714",x"bbeb",x"b08b",x"98b5",x"3956",x"288b",x"234d",x"3931",x"36eb",x"bbf5",x"ae59",x"2467",x"395a",x"289e"),
(x"2237",x"3940",x"36eb",x"bab1",x"b862",x"21f0",x"395b",x"285c",x"214b",x"3944",x"3714",x"b95a",x"b9f1",x"2025",x"3956",x"2845",x"227e",x"393d",x"3712",x"bb76",x"b5c5",x"204d",x"3956",x"2866"),
(x"1f6a",x"3948",x"36eb",x"b7e1",x"baf5",x"269a",x"395b",x"2826",x"1f1f",x"3949",x"3714",x"b5bf",x"bb76",x"27db",x"3956",x"2820",x"214b",x"3944",x"3714",x"b95a",x"b9f1",x"2025",x"3956",x"2845"),
(x"142d",x"394c",x"36eb",x"b03c",x"bbeb",x"299b",x"395b",x"27de",x"11db",x"394d",x"3715",x"2836",x"bbfd",x"294f",x"3956",x"27d1",x"1f1f",x"3949",x"3714",x"b5bf",x"bb76",x"27db",x"3956",x"2820"),
(x"9d76",x"3949",x"36eb",x"3868",x"baab",x"296a",x"395b",x"2770",x"9d99",x"394a",x"3716",x"386f",x"baa7",x"2604",x"3956",x"2765",x"11db",x"394d",x"3715",x"2836",x"bbfd",x"294f",x"3956",x"27d1"),
(x"9d76",x"3949",x"36eb",x"3868",x"baab",x"296a",x"395b",x"2770",x"a11a",x"393d",x"36eb",x"3af3",x"b7df",x"2b38",x"395b",x"26eb",x"a14f",x"393d",x"3714",x"3b01",x"b7b5",x"2839",x"3956",x"26e0"),
(x"a1ea",x"3933",x"36eb",x"3bf9",x"ad11",x"2511",x"395b",x"2695",x"a1ee",x"3932",x"3714",x"3be6",x"310f",x"9bfc",x"3956",x"267f",x"a14f",x"393d",x"3714",x"3b01",x"b7b5",x"2839",x"3956",x"26e0"),
(x"a11a",x"3929",x"36eb",x"390c",x"3a34",x"2532",x"395c",x"2642",x"a0ed",x"3929",x"3715",x"3928",x"3a1d",x"1553",x"3956",x"262a",x"a1ee",x"3932",x"3714",x"3be6",x"310f",x"9bfc",x"3956",x"267f"),
(x"a11a",x"3929",x"36eb",x"390c",x"3a34",x"2532",x"395c",x"2642",x"9d99",x"3929",x"36eb",x"b5dd",x"3b6d",x"2be9",x"395c",x"25f5",x"9ddf",x"3928",x"3714",x"afe4",x"3bee",x"28fd",x"3957",x"25e8"),
(x"9d99",x"3929",x"36eb",x"b5dd",x"3b6d",x"2be9",x"395c",x"25f5",x"99c6",x"392e",x"36eb",x"b2b1",x"3bc8",x"2e54",x"395c",x"25b8",x"9908",x"392c",x"3711",x"b64f",x"3b52",x"2d1b",x"3958",x"25a8"),
(x"199d",x"390f",x"36eb",x"3bf6",x"aa70",x"2d61",x"395b",x"2417",x"18c5",x"3910",x"3713",x"3bc2",x"b3a5",x"298a",x"3956",x"2437",x"1b8a",x"3913",x"3711",x"3a7a",x"b8b0",x"283c",x"3957",x"245d"),
(x"99c6",x"392e",x"36eb",x"b2b1",x"3bc8",x"2e54",x"395c",x"25b8",x"1ab2",x"392e",x"36eb",x"337e",x"3bba",x"2ef6",x"395c",x"2550",x"1937",x"392d",x"3710",x"3416",x"3bad",x"2f8d",x"3958",x"2552"),
(x"21a6",x"3888",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b24",x"3a53",x"221a",x"3885",x"3713",x"b583",x"3b63",x"3153",x"3b26",x"3a4f",x"1fdf",x"387c",x"370f",x"ba9b",x"3854",x"30fa",x"3b23",x"3a4e"),
(x"2166",x"37ce",x"36eb",x"3b89",x"3473",x"31fc",x"395b",x"302b",x"2222",x"3797",x"36eb",x"3b99",x"b315",x"330d",x"395c",x"300e",x"20de",x"3798",x"3715",x"3bc5",x"ab9a",x"3358",x"3957",x"300b"),
(x"1de8",x"3919",x"3710",x"2856",x"29ab",x"3bfc",x"391e",x"3963",x"1b8a",x"3913",x"3711",x"340c",x"a6c2",x"3bbc",x"391c",x"3960",x"9a89",x"390e",x"3718",x"2b65",x"3528",x"3b8f",x"3914",x"395d"),
(x"9e52",x"37c7",x"36eb",x"bbe3",x"ace8",x"30c3",x"3955",x"2f4a",x"9f80",x"37ae",x"3712",x"bbcf",x"3081",x"3141",x"3953",x"2f77",x"a0ba",x"37ad",x"36eb",x"bbdb",x"9c67",x"320a",x"3957",x"2f62"),
(x"9e52",x"37c7",x"36eb",x"bbe3",x"ace8",x"30c3",x"3955",x"2f4a",x"9de0",x"37c2",x"3715",x"bbd7",x"31f9",x"2c2a",x"3951",x"2f66",x"9f80",x"37ae",x"3712",x"bbcf",x"3081",x"3141",x"3953",x"2f77"),
(x"a081",x"385d",x"36eb",x"b958",x"b9de",x"2fdf",x"3977",x"28c9",x"a2ed",x"386d",x"36eb",x"bb75",x"b5a2",x"2d46",x"3977",x"287b",x"a294",x"386e",x"3710",x"bb6b",x"b5ba",x"2efe",x"3972",x"287b"),
(x"1e0f",x"392a",x"36eb",x"3aa4",x"3859",x"2fe5",x"395c",x"2513",x"1d11",x"3928",x"3711",x"3a7e",x"3887",x"3089",x"3958",x"2517",x"1937",x"392d",x"3710",x"3416",x"3bad",x"2f8d",x"3958",x"2552"),
(x"990f",x"3909",x"36eb",x"bbe6",x"b08e",x"2c41",x"398e",x"2c46",x"9747",x"3909",x"3718",x"bbe6",x"b09e",x"2baa",x"398a",x"2c2f",x"9613",x"38f6",x"3715",x"bbfa",x"2710",x"2c48",x"3988",x"2c55"),
(x"1e0f",x"392a",x"36eb",x"3aa4",x"3859",x"2fe5",x"395c",x"2513",x"1f98",x"3921",x"36eb",x"3bf4",x"1edc",x"2ebb",x"395c",x"24c5",x"1ea1",x"3921",x"3710",x"3bcc",x"3227",x"2f2f",x"3958",x"24db"),
(x"1e92",x"387d",x"36eb",x"bb7d",x"3521",x"3096",x"3b21",x"3a52",x"1fdf",x"387c",x"370f",x"ba9b",x"3854",x"30fa",x"3b23",x"3a4e",x"2010",x"3876",x"370e",x"bb25",x"b70d",x"2d6a",x"3b22",x"3a4d"),
(x"247a",x"38ba",x"36eb",x"36fe",x"3b25",x"2ea4",x"3997",x"2711",x"2458",x"38b7",x"3714",x"3972",x"39bb",x"30de",x"3992",x"2716",x"2074",x"38bd",x"3711",x"34dc",x"3b97",x"2d60",x"3993",x"27ac"),
(x"1bc8",x"3913",x"36eb",x"39db",x"b96c",x"2c1a",x"395b",x"2439",x"1b8a",x"3913",x"3711",x"3a7a",x"b8b0",x"283c",x"3957",x"245d",x"1de8",x"3919",x"3710",x"3b2f",x"b6d9",x"2e52",x"3957",x"2492"),
(x"1c1b",x"3851",x"36eb",x"b776",x"bb0b",x"2d41",x"3977",x"2941",x"a081",x"385d",x"36eb",x"b958",x"b9de",x"2fdf",x"3977",x"28c9",x"9faa",x"385f",x"3712",x"b84e",x"bab0",x"2ec8",x"3972",x"28c9"),
(x"9943",x"38f3",x"36eb",x"b9df",x"3964",x"2d28",x"398c",x"2c6f",x"989a",x"38f6",x"36eb",x"bbfa",x"20b5",x"2cb4",x"398c",x"2c6a",x"9613",x"38f6",x"3715",x"bbfa",x"2710",x"2c48",x"3988",x"2c55"),
(x"2166",x"386c",x"36eb",x"bad3",x"b822",x"2c4d",x"3b1c",x"3a4f",x"1f2f",x"3877",x"36eb",x"bb19",x"b744",x"2cf7",x"3b1f",x"3a51",x"2010",x"3876",x"370e",x"bb25",x"b70d",x"2d6a",x"3b22",x"3a4d"),
(x"95be",x"381e",x"36eb",x"3bfe",x"9e8d",x"2828",x"3958",x"3068",x"17f3",x"380a",x"36eb",x"3b4a",x"3677",x"2cf9",x"3959",x"3053",x"1624",x"3809",x"370e",x"3b5f",x"35f1",x"2f4d",x"3955",x"304d"),
(x"1c1b",x"3851",x"36eb",x"b776",x"bb0b",x"2d41",x"3977",x"2941",x"1b46",x"3853",x"3716",x"b7e9",x"baf1",x"2aa7",x"3972",x"2932",x"1d2c",x"3850",x"3716",x"bbde",x"b1b6",x"2825",x"3971",x"2944"),
(x"a0ef",x"38e8",x"36eb",x"b9ed",x"394b",x"2f45",x"398a",x"2c92",x"9943",x"38f3",x"36eb",x"b9df",x"3964",x"2d28",x"398c",x"2c6f",x"98e9",x"38f1",x"3715",x"b95d",x"39e3",x"2de3",x"3987",x"2c5d"),
(x"1f03",x"38c0",x"3711",x"3b12",x"3763",x"2ca3",x"3993",x"27d5",x"1e50",x"38c4",x"3712",x"3bf7",x"a83c",x"2d8f",x"3993",x"27f6",x"1f30",x"38c5",x"36eb",x"3bf8",x"2379",x"2d44",x"3997",x"27f5"),
(x"201d",x"38be",x"36eb",x"37d8",x"3af6",x"2a35",x"3997",x"27b6",x"2074",x"38bd",x"3711",x"34dc",x"3b97",x"2d60",x"3993",x"27ac",x"1f03",x"38c0",x"3711",x"3b12",x"3763",x"2ca3",x"3993",x"27d5"),
(x"216e",x"386a",x"36eb",x"b9e9",x"3955",x"2e31",x"3988",x"1d1f",x"2166",x"386c",x"36eb",x"bad3",x"b822",x"2c4d",x"3988",x"1cd9",x"219e",x"386d",x"3713",x"bb5b",x"b634",x"2c03",x"3983",x"1d26"),
(x"95be",x"381e",x"36eb",x"3bfe",x"9e8d",x"2828",x"3958",x"3068",x"9631",x"381e",x"3716",x"3bff",x"a0b5",x"2138",x"3952",x"3062",x"16e7",x"3832",x"370f",x"3ad7",x"b821",x"29e6",x"3952",x"3079"),
(x"1cd4",x"3850",x"36eb",x"bb24",x"371c",x"2cde",x"3977",x"294a",x"1d2c",x"3850",x"3716",x"bbde",x"b1b6",x"2825",x"3971",x"2944",x"1ba5",x"384b",x"3714",x"b9e8",x"3951",x"2f27",x"3972",x"295e"),
(x"a0ef",x"38e8",x"36eb",x"b9ed",x"394b",x"2f45",x"398a",x"2c92",x"9ff6",x"38e8",x"3719",x"b9a6",x"3994",x"2fc6",x"3985",x"2c77",x"9fe7",x"38e6",x"3719",x"b250",x"bbca",x"2f22",x"3985",x"2c7b"),
(x"1f30",x"38c5",x"36eb",x"3bf8",x"2379",x"2d44",x"3997",x"27f5",x"1e50",x"38c4",x"3712",x"3bf7",x"a83c",x"2d8f",x"3993",x"27f6",x"1f3f",x"38cf",x"3712",x"3b92",x"b509",x"2cb0",x"3993",x"2829"),
(x"2072",x"3865",x"3710",x"b833",x"3ac7",x"2d1d",x"3984",x"1e78",x"1ce8",x"3862",x"3713",x"b0a8",x"3bea",x"22dc",x"3984",x"1f99",x"1c5d",x"3862",x"36eb",x"b046",x"3be8",x"2cb7",x"3989",x"1f14"),
(x"216e",x"386a",x"36eb",x"b9e9",x"3955",x"2e31",x"3988",x"1d1f",x"21a8",x"386a",x"3713",x"bb09",x"3791",x"2ab8",x"3983",x"1da7",x"2072",x"3865",x"3710",x"b833",x"3ac7",x"2d1d",x"3984",x"1e78"),
(x"1fba",x"383a",x"36eb",x"373f",x"bb1a",x"2d3c",x"3956",x"308c",x"17ea",x"3831",x"36eb",x"3ab4",x"b859",x"2a66",x"3956",x"307d",x"16e7",x"3832",x"370f",x"3ad7",x"b821",x"29e6",x"3952",x"3079"),
(x"1986",x"384c",x"36eb",x"b97a",x"39b6",x"3099",x"3977",x"2960",x"1ba5",x"384b",x"3714",x"b9e8",x"3951",x"2f27",x"3972",x"295e",x"9aec",x"383c",x"3717",x"ba77",x"3889",x"310e",x"3972",x"29b5"),
(x"9950",x"38e5",x"36eb",x"bb01",x"b745",x"3141",x"3987",x"2cac",x"a09e",x"38e4",x"36eb",x"b2cb",x"bbc1",x"2fc5",x"3989",x"2c99",x"9fe7",x"38e6",x"3719",x"b250",x"bbca",x"2f22",x"3985",x"2c7b"),
(x"1fbf",x"38cd",x"36eb",x"3b57",x"b625",x"2e99",x"3997",x"281d",x"1f3f",x"38cf",x"3712",x"3b92",x"b509",x"2cb0",x"3993",x"2829",x"2353",x"38f1",x"3711",x"3b70",x"b585",x"3014",x"3994",x"28c4"),
(x"11f0",x"3862",x"3712",x"32e8",x"3bcb",x"2c10",x"3985",x"2052",x"9ad5",x"3864",x"3711",x"3934",x"3a0d",x"2c16",x"3986",x"20db",x"9a03",x"3866",x"36eb",x"374a",x"3b15",x"2de4",x"398a",x"2082"),
(x"1c5d",x"3862",x"36eb",x"b046",x"3be8",x"2cb7",x"3989",x"1f14",x"1ce8",x"3862",x"3713",x"b0a8",x"3bea",x"22dc",x"3984",x"1f99",x"11f0",x"3862",x"3712",x"32e8",x"3bcb",x"2c10",x"3985",x"2052"),
(x"1fba",x"383a",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b48",x"3a50",x"1f0d",x"383c",x"3713",x"37c2",x"baf3",x"2e28",x"3b45",x"3a4b",x"2079",x"383b",x"3712",x"b722",x"bb24",x"2bf9",x"3b44",x"3a4c"),
(x"9d26",x"383d",x"36eb",x"baff",x"373c",x"3197",x"3977",x"29bc",x"9aec",x"383c",x"3717",x"ba77",x"3889",x"310e",x"3972",x"29b5",x"a039",x"3821",x"3713",x"bbc6",x"31be",x"30de",x"3972",x"2a2e"),
(x"2422",x"38f3",x"36eb",x"3b99",x"b45f",x"30d6",x"3999",x"28c9",x"2353",x"38f1",x"3711",x"3b70",x"b585",x"3014",x"3994",x"28c4",x"2467",x"3910",x"3711",x"3be4",x"ad1d",x"308c",x"3995",x"294b"),
(x"a09f",x"3872",x"36eb",x"3aaf",x"3860",x"2a70",x"398b",x"2196",x"9a03",x"3866",x"36eb",x"374a",x"3b15",x"2de4",x"398a",x"2082",x"9ad5",x"3864",x"3711",x"3934",x"3a0d",x"2c16",x"3986",x"20db"),
(x"20b1",x"3839",x"36eb",x"b8ae",x"ba73",x"2d49",x"3b47",x"3a50",x"2079",x"383b",x"3712",x"b722",x"bb24",x"2bf9",x"3b44",x"3a4c",x"21e0",x"3837",x"3711",x"b5dd",x"bb65",x"2eae",x"3b43",x"3a4d"),
(x"a0d9",x"3806",x"36eb",x"bbea",x"2e0a",x"2f12",x"3976",x"2aaa",x"a139",x"3821",x"36eb",x"bbbf",x"3113",x"322d",x"3977",x"2a39",x"a039",x"3821",x"3713",x"bbc6",x"31be",x"30de",x"3972",x"2a2e"),
(x"9950",x"38e5",x"36eb",x"bb01",x"b745",x"3141",x"398c",x"2f51",x"9dca",x"38de",x"3715",x"b9d1",x"3974",x"2cc6",x"398f",x"2f7b",x"9fd8",x"38dc",x"36eb",x"ba0e",x"3929",x"2e76",x"3990",x"2f4e"),
(x"9950",x"38e5",x"36eb",x"bb01",x"b745",x"3141",x"398c",x"2f51",x"9920",x"38e4",x"3718",x"baf6",x"37e0",x"2460",x"398d",x"2f80",x"9dca",x"38de",x"3715",x"b9d1",x"3974",x"2cc6",x"398f",x"2f7b"),
(x"24b3",x"3933",x"36eb",x"3be8",x"2d66",x"3010",x"399a",x"29d7",x"24be",x"3910",x"36eb",x"3be6",x"ac77",x"308c",x"3999",x"2946",x"2467",x"3910",x"3711",x"3be4",x"ad1d",x"308c",x"3995",x"294b"),
(x"a166",x"3882",x"36eb",x"3bfa",x"2c62",x"2617",x"398d",x"2295",x"a09f",x"3872",x"36eb",x"3aaf",x"3860",x"2a70",x"398b",x"2196",x"a0d7",x"3872",x"3717",x"3b6f",x"35e4",x"261e",x"3986",x"2216"),
(x"21ab",x"3835",x"36eb",x"ae28",x"bbe6",x"3005",x"3b46",x"3a51",x"21e0",x"3837",x"3711",x"b5dd",x"bb65",x"2eae",x"3b43",x"3a4d",x"23f2",x"3838",x"3712",x"35a6",x"bb63",x"30cc",x"3b41",x"3a4e"),
(x"a0d9",x"3806",x"36eb",x"bbea",x"2e0a",x"2f12",x"3976",x"2aaa",x"a08e",x"3806",x"3717",x"bbf0",x"2f0f",x"2aec",x"3970",x"2a9d",x"a1a0",x"37df",x"370f",x"bbdd",x"30de",x"2e6c",x"3971",x"2afe"),
(x"9fd8",x"38dc",x"36eb",x"ba0e",x"3929",x"2e76",x"3990",x"2f4e",x"9dca",x"38de",x"3715",x"b9d1",x"3974",x"2cc6",x"398f",x"2f7b",x"a0a3",x"38d3",x"3718",x"bb13",x"3732",x"2fec",x"3992",x"2f7c"),
(x"24b3",x"3933",x"36eb",x"3be8",x"2d66",x"3010",x"399a",x"29d7",x"2469",x"3932",x"3714",x"3bec",x"2d02",x"2f4a",x"3995",x"29d9",x"23cf",x"3942",x"3712",x"3b45",x"3640",x"30a6",x"3995",x"2a1c"),
(x"1f98",x"3921",x"36eb",x"3bf4",x"1edc",x"2ebb",x"395c",x"24c5",x"1edf",x"3917",x"36eb",x"3b02",x"b777",x"2fc8",x"395c",x"2477",x"1de8",x"3919",x"3710",x"3b2f",x"b6d9",x"2e52",x"3957",x"2492"),
(x"a0d8",x"3897",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"398e",x"23e2",x"a166",x"3882",x"36eb",x"3bfa",x"2c62",x"2617",x"398d",x"2295",x"a180",x"3883",x"3715",x"3bfe",x"a412",x"2867",x"3988",x"231a"),
(x"244f",x"3835",x"36eb",x"3913",x"ba0d",x"310f",x"3b43",x"3a52",x"23f2",x"3838",x"3712",x"35a6",x"bb63",x"30cc",x"3b41",x"3a4e",x"2498",x"383f",x"3711",x"3bb2",x"b32f",x"30f4",x"3b3f",x"3a4f"),
(x"a243",x"37e1",x"36eb",x"bbe4",x"2adf",x"30ee",x"3975",x"2b06",x"a1a0",x"37df",x"370f",x"bbdd",x"30de",x"2e6c",x"3971",x"2afe",x"a12d",x"37d1",x"370d",x"bb0d",x"b70c",x"3169",x"3971",x"2b1d"),
(x"a164",x"38d4",x"36eb",x"bbbf",x"3333",x"2ed0",x"3992",x"2f4c",x"a0a3",x"38d3",x"3718",x"bb13",x"3732",x"2fec",x"3992",x"2f7c",x"a0f6",x"38cb",x"3712",x"bbf0",x"ac20",x"2e95",x"3994",x"2f75"),
(x"2427",x"3945",x"36eb",x"3ab2",x"3834",x"30cb",x"399a",x"2a24",x"23cf",x"3942",x"3712",x"3b45",x"3640",x"30a6",x"3995",x"2a1c",x"20a5",x"3951",x"3715",x"393c",x"39e9",x"3110",x"3994",x"2a6f"),
(x"9d2f",x"38a7",x"36eb",x"3ac2",x"b833",x"2e8a",x"3990",x"2480",x"a0d8",x"3897",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"398e",x"23e2",x"a123",x"3899",x"3714",x"3b81",x"b558",x"2da5",x"398a",x"243a"),
(x"24ee",x"383f",x"36eb",x"3be5",x"2dbc",x"3036",x"3b40",x"3a53",x"2498",x"383f",x"3711",x"3bb2",x"b32f",x"30f4",x"3b3f",x"3a4f",x"242c",x"384b",x"3712",x"3ae4",x"37c3",x"30c9",x"3b3c",x"3a4f"),
(x"a088",x"37c6",x"36eb",x"b571",x"bb6d",x"30cc",x"3974",x"2b4c",x"a1da",x"37ca",x"36eb",x"baf6",x"b714",x"32f0",x"3975",x"2b36",x"a12d",x"37d1",x"370d",x"bb0d",x"b70c",x"3169",x"3971",x"2b1d"),
(x"a13e",x"38c8",x"36eb",x"bbbf",x"b371",x"2dad",x"3995",x"2f4c",x"a0f6",x"38cb",x"3712",x"bbf0",x"ac20",x"2e95",x"3994",x"2f75",x"a072",x"38c8",x"3712",x"b297",x"bbcc",x"2d84",x"3995",x"2f76"),
(x"20e4",x"3955",x"36eb",x"37cb",x"3ae6",x"3068",x"3999",x"2a7b",x"20a5",x"3951",x"3715",x"393c",x"39e9",x"3110",x"3994",x"2a6f",x"1788",x"3956",x"3715",x"1ef6",x"3bee",x"302a",x"3994",x"2ab0"),
(x"9470",x"38b1",x"36eb",x"39cd",x"b979",x"2caa",x"3991",x"24e4",x"9d2f",x"38a7",x"36eb",x"3ac2",x"b833",x"2e8a",x"3990",x"2480",x"9e13",x"38a8",x"3715",x"3a65",x"b8c1",x"2d9c",x"398b",x"24c4"),
(x"2454",x"384e",x"36eb",x"3902",x"3a23",x"3069",x"3b3c",x"3a54",x"242c",x"384b",x"3712",x"3ae4",x"37c3",x"30c9",x"3b3c",x"3a4f",x"2226",x"384e",x"3713",x"3607",x"3b5e",x"2e4d",x"3b39",x"3a4f"),
(x"9e52",x"37c7",x"36eb",x"bbe3",x"ace8",x"30c3",x"3974",x"2b61",x"a088",x"37c6",x"36eb",x"b571",x"bb6d",x"30cc",x"3974",x"2b4c",x"a05e",x"37cb",x"3713",x"b451",x"bbac",x"2d81",x"3970",x"2b2a"),
(x"9ce6",x"38c7",x"36eb",x"ac58",x"bbf7",x"2bc1",x"3998",x"2f50",x"a0e1",x"38c6",x"36eb",x"aeda",x"bbea",x"2e47",x"3996",x"2f4c",x"a072",x"38c8",x"3712",x"b297",x"bbcc",x"2d84",x"3995",x"2f76"),
(x"9dfd",x"3955",x"36eb",x"b66a",x"3b44",x"2f81",x"3998",x"2b02",x"177f",x"3959",x"36eb",x"16f6",x"3bf5",x"2e99",x"3999",x"2abf",x"1788",x"3956",x"3715",x"1ef6",x"3bee",x"302a",x"3994",x"2ab0"),
(x"11e3",x"38b4",x"36eb",x"b5a5",x"bb74",x"2d53",x"3992",x"2508",x"9470",x"38b1",x"36eb",x"39cd",x"b979",x"2caa",x"3991",x"24e4",x"9607",x"38b2",x"3717",x"3939",x"ba0b",x"29e0",x"398c",x"252b"),
(x"2164",x"3852",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b39",x"3a54",x"21e1",x"3850",x"36eb",x"33f1",x"3bbc",x"2b58",x"3b39",x"3a54",x"2226",x"384e",x"3713",x"3607",x"3b5e",x"2e4d",x"3b39",x"3a4f"),
(x"9de0",x"37c2",x"3715",x"2587",x"b07a",x"3beb",x"390c",x"38b2",x"2043",x"37cb",x"3715",x"99bc",x"26cf",x"3bff",x"391b",x"38b3",x"9f80",x"37ae",x"3712",x"a9f0",x"ab1d",x"3bfa",x"390a",x"38ad"),
(x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4",x"1624",x"3809",x"370e",x"3004",x"271d",x"3bef",x"3916",x"38c8",x"2043",x"37cb",x"3715",x"99bc",x"26cf",x"3bff",x"391b",x"38b3"),
(x"9e25",x"37c9",x"3716",x"20ea",x"2786",x"3bfe",x"390c",x"38b4",x"2043",x"37cb",x"3715",x"99bc",x"26cf",x"3bff",x"391b",x"38b3",x"9de0",x"37c2",x"3715",x"2587",x"b07a",x"3beb",x"390c",x"38b2"),
(x"a08e",x"3806",x"3717",x"2bf6",x"a5ae",x"3bfb",x"390b",x"38c7",x"9631",x"381e",x"3716",x"2adf",x"26b5",x"3bfc",x"3914",x"38d4",x"1624",x"3809",x"370e",x"3004",x"271d",x"3bef",x"3916",x"38c8"),
(x"9ce6",x"38c7",x"36eb",x"ac58",x"bbf7",x"2bc1",x"3998",x"2f50",x"9d58",x"38c8",x"3717",x"aa07",x"bbfc",x"284d",x"3997",x"2f7e",x"9b02",x"38c7",x"3716",x"b8f4",x"ba42",x"2c09",x"3998",x"2f7d"),
(x"a395",x"3947",x"36eb",x"b9f2",x"3938",x"30b5",x"3997",x"2b5e",x"9dfd",x"3955",x"36eb",x"b66a",x"3b44",x"2f81",x"3998",x"2b02",x"9e4d",x"3951",x"3713",x"b82e",x"3aba",x"306c",x"3993",x"2af7"),
(x"1acb",x"38b1",x"3714",x"b9a7",x"b99e",x"2d1e",x"398e",x"2580",x"1e07",x"38ab",x"3714",x"b97e",x"b9c5",x"2dbf",x"398f",x"25bd",x"1e32",x"38a8",x"36eb",x"b976",x"b9cc",x"2dcc",x"3993",x"2580"),
(x"11e3",x"38b4",x"36eb",x"b5a5",x"bb74",x"2d53",x"3992",x"2508",x"125b",x"38b5",x"3717",x"ac93",x"bbf9",x"2918",x"398d",x"2556",x"1acb",x"38b1",x"3714",x"b9a7",x"b99e",x"2d1e",x"398e",x"2580"),
(x"2164",x"3852",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b39",x"3a54",x"212c",x"3852",x"3716",x"3ac7",x"b83c",x"283f",x"3b38",x"3a4f",x"2360",x"3856",x"3711",x"38c8",x"ba4e",x"30a8",x"3b35",x"3a50"),
(x"a493",x"3934",x"36eb",x"bbc4",x"327a",x"3012",x"3995",x"2bae",x"a395",x"3947",x"36eb",x"b9f2",x"3938",x"30b5",x"3997",x"2b5e",x"a2e7",x"3945",x"3715",x"bae0",x"37cf",x"30d4",x"3992",x"2b45"),
(x"1e32",x"38a8",x"36eb",x"b976",x"b9cc",x"2dcc",x"3993",x"2580",x"1e07",x"38ab",x"3714",x"b97e",x"b9c5",x"2dbf",x"398f",x"25bd",x"2116",x"38a4",x"3716",x"b7d5",x"baf0",x"2d8e",x"3990",x"260f"),
(x"2433",x"3855",x"36eb",x"39ec",x"b92b",x"31e4",x"3b35",x"3a55",x"2360",x"3856",x"3711",x"38c8",x"ba4e",x"30a8",x"3b35",x"3a50",x"24fa",x"3866",x"370f",x"3b4b",x"b5cc",x"3223",x"3b30",x"3a51"),
(x"a0ba",x"37ad",x"36eb",x"bbdb",x"9c67",x"320a",x"3957",x"2f62",x"9f80",x"37ae",x"3712",x"bbcf",x"3081",x"3141",x"3953",x"2f77",x"9e24",x"3783",x"370e",x"bb7b",x"b4a9",x"3270",x"3956",x"2f9c"),
(x"9959",x"38c4",x"3715",x"ba5f",x"3873",x"3388",x"396f",x"25f6",x"9abe",x"38bf",x"3714",x"3879",x"b47b",x"3a3d",x"396f",x"261d",x"9ec5",x"38b7",x"3718",x"bac6",x"37dc",x"3286",x"3970",x"2672"),
(x"a46a",x"3921",x"36eb",x"bb6e",x"b575",x"309f",x"3993",x"2bf8",x"a493",x"3934",x"36eb",x"bbc4",x"327a",x"3012",x"3995",x"2bae",x"a44d",x"3933",x"3715",x"bbec",x"2be2",x"2fce",x"3990",x"2b92"),
(x"2002",x"38f9",x"3714",x"305e",x"a1a1",x"3bec",x"3920",x"3951",x"2467",x"3910",x"3711",x"2cd1",x"a504",x"3bf9",x"392a",x"395e",x"2353",x"38f1",x"3711",x"3115",x"a7d5",x"3be4",x"3927",x"394c"),
(x"2002",x"38f9",x"3714",x"305e",x"a1a1",x"3bec",x"3920",x"3951",x"22b8",x"3913",x"3713",x"30f4",x"99bc",x"3be7",x"3926",x"3960",x"2467",x"3910",x"3711",x"2cd1",x"a504",x"3bf9",x"392a",x"395e"),
(x"20ef",x"38a3",x"36eb",x"b53f",x"bb87",x"2d28",x"3994",x"25c5",x"2116",x"38a4",x"3716",x"b7d5",x"baf0",x"2d8e",x"3990",x"260f",x"2323",x"38a3",x"3716",x"2345",x"bbf7",x"2dcc",x"3990",x"2650"),
(x"2563",x"3866",x"36eb",x"3bbc",x"b212",x"3175",x"3b30",x"3a55",x"24fa",x"3866",x"370f",x"3b4b",x"b5cc",x"3223",x"3b30",x"3a51",x"2517",x"3879",x"370f",x"3bd3",x"2f46",x"3182",x"3b2b",x"3a50"),
(x"a0d7",x"38b5",x"36eb",x"bafe",x"375c",x"30f4",x"3975",x"2683",x"9ec5",x"38b7",x"3718",x"bac6",x"37dc",x"3286",x"3970",x"2672",x"a29f",x"389f",x"3714",x"bb6b",x"3587",x"3096",x"3971",x"2754"),
(x"a46a",x"3921",x"36eb",x"bb6e",x"b575",x"309f",x"3993",x"2bf8",x"a409",x"3922",x"3717",x"bb55",x"b5fd",x"307e",x"398e",x"2bd3",x"a18f",x"3914",x"3711",x"b8a4",x"ba69",x"309a",x"398d",x"2c0c"),
(x"2357",x"38a1",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3995",x"2610",x"2323",x"38a3",x"3716",x"2345",x"bbf7",x"2dcc",x"3990",x"2650",x"245f",x"38a6",x"3714",x"3976",x"b9c0",x"3023",x"3991",x"2689"),
(x"2574",x"387a",x"36eb",x"3b61",x"35a0",x"3119",x"3b2b",x"3a55",x"2517",x"3879",x"370f",x"3bd3",x"2f46",x"3182",x"3b2b",x"3a50",x"2437",x"3883",x"370f",x"3891",x"3a72",x"30f5",x"3b28",x"3a50"),
(x"9f92",x"377e",x"36eb",x"bade",x"b7ab",x"31d3",x"395a",x"2f8e",x"9e24",x"3783",x"370e",x"bb7b",x"b4a9",x"3270",x"3956",x"2f9c",x"0f4a",x"3761",x"3712",x"b8b5",x"ba3e",x"32bc",x"3958",x"2fc7"),
(x"a348",x"389f",x"36eb",x"bbba",x"3376",x"2f14",x"3976",x"2750",x"a29f",x"389f",x"3714",x"bb6b",x"3587",x"3096",x"3971",x"2754",x"a3b3",x"3886",x"3712",x"bbf0",x"2a00",x"2f46",x"3972",x"2814"),
(x"9bc5",x"390e",x"36eb",x"b60d",x"bb5a",x"2ef3",x"398f",x"2c3d",x"a22e",x"3911",x"36eb",x"b884",x"ba69",x"3249",x"3991",x"2c1f",x"a18f",x"3914",x"3711",x"b8a4",x"ba69",x"309a",x"398d",x"2c0c"),
(x"24b8",x"38a5",x"36eb",x"3acc",x"b812",x"3064",x"3996",x"265b",x"245f",x"38a6",x"3714",x"3976",x"b9c0",x"3023",x"3991",x"2689",x"24ba",x"38af",x"3712",x"3be0",x"ae5e",x"30a3",x"3992",x"26ce"),
(x"21a6",x"3888",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b24",x"3a53",x"2449",x"3886",x"36eb",x"386e",x"3a87",x"313e",x"3b27",x"3a54",x"2437",x"3883",x"370f",x"3891",x"3a72",x"30f5",x"3b28",x"3a50"),
(x"1dd1",x"3756",x"36eb",x"3996",x"b95f",x"33ec",x"395d",x"2fd5",x"1222",x"3756",x"36eb",x"b8a6",x"ba54",x"3207",x"395d",x"2fc0",x"0f4a",x"3761",x"3712",x"b8b5",x"ba3e",x"32bc",x"3958",x"2fc7"),
(x"a41c",x"3885",x"36eb",x"bbef",x"ad0b",x"2e69",x"3977",x"2816",x"a3b3",x"3886",x"3712",x"bbf0",x"2a00",x"2f46",x"3972",x"2814",x"a294",x"386e",x"3710",x"bb6b",x"b5ba",x"2efe",x"3972",x"287b"),
(x"990f",x"3909",x"36eb",x"bbe6",x"b08e",x"2c41",x"398e",x"2c46",x"9bc5",x"390e",x"36eb",x"b60d",x"bb5a",x"2ef3",x"398f",x"2c3d",x"9a89",x"390e",x"3718",x"b8ae",x"ba78",x"2b7c",x"398a",x"2c25"),
(x"2515",x"38b0",x"36eb",x"3bcf",x"3174",x"303e",x"3997",x"26b6",x"24ba",x"38af",x"3712",x"3be0",x"ae5e",x"30a3",x"3992",x"26ce",x"2458",x"38b7",x"3714",x"3972",x"39bb",x"30de",x"3992",x"2716"),
(x"2467",x"3910",x"3711",x"2cd1",x"a504",x"3bf9",x"392a",x"395e",x"22b8",x"3913",x"3713",x"30f4",x"99bc",x"3be7",x"3926",x"3960",x"235a",x"3925",x"3710",x"a828",x"a60a",x"3bfe",x"3928",x"396a"),
(x"235a",x"3925",x"3710",x"a828",x"a60a",x"3bfe",x"3928",x"396a",x"2469",x"3932",x"3714",x"aeb0",x"a8fa",x"3bf3",x"392b",x"3971",x"2467",x"3910",x"3711",x"2cd1",x"a504",x"3bf9",x"392a",x"395e"),
(x"23cf",x"3942",x"3712",x"2587",x"a08e",x"3bff",x"3929",x"397a",x"2325",x"3935",x"3714",x"a946",x"9ffc",x"3bfe",x"3928",x"3972",x"227e",x"393d",x"3712",x"a953",x"a7ae",x"3bfd",x"3927",x"3977"),
(x"23cf",x"3942",x"3712",x"2587",x"a08e",x"3bff",x"3929",x"397a",x"2469",x"3932",x"3714",x"aeb0",x"a8fa",x"3bf3",x"392b",x"3971",x"2325",x"3935",x"3714",x"a946",x"9ffc",x"3bfe",x"3928",x"3972"),
(x"20a5",x"3951",x"3715",x"20ea",x"aafd",x"3bfc",x"3923",x"3983",x"23cf",x"3942",x"3712",x"2587",x"a08e",x"3bff",x"3929",x"397a",x"214b",x"3944",x"3714",x"28bf",x"ac20",x"3bfa",x"3924",x"397b"),
(x"1788",x"3956",x"3715",x"a7e2",x"a9b2",x"3bfc",x"391c",x"3986",x"20a5",x"3951",x"3715",x"20ea",x"aafd",x"3bfc",x"3923",x"3983",x"1f1f",x"3949",x"3714",x"a31d",x"ab5f",x"3bfc",x"3921",x"397e"),
(x"9e4d",x"3951",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3913",x"3984",x"1788",x"3956",x"3715",x"a7e2",x"a9b2",x"3bfc",x"391c",x"3986",x"11db",x"394d",x"3715",x"a70a",x"2779",x"3bfe",x"391a",x"3981"),
(x"a2e7",x"3945",x"3715",x"2266",x"1d87",x"3bff",x"390b",x"397d",x"9e4d",x"3951",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3913",x"3984",x"9d99",x"394a",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3914",x"397f"),
(x"a44d",x"3933",x"3715",x"288e",x"27ce",x"3bfd",x"3907",x"3973",x"a2e7",x"3945",x"3715",x"2266",x"1d87",x"3bff",x"390b",x"397d",x"a14f",x"393d",x"3714",x"28e0",x"a99e",x"3bfc",x"390e",x"3979"),
(x"a0ed",x"3929",x"3715",x"2c67",x"a8a5",x"3bf9",x"390e",x"396d",x"a409",x"3922",x"3717",x"2d04",x"a793",x"3bf8",x"3907",x"396a",x"a44d",x"3933",x"3715",x"288e",x"27ce",x"3bfd",x"3907",x"3973"),
(x"a18f",x"3914",x"3711",x"28d9",x"252b",x"3bfe",x"390c",x"3962",x"a409",x"3922",x"3717",x"2d04",x"a793",x"3bf8",x"3907",x"396a",x"a0ed",x"3929",x"3715",x"2c67",x"a8a5",x"3bf9",x"390e",x"396d"),
(x"1d11",x"3928",x"3711",x"2bef",x"28a8",x"3bfa",x"391e",x"396c",x"9ddf",x"3928",x"3714",x"2a45",x"ab10",x"3bfa",x"3912",x"396c",x"9908",x"392c",x"3711",x"2a66",x"331a",x"3bca",x"3916",x"396f"),
(x"9a89",x"390e",x"3718",x"2b65",x"3528",x"3b8f",x"3914",x"395d",x"1b8a",x"3913",x"3711",x"340c",x"a6c2",x"3bbc",x"391c",x"3960",x"18c5",x"3910",x"3713",x"341f",x"2c3a",x"3bb6",x"391a",x"395e"),
(x"1832",x"3906",x"3714",x"2de0",x"24c2",x"3bf6",x"391a",x"3958",x"9747",x"3909",x"3718",x"3420",x"9418",x"3bba",x"3916",x"395a",x"18c5",x"3910",x"3713",x"341f",x"2c3a",x"3bb6",x"391a",x"395e"),
(x"1832",x"3906",x"3714",x"2de0",x"24c2",x"3bf6",x"391a",x"3958",x"9613",x"38f6",x"3715",x"27ae",x"24ea",x"3bfe",x"3916",x"394f",x"9747",x"3909",x"3718",x"3420",x"9418",x"3bba",x"3916",x"395a"),
(x"9ddf",x"3928",x"3714",x"2a45",x"ab10",x"3bfa",x"3912",x"396c",x"1de8",x"3919",x"3710",x"2856",x"29ab",x"3bfc",x"391e",x"3963",x"a18f",x"3914",x"3711",x"28d9",x"252b",x"3bfe",x"390c",x"3962"),
(x"1d11",x"3928",x"3711",x"2bef",x"28a8",x"3bfa",x"391e",x"396c",x"1ea1",x"3921",x"3710",x"2a8d",x"a973",x"3bfb",x"391f",x"3968",x"1de8",x"3919",x"3710",x"2856",x"29ab",x"3bfc",x"391e",x"3963"),
(x"1832",x"3906",x"3714",x"3bf3",x"2e23",x"2b27",x"3956",x"23d5",x"18c5",x"3910",x"3713",x"3bc2",x"b3a5",x"298a",x"3956",x"2437",x"199d",x"390f",x"36eb",x"3bf6",x"aa70",x"2d61",x"395b",x"2417"),
(x"1c29",x"38ee",x"36eb",x"346a",x"3b91",x"316a",x"395a",x"2202",x"1c29",x"38ee",x"3718",x"39e5",x"3968",x"0000",x"3954",x"2241",x"1832",x"3906",x"3714",x"3bf3",x"2e23",x"2b27",x"3956",x"23d5"),
(x"b7a8",x"3ca1",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a",x"b783",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b790",x"3ca0",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3107"),
(x"b34f",x"3c93",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20",x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b351",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b368",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b351",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b340",x"3c77",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2a0e"),
(x"b34f",x"3c83",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20",x"b351",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b87d",x"3540",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d",x"b87d",x"3540",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b88f",x"352f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25"),
(x"b441",x"35ca",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19",x"b441",x"35ca",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b40d",x"35e8",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25"),
(x"b4e1",x"3555",x"3710",x"33d2",x"3bc1",x"868d",x"3a87",x"3b28",x"b4e1",x"3555",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4d8",x"354d",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a"),
(x"b568",x"35f7",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21",x"b568",x"35f7",x"36da",x"bb03",x"37b2",x"0000",x"3a97",x"3a21",x"b569",x"3600",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23"),
(x"b88f",x"352f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25",x"b88f",x"352f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b89e",x"351b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b"),
(x"b50c",x"35c6",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3",x"b50c",x"35c6",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b451",x"35c5",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16"),
(x"b4d8",x"354d",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a",x"b4d8",x"354d",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4da",x"3540",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c"),
(x"b84a",x"362a",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01",x"b84a",x"362a",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b83a",x"361d",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa"),
(x"b89e",x"351b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b",x"b89e",x"351b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b8a3",x"3519",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d"),
(x"b451",x"35c5",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16",x"b451",x"35c5",x"36da",x"a987",x"3bfe",x"068d",x"3a54",x"3a16",x"b441",x"35ca",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19"),
(x"b4da",x"3540",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c",x"b4da",x"3540",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4f2",x"3527",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33"),
(x"b85e",x"3620",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09",x"b85e",x"3620",x"36da",x"b5f3",x"3b6d",x"0a8d",x"3be3",x"3a09",x"b84a",x"362a",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01"),
(x"b116",x"35af",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70",x"b116",x"35af",x"36da",x"3bdf",x"31b0",x"8000",x"3a6e",x"3b70",x"b116",x"358c",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77"),
(x"b526",x"35ca",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee",x"b526",x"35ca",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b50c",x"35c6",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3"),
(x"b4f2",x"3527",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33",x"b4f2",x"3527",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f5",x"351a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35"),
(x"b865",x"360e",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e",x"b865",x"360e",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b85e",x"3620",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09"),
(x"b52c",x"35cf",x"3710",x"3bfc",x"ab6c",x"0000",x"3a5f",x"39ec",x"b52c",x"35cf",x"36da",x"3b0d",x"378c",x"0000",x"3a54",x"39ec",x"b526",x"35ca",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee"),
(x"b4f5",x"351a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35",x"b4f5",x"351a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f9",x"350c",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38"),
(x"b867",x"3602",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11",x"b867",x"3602",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b865",x"360e",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e"),
(x"b528",x"35d4",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60",x"b528",x"35d4",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b52c",x"35cf",x"3710",x"3bfc",x"ab6c",x"0000",x"3aa1",x"3a61"),
(x"b4f9",x"350c",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38",x"b4f9",x"350c",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b50d",x"3503",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c"),
(x"b86e",x"35fa",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14",x"b86e",x"35fa",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b867",x"3602",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11"),
(x"b51a",x"35db",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d",x"b51a",x"35db",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b528",x"35d4",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60"),
(x"b50d",x"3503",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c",x"b50d",x"3503",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b52b",x"3507",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42"),
(x"b87d",x"35fb",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a",x"b87d",x"35fb",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b86e",x"35fa",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14"),
(x"b4e1",x"35e6",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52",x"b4e1",x"35e6",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b51a",x"35db",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d"),
(x"b52b",x"3507",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42",x"b52b",x"3507",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b544",x"3511",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47"),
(x"b88f",x"360c",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22",x"b88f",x"360c",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b87d",x"35fb",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a"),
(x"b4d8",x"35ef",x"3710",x"3be5",x"b11d",x"0000",x"3aa1",x"3a50",x"b4d8",x"35ef",x"36da",x"3af9",x"b7d7",x"8000",x"3a97",x"3a50",x"b4e1",x"35e6",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52"),
(x"b544",x"3511",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47",x"b544",x"3511",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b558",x"3511",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b"),
(x"b89e",x"3620",x"3710",x"36ef",x"3b35",x"0000",x"3bd9",x"3a29",x"b89e",x"3620",x"36da",x"380f",x"3ae4",x"8000",x"3be3",x"3a29",x"b88f",x"360c",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22"),
(x"b4da",x"35fb",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d",x"b4da",x"35fb",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4d8",x"35ef",x"3710",x"3be5",x"b11d",x"0000",x"3aa1",x"3a50"),
(x"b558",x"3511",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b",x"b558",x"3511",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b568",x"3518",x"3710",x"b810",x"bae4",x"8000",x"3a87",x"3b4e"),
(x"b8a3",x"3622",x"3710",x"286a",x"3bfe",x"868d",x"3bd9",x"3a2b",x"b8a3",x"3622",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b89e",x"3620",x"3710",x"36ef",x"3b35",x"0000",x"3bd9",x"3a29"),
(x"b4f2",x"3615",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47",x"b4f2",x"3615",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4da",x"35fb",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d"),
(x"b568",x"3544",x"3710",x"bb03",x"b7b2",x"0000",x"3a87",x"3b59",x"b568",x"3544",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b581",x"355c",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f"),
(x"b8ff",x"3627",x"3710",x"2581",x"3bff",x"1553",x"3bd9",x"3a4f",x"b8ff",x"3627",x"36da",x"26a7",x"3bff",x"8000",x"3be3",x"3a4f",x"b8a3",x"3622",x"3710",x"286a",x"3bfe",x"868d",x"3bd9",x"3a2b"),
(x"b931",x"35cd",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4",x"b931",x"35cd",x"36da",x"bbff",x"a4d0",x"0000",x"3a18",x"33f3",x"b931",x"3629",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9"),
(x"b4f5",x"3621",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44",x"b4f5",x"3621",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f2",x"3615",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47"),
(x"b581",x"355c",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f",x"b581",x"355c",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b5a1",x"3568",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66"),
(x"b4f9",x"362f",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41",x"b4f9",x"362f",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f5",x"3621",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44"),
(x"b5a1",x"3568",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66",x"b5a1",x"3568",x"36da",x"b72d",x"bb26",x"0000",x"3a7c",x"3b66",x"b5bd",x"3578",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c"),
(x"b50d",x"3638",x"3710",x"2546",x"3bff",x"068d",x"3aa1",x"3a3d",x"b50d",x"3638",x"36da",x"324b",x"3bd8",x"0000",x"3a97",x"3a3d",x"b4f9",x"362f",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41"),
(x"b5bd",x"3578",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c",x"b5bd",x"3578",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5ce",x"357b",x"3710",x"2aec",x"bbfc",x"0000",x"3a87",x"3b6f"),
(x"b52b",x"3634",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37",x"b52b",x"3634",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b50d",x"3638",x"3710",x"2546",x"3bff",x"068d",x"3aa1",x"3a3d"),
(x"b5ce",x"357b",x"3710",x"2aec",x"bbfc",x"0000",x"3a87",x"3b6f",x"b5ce",x"357b",x"36da",x"2f27",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b62a",x"356e",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81"),
(x"b544",x"362a",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32",x"b544",x"362a",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b52b",x"3634",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37"),
(x"b575",x"3526",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52",x"b575",x"3526",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3530",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54"),
(x"b558",x"362a",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f",x"b558",x"362a",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b544",x"362a",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32"),
(x"b62a",x"356e",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81",x"b62a",x"356e",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b63d",x"356c",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84"),
(x"b568",x"3623",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b",x"b568",x"3623",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b558",x"362a",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f"),
(x"b63d",x"356c",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84",x"b63d",x"356c",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b669",x"3574",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d"),
(x"b8a3",x"3519",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d",x"b8a3",x"3519",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b906",x"3513",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53"),
(x"b581",x"35e0",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a",x"b581",x"35e0",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b568",x"35f7",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21"),
(x"b669",x"3574",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d",x"b669",x"3574",x"36da",x"a666",x"bbff",x"0000",x"3a7c",x"3b8d",x"b721",x"3575",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf"),
(x"b5a1",x"35d3",x"3710",x"b72d",x"3b26",x"0000",x"3aa1",x"3a14",x"b5a1",x"35d3",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b581",x"35e0",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a"),
(x"b568",x"3518",x"3710",x"b810",x"bae4",x"8000",x"3a87",x"3b4e",x"b568",x"3518",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b575",x"3526",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52"),
(x"b116",x"358c",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77",x"b116",x"358c",x"36da",x"3b51",x"b675",x"8000",x"3a6e",x"3b77",x"b135",x"357a",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b"),
(x"b93a",x"35c9",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"3861",x"b93a",x"35c9",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"385a",x"b931",x"35cd",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b5bd",x"35c3",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e",x"b5bd",x"35c3",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5a1",x"35d3",x"3710",x"b72d",x"3b26",x"0000",x"3aa1",x"3a14"),
(x"b721",x"3575",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf",x"b721",x"3575",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b72d",x"3572",x"3710",x"3778",x"bb13",x"0000",x"3a87",x"3bb2"),
(x"b135",x"357a",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b",x"b135",x"357a",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b161",x"3571",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80"),
(x"b5ce",x"35c0",x"3710",x"2f27",x"3bf3",x"0000",x"3aa1",x"3a0b",x"b5ce",x"35c0",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5bd",x"35c3",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e"),
(x"b72d",x"3572",x"3710",x"3778",x"bb13",x"0000",x"3a95",x"39fb",x"b72d",x"3572",x"36da",x"3a45",x"b8f8",x"0000",x"3a8a",x"39fb",x"b72e",x"356a",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd"),
(x"b161",x"3571",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80",x"b161",x"3571",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b1a1",x"356f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86"),
(x"b62a",x"35cd",x"3710",x"2fb9",x"3bf1",x"0000",x"3aa1",x"39f9",x"b62a",x"35cd",x"36da",x"303a",x"3bed",x"8000",x"3a97",x"39f9",x"b5ce",x"35c0",x"3710",x"2f27",x"3bf3",x"0000",x"3aa1",x"3a0b"),
(x"b72e",x"356a",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd",x"b72e",x"356a",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b721",x"3562",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00"),
(x"b1a1",x"356f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86",x"b1a1",x"356f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1c1",x"356b",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89"),
(x"b575",x"360b",x"3710",x"ba67",x"b8cb",x"868d",x"3aa1",x"3a26",x"b575",x"360b",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"3615",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28"),
(x"b721",x"3562",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00",x"b721",x"3562",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b6fb",x"3550",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08"),
(x"b906",x"3513",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53",x"b906",x"3513",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b931",x"3514",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63"),
(x"b1c1",x"356b",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89",x"b1c1",x"356b",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1fd",x"3558",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90"),
(x"b63d",x"35cf",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5",x"b63d",x"35cf",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b62a",x"35cd",x"3710",x"2fb9",x"3bf1",x"0000",x"3aa1",x"39f9"),
(x"b6fb",x"3550",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08",x"b6fb",x"3550",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6ef",x"3541",x"3710",x"3b57",x"3658",x"868d",x"3a95",x"3a0c"),
(x"b1fd",x"3558",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90",x"b1fd",x"3558",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b22d",x"3552",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94"),
(x"b906",x"3513",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53",x"b931",x"3514",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63",x"b90c",x"3513",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55"),
(x"b90c",x"3513",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55",x"b92b",x"3513",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b912",x"3513",x"373c",x"184d",x"bbff",x"26c8",x"3a8e",x"3a57"),
(x"b912",x"3513",x"373c",x"184d",x"bbff",x"26c8",x"3a8e",x"3a57",x"b924",x"3514",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b918",x"3514",x"374b",x"2511",x"bbff",x"2259",x"3a91",x"3a59"),
(x"b8ff",x"3627",x"3710",x"257a",x"3bff",x"15bc",x"3bd9",x"3a4f",x"b907",x"3627",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b931",x"3629",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63"),
(x"b907",x"3627",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b90b",x"3627",x"3722",x"2773",x"3bfe",x"22dc",x"3bd6",x"3a54",x"b92f",x"3629",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62"),
(x"b90b",x"3627",x"3722",x"2773",x"3bfe",x"22dc",x"3bd6",x"3a54",x"b911",x"3628",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b92c",x"3629",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60"),
(x"b911",x"3628",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b918",x"3627",x"374b",x"270a",x"3bfd",x"287a",x"3bce",x"3a59",x"b925",x"3628",x"3749",x"257a",x"3bfd",x"28f7",x"3bcf",x"3a5e"),
(x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b8a3",x"3519",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b906",x"3513",x"3710",x"2e12",x"a66c",x"3bf6",x"39f2",x"333e"),
(x"b907",x"3627",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340",x"b8ff",x"3627",x"3710",x"2904",x"26d5",x"3bfd",x"3a2d",x"3331",x"b906",x"35cc",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d"),
(x"b906",x"35cc",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b8a3",x"3622",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b8a3",x"3519",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b8a3",x"3622",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b89e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b89e",x"3620",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3284",x"b88f",x"360c",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b89e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b88f",x"352f",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"3269",x"b88f",x"360c",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b87d",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248"),
(x"b87d",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248",x"b87d",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b86e",x"3541",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b86e",x"35fa",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"322d",x"b867",x"3602",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b86e",x"3541",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b867",x"3539",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"3222",x"b867",x"3602",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b865",x"352d",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d"),
(x"b865",x"352d",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d",x"b865",x"360e",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b85e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211"),
(x"b85e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211",x"b85e",x"3620",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b84a",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"b84a",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed",x"b84a",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b83a",x"351e",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b83a",x"361d",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"31d0",x"b820",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b83a",x"351e",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b820",x"3554",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"31a2",x"b820",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b801",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b"),
(x"b801",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b",x"b801",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b7c0",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130"),
(x"b77b",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b783",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b72e",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b783",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b77b",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b72e",x"356a",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae"),
(x"b77b",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b72e",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae",x"b776",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b72d",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b72e",x"356a",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b776",x"355b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"b783",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b7a4",x"351f",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7a8",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a"),
(x"b7bd",x"35ff",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d",x"b7a4",x"361c",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b7a8",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a"),
(x"b7c7",x"3608",x"3710",x"8000",x"0000",x"3c00",x"3a26",x"3136",x"b7c7",x"360d",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3135",x"b7bd",x"35ff",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d"),
(x"b7a4",x"351f",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7c7",x"352e",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3135",x"b7bd",x"353c",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d"),
(x"b783",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b72e",x"356a",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b73e",x"350e",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"b783",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b73e",x"362d",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b72e",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b73e",x"362d",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b705",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b721",x"35da",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"b705",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b6f1",x"3610",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"3076",x"b6fb",x"35eb",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080"),
(x"b73e",x"350e",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc",x"b721",x"3562",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b705",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088"),
(x"b705",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088",x"b6fb",x"3550",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b6f1",x"352c",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3076"),
(x"b72d",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b776",x"355b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b72d",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"b776",x"355b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b77a",x"3565",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b776",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b77a",x"3565",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b794",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b77a",x"35d6",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"b794",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"3109",x"b794",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b7c0",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130"),
(x"b72d",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"30ad",x"b72d",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b721",x"3575",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b721",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30a2",x"b669",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b721",x"3575",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b669",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2ffc",x"b669",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b63d",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"b63d",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac",x"b63d",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b62a",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"b568",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30",x"b568",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b52c",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"b526",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2dbb",x"b526",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb",x"b52c",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"b52c",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5",x"b528",x"3567",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b568",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b569",x"3600",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33",x"b528",x"35d4",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b568",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"b4f2",x"3527",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b544",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b528",x"3567",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"b4f2",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e",x"b528",x"35d4",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b544",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"b4da",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33",x"b51a",x"35db",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b4f2",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b528",x"3567",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b51a",x"3560",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4f2",x"3527",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"b51a",x"3560",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4e1",x"3555",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"2d40",x"b4da",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"b4d8",x"35ef",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2d2f",x"b4e1",x"35e6",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2d40",x"b4da",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"b575",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47",x"b558",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b569",x"3600",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"b575",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2e49",x"b568",x"3623",x"3710",x"8000",x"0000",x"3c00",x"3a2c",x"2e32",x"b575",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"b544",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b558",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b569",x"353b",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"b558",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b568",x"3518",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2e32",x"b575",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"b544",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b4f2",x"3527",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b52b",x"3507",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"b52b",x"3507",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4",x"b4f5",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b50d",x"3503",x"3710",x"8000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"b544",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0",x"b52b",x"3634",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b4f2",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b52b",x"3634",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b50d",x"3638",x"3710",x"8000",x"0000",x"3c00",x"3a30",x"2d8e",x"b4f5",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"b581",x"355c",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2e5e",x"b581",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e",x"b568",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b581",x"355c",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2e5e",x"b5a1",x"3568",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b581",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"b5a1",x"3568",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b5bd",x"3578",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9",x"b5a1",x"35d3",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"b5ce",x"357b",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2ee7",x"b5ce",x"35c0",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7",x"b5bd",x"3578",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"b5ce",x"357b",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2ee7",x"b62a",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b",x"b5ce",x"35c0",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"b526",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2dbb",x"b50c",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d",x"b526",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"b368",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b340",x"35ee",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"2a04",x"b351",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b407",x"35f1",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76",x"b3a5",x"3610",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b368",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b3a5",x"352b",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b3a5",x"352b",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b3d2",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b407",x"354a",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"b3d2",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b3f4",x"352a",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b409",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"b3f4",x"352a",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b40b",x"3528",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b84",x"b413",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"b409",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d",x"b3d2",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b407",x"35f1",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"b413",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0",x"b3f4",x"3612",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b409",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"b413",x"360e",x"3710",x"068d",x"0000",x"3c00",x"3a27",x"2ba0",x"b40b",x"3613",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b84",x"b413",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"b34f",x"357c",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20",x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b34f",x"35bf",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b441",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b441",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b451",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b441",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"b451",x"35c5",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2c3f",x"b451",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b50c",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"b34f",x"35bf",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20",x"b326",x"35bd",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b34f",x"357c",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"b326",x"35bd",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b2d6",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b326",x"357e",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"b2d6",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b2aa",x"35cd",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b2d6",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949"),
(x"b2aa",x"35cd",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b261",x"35e2",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b2aa",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"b261",x"35e2",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b22d",x"35e9",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a",x"b261",x"3559",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878"),
(x"b1fd",x"35e3",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"278b",x"b1fd",x"3558",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b",x"b22d",x"35e9",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"b1fd",x"35e3",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"278b",x"b1c1",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3",x"b1fd",x"3558",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b"),
(x"b1a1",x"35cc",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2643",x"b1a1",x"356f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643",x"b1c1",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"b1a1",x"35cc",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2643",x"b161",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b1a1",x"356f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643"),
(x"b161",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b135",x"35c1",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b161",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f"),
(x"b135",x"35c1",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b116",x"35af",x"3710",x"8000",x"0000",x"3c00",x"3a13",x"2451",x"b135",x"357a",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"b906",x"35cc",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b90b",x"35ce",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b907",x"3627",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340"),
(x"b90b",x"35ce",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b913",x"35cf",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b90b",x"3627",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c"),
(x"b911",x"3628",x"373c",x"3ac9",x"a6b5",x"383a",x"3a2d",x"3366",x"b913",x"35cf",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b918",x"3627",x"374b",x"38ec",x"a7f6",x"3a4c",x"3a2d",x"3378"),
(x"b918",x"3627",x"374b",x"38ec",x"a7f6",x"3a4c",x"3a2d",x"3378",x"b919",x"35cf",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b91f",x"3628",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385"),
(x"b91f",x"3628",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385",x"b920",x"35ce",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b925",x"3628",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b925",x"35ce",x"3746",x"b918",x"a84d",x"3a28",x"3a1a",x"338e",x"b92a",x"35ce",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b925",x"3628",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b92a",x"35ce",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b92f",x"3629",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b92c",x"3629",x"373a",x"baa5",x"a5fd",x"3872",x"3a2d",x"33a3"),
(x"b931",x"3629",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9",x"b92f",x"3629",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b931",x"35cd",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4"),
(x"b90e",x"3574",x"370e",x"b4eb",x"a6e9",x"3b9c",x"3a06",x"334b",x"b90d",x"35c9",x"3711",x"b36d",x"a40b",x"3bc7",x"3a19",x"3349",x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b906",x"35cc",x"3713",x"2edc",x"bb7b",x"3565",x"3b16",x"387a",x"b90d",x"35c9",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"387b",x"b90b",x"35ce",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879"),
(x"b90b",x"35ce",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879",x"b90d",x"35c9",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"387b",x"b90f",x"35c9",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879"),
(x"b90b",x"35ce",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3879",x"b90f",x"35c9",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879",x"b913",x"35cf",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875"),
(x"b913",x"35cf",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875",x"b913",x"35c8",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b919",x"35cf",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873"),
(x"b919",x"35cf",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873",x"b91a",x"35c8",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b920",x"35ce",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871"),
(x"b920",x"35ce",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871",x"b922",x"35c8",x"3751",x"9a8d",x"39ac",x"39a3",x"3b24",x"3871",x"b928",x"35c8",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e"),
(x"b920",x"35ce",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871",x"b928",x"35c8",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e",x"b925",x"35ce",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e"),
(x"b925",x"35ce",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e",x"b92f",x"35c8",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b92a",x"35ce",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"386b"),
(x"b92a",x"35ce",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"386b",x"b935",x"35c8",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b931",x"35cd",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b92a",x"356e",x"3733",x"b800",x"ba99",x"3437",x"3bb7",x"3993",x"b930",x"3577",x"3738",x"b75b",x"bae5",x"32d3",x"3bb5",x"3992",x"b92b",x"3577",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b924",x"3577",x"374d",x"b1ce",x"b808",x"3ac1",x"3bb5",x"3999",x"b922",x"356e",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998",x"b92b",x"3577",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b924",x"3577",x"374d",x"b1ce",x"b808",x"3ac1",x"3bb5",x"3999",x"b91b",x"3577",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b922",x"356e",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998"),
(x"b912",x"3513",x"373c",x"3aea",x"2832",x"3802",x"39f2",x"336a",x"b918",x"3514",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b",x"b913",x"356e",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369"),
(x"b938",x"3576",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a",x"b930",x"3577",x"3738",x"b75b",x"bae5",x"32d3",x"3bb5",x"3992",x"b930",x"356e",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c"),
(x"b935",x"35c8",x"3725",x"bb50",x"a638",x"3678",x"3be8",x"39de",x"b938",x"3576",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b93a",x"35c9",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3be8",x"39da"),
(x"b938",x"3576",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b935",x"35c8",x"3725",x"bb50",x"a638",x"3678",x"3be8",x"39de",x"b930",x"3577",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3"),
(x"b930",x"3577",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3",x"b92f",x"35c8",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b92b",x"3577",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6"),
(x"b92b",x"3577",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6",x"b928",x"35c8",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b924",x"3577",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b922",x"35c8",x"3751",x"a11e",x"aa52",x"3bfd",x"3be8",x"39eb",x"b91a",x"35c8",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b924",x"3577",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b91a",x"35c8",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b913",x"35c8",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b91b",x"3577",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed"),
(x"b90f",x"35c9",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7",x"b90d",x"35c9",x"3711",x"3be1",x"a6cf",x"3179",x"3be9",x"39fb",x"b90e",x"3574",x"370e",x"3bcb",x"a949",x"330f",x"3bf9",x"39fa"),
(x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b906",x"3513",x"3710",x"2e12",x"a66c",x"3bf6",x"39f2",x"333e",x"b90c",x"3513",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352"),
(x"b91b",x"3577",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b913",x"3575",x"373a",x"3ae3",x"2b4b",x"380a",x"3bb9",x"399f",x"b91b",x"356e",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b"),
(x"b907",x"3571",x"3713",x"2f5f",x"3bdb",x"30c1",x"3bc0",x"39a6",x"b913",x"356e",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b90e",x"3574",x"370e",x"3754",x"3ae5",x"32eb",x"3bbd",x"39a7"),
(x"b91f",x"3513",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387",x"b91b",x"356e",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b918",x"3514",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b"),
(x"b924",x"3514",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392",x"b922",x"356e",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b91f",x"3513",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387"),
(x"b92b",x"3513",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa",x"b92a",x"356e",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b924",x"3514",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392"),
(x"b931",x"3514",x"3710",x"bbe9",x"26a1",x"309e",x"39f4",x"33ca",x"b930",x"356e",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0",x"b92b",x"3513",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa"),
(x"b83a",x"361d",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa",x"b83a",x"361d",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b820",x"35e8",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec"),
(x"b51a",x"3560",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d",x"b51a",x"3560",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b4e1",x"3555",x"3710",x"33d2",x"3bc1",x"868d",x"3a87",x"3b28"),
(x"b40d",x"35e8",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25",x"b40d",x"35e8",x"36da",x"b8bf",x"3a70",x"868d",x"3a54",x"3a25",x"b407",x"35f1",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27"),
(x"b86e",x"3541",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17",x"b86e",x"3541",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b87d",x"3540",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d"),
(x"b569",x"3600",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23",x"b569",x"3600",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b575",x"360b",x"3710",x"ba67",x"b8cb",x"868d",x"3aa1",x"3a26"),
(x"b528",x"3567",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a",x"b528",x"3567",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b51a",x"3560",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d"),
(x"b407",x"35f1",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27",x"b407",x"35f1",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b409",x"35f7",x"3710",x"bb1a",x"b75d",x"8000",x"3a5f",x"3a28"),
(x"b867",x"3539",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14",x"b867",x"3539",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b86e",x"3541",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17"),
(x"b820",x"35e8",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec",x"b820",x"35e8",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b801",x"35ca",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de"),
(x"b52c",x"356c",x"3710",x"3b0d",x"b78c",x"0000",x"3a87",x"3b19",x"b52c",x"356c",x"36da",x"3bfc",x"2b6c",x"0000",x"3a7c",x"3b19",x"b528",x"3567",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a"),
(x"b409",x"35f7",x"3710",x"bb1a",x"b75d",x"8000",x"3a5f",x"3a28",x"b409",x"35f7",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b413",x"3605",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b"),
(x"b865",x"352d",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12",x"b865",x"352d",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b867",x"3539",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14"),
(x"b801",x"35ca",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de",x"b801",x"35ca",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b7c0",x"35c2",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1"),
(x"b526",x"3571",x"3710",x"33bb",x"bbc3",x"0000",x"3b06",x"3a0f",x"b526",x"3571",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b52c",x"356c",x"3710",x"3b0d",x"b78c",x"0000",x"3b06",x"3a11"),
(x"b413",x"3605",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b",x"b413",x"3605",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"360e",x"3710",x"bb8c",x"354a",x"0000",x"3a5f",x"3a2d"),
(x"b85e",x"351b",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d",x"b85e",x"351b",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b865",x"352d",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12"),
(x"b7c0",x"35c2",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1",x"b7c0",x"35c2",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b794",x"35c9",x"3710",x"b357",x"3bc9",x"0000",x"3bd9",x"39c8"),
(x"b50c",x"3576",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a",x"b50c",x"3576",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b526",x"3571",x"3710",x"33bb",x"bbc3",x"0000",x"3b06",x"3a0f"),
(x"b413",x"360e",x"3710",x"bb8c",x"354a",x"0000",x"3a5f",x"3a2d",x"b413",x"360e",x"36da",x"ba12",x"3935",x"068d",x"3a54",x"3a2d",x"b40b",x"3613",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e"),
(x"b84a",x"3511",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05",x"b84a",x"3511",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b85e",x"351b",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d"),
(x"b794",x"35c9",x"3710",x"b357",x"3bc9",x"0000",x"3bd9",x"39c8",x"b794",x"35c9",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b77a",x"35d6",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2"),
(x"b441",x"3571",x"3710",x"b7a4",x"bb07",x"0000",x"3b06",x"39e4",x"b441",x"3571",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b451",x"3576",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7"),
(x"b40b",x"3613",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e",x"b40b",x"3613",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b3f4",x"3612",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32"),
(x"b83a",x"351e",x"3710",x"3953",x"b9f7",x"868d",x"3a85",x"39ff",x"b83a",x"351e",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b84a",x"3511",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05"),
(x"b77a",x"35d6",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2",x"b77a",x"35d6",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b776",x"35e0",x"3710",x"bbee",x"3038",x"0000",x"3bd9",x"39c0"),
(x"b451",x"3576",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7",x"b451",x"3576",x"36da",x"a0ea",x"bc00",x"0000",x"3afb",x"39e7",x"b50c",x"3576",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a"),
(x"b3f4",x"3612",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32",x"b3f4",x"3612",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3d2",x"360b",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35"),
(x"b569",x"353b",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57",x"b569",x"353b",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b568",x"3544",x"3710",x"bb03",x"b7b2",x"0000",x"3a87",x"3b59"),
(x"b776",x"35e0",x"3710",x"bbee",x"3038",x"0000",x"3bd9",x"39c0",x"b776",x"35e0",x"36da",x"bbce",x"b2fb",x"0000",x"3be3",x"39c0",x"b77b",x"35e8",x"3710",x"b937",x"ba10",x"0000",x"3bd9",x"39be"),
(x"b40d",x"3553",x"3710",x"b8bf",x"ba70",x"8000",x"3b06",x"39d8",x"b40d",x"3553",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b441",x"3571",x"3710",x"b7a4",x"bb07",x"0000",x"3b06",x"39e4"),
(x"b3d2",x"360b",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35",x"b3d2",x"360b",x"36da",x"abf6",x"3bfc",x"0000",x"3a54",x"3a35",x"b3a5",x"3610",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39"),
(x"b820",x"3554",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1",x"b820",x"3554",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b83a",x"351e",x"3710",x"3953",x"b9f7",x"868d",x"3a85",x"39ff"),
(x"b77b",x"35e8",x"3710",x"b937",x"ba10",x"0000",x"3a87",x"3ac5",x"b77b",x"35e8",x"36da",x"b853",x"baba",x"0000",x"3a7d",x"3ac5",x"b790",x"35f3",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9"),
(x"b407",x"354a",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6",x"b407",x"354a",x"36da",x"bb61",x"b629",x"0000",x"3afb",x"39d6",x"b40d",x"3553",x"3710",x"b8bf",x"ba70",x"8000",x"3b06",x"39d8"),
(x"b3a5",x"3610",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39",x"b3a5",x"3610",x"36da",x"32b5",x"3bd2",x"8000",x"3a54",x"3a39",x"b368",x"3605",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40"),
(x"b575",x"3530",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54",x"b575",x"3530",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b569",x"353b",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57"),
(x"b790",x"35f3",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9",x"b790",x"35f3",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b7a8",x"35f7",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace"),
(x"b409",x"3544",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5",x"b409",x"3544",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b407",x"354a",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6"),
(x"b368",x"3605",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40",x"b368",x"3605",x"36da",x"3912",x"3a2f",x"8000",x"3a54",x"3a40",x"b340",x"35ee",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45"),
(x"b801",x"3572",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4",x"b801",x"3572",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b820",x"3554",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1"),
(x"b7a8",x"35f7",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace",x"b7a8",x"35f7",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7bd",x"35ff",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2"),
(x"b413",x"3536",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2",x"b413",x"3536",x"36da",x"bb08",x"37a1",x"868d",x"3afb",x"39d2",x"b409",x"3544",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5"),
(x"b340",x"35ee",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45",x"b340",x"35ee",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b33a",x"35d9",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49"),
(x"b7c0",x"3579",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7",x"b7c0",x"3579",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b801",x"3572",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4"),
(x"b7bd",x"35ff",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2",x"b7bd",x"35ff",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7c7",x"3608",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5"),
(x"b931",x"3514",x"3710",x"bbe9",x"26a1",x"309e",x"39f4",x"33ca",x"b931",x"3514",x"36da",x"bbff",x"26b5",x"0000",x"39f5",x"33fa",x"b930",x"356e",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0"),
(x"b413",x"352d",x"3710",x"ba12",x"b935",x"868d",x"3b06",x"39d0",x"b413",x"352d",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"3536",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2"),
(x"b33a",x"35d9",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49",x"b33a",x"35d9",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b351",x"35c7",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d"),
(x"b794",x"3572",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf",x"b794",x"3572",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b7c0",x"3579",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7"),
(x"b7c7",x"3608",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5",x"b7c7",x"3608",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"360d",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6"),
(x"b40b",x"3528",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce",x"b40b",x"3528",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b413",x"352d",x"3710",x"ba12",x"b935",x"868d",x"3b06",x"39d0"),
(x"b351",x"35c7",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d",x"b351",x"35c7",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b34f",x"35bf",x"3710",x"3913",x"3a2f",x"0000",x"3a5f",x"3a4f"),
(x"b77a",x"3565",x"3710",x"b97c",x"b9d2",x"0000",x"3a85",x"39c9",x"b77a",x"3565",x"36da",x"b83f",x"bac7",x"0000",x"3a7b",x"39c9",x"b794",x"3572",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf"),
(x"b7c7",x"360d",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6",x"b7c7",x"360d",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7a4",x"361c",x"3710",x"b655",x"3b58",x"8000",x"3a87",x"3add"),
(x"b3f4",x"352a",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb",x"b3f4",x"352a",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b40b",x"3528",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce"),
(x"b34f",x"35bf",x"3710",x"3913",x"3a2f",x"0000",x"3a79",x"3b35",x"b34f",x"35bf",x"36da",x"3448",x"3bb5",x"0000",x"3a6e",x"3b35",x"b326",x"35bd",x"3710",x"a5e3",x"3bff",x"0000",x"3a79",x"3b39"),
(x"b776",x"355b",x"3710",x"bbce",x"32fc",x"0000",x"3a95",x"3a4d",x"b776",x"355b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b77a",x"3565",x"3710",x"b97c",x"b9d2",x"0000",x"3a95",x"3a50"),
(x"b7a4",x"361c",x"3710",x"b655",x"3b58",x"8000",x"3a87",x"3add",x"b7a4",x"361c",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b783",x"362a",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4"),
(x"b3d2",x"3530",x"3710",x"abf6",x"bbfc",x"0000",x"3b06",x"39c8",x"b3d2",x"3530",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3f4",x"352a",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb"),
(x"b326",x"35bd",x"3710",x"a5e3",x"3bff",x"0000",x"3a79",x"3b39",x"b326",x"35bd",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b2d6",x"35c2",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41"),
(x"b77b",x"3553",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c",x"b77b",x"3553",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b776",x"355b",x"3710",x"bbce",x"32fc",x"0000",x"3a95",x"3a4d"),
(x"b783",x"362a",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4",x"b783",x"362a",x"36da",x"afa0",x"3bf1",x"068d",x"3a7d",x"3ae4",x"b73e",x"362d",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1"),
(x"b3a5",x"352b",x"3710",x"32b5",x"bbd2",x"068d",x"3b06",x"39c3",x"b3a5",x"352b",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3d2",x"3530",x"3710",x"abf6",x"bbfc",x"0000",x"3b06",x"39c8"),
(x"b2d6",x"35c2",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41",x"b2d6",x"35c2",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2aa",x"35cd",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46"),
(x"b790",x"3548",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47",x"b790",x"3548",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b77b",x"3553",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c"),
(x"b73e",x"362d",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1",x"b73e",x"362d",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b705",x"3621",x"3710",x"34b8",x"3ba4",x"868d",x"3a87",x"3afc"),
(x"b368",x"3536",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd",x"b368",x"3536",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b3a5",x"352b",x"3710",x"32b5",x"bbd2",x"068d",x"3b06",x"39c3"),
(x"b2aa",x"35cd",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46",x"b2aa",x"35cd",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b261",x"35e2",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e"),
(x"b7a8",x"3544",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43",x"b7a8",x"3544",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b790",x"3548",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47"),
(x"b705",x"3621",x"3710",x"34b8",x"3ba4",x"868d",x"3a87",x"3afc",x"b705",x"3621",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b6f1",x"3610",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01"),
(x"b340",x"354d",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7",x"b340",x"354d",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b368",x"3536",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd"),
(x"b261",x"35e2",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e",x"b261",x"35e2",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b22d",x"35e9",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53"),
(x"b7bd",x"353c",x"3710",x"b821",x"3ad9",x"8000",x"3a95",x"3a3e",x"b7bd",x"353c",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7a8",x"3544",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43"),
(x"b6f1",x"3610",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01",x"b6f1",x"3610",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6ef",x"35fa",x"3710",x"3be9",x"b0b7",x"0000",x"3a87",x"3b05"),
(x"b33a",x"3562",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3",x"b33a",x"3562",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b340",x"354d",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7"),
(x"b22d",x"35e9",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53",x"b22d",x"35e9",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b1fd",x"35e3",x"3710",x"35da",x"3b72",x"0000",x"3a79",x"3b57"),
(x"b7c7",x"3533",x"3710",x"bb43",x"36b3",x"0000",x"3a95",x"3a3c",x"b7c7",x"3533",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7bd",x"353c",x"3710",x"b821",x"3ad9",x"8000",x"3a95",x"3a3e"),
(x"b6ef",x"35fa",x"3710",x"3be9",x"b0b7",x"0000",x"3a87",x"3b05",x"b6ef",x"35fa",x"36da",x"3b57",x"b658",x"068d",x"3a7d",x"3b05",x"b6fb",x"35eb",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08"),
(x"b351",x"3574",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af",x"b351",x"3574",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b33a",x"3562",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3"),
(x"b1fd",x"35e3",x"3710",x"35da",x"3b72",x"0000",x"3a79",x"3b57",x"b1fd",x"35e3",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1c1",x"35d1",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e"),
(x"b7c7",x"352e",x"3710",x"b744",x"bb20",x"8a8d",x"3a95",x"3a3b",x"b7c7",x"352e",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"3533",x"3710",x"bb43",x"36b3",x"0000",x"3a95",x"3a3c"),
(x"b6fb",x"35eb",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08",x"b6fb",x"35eb",x"36da",x"37ed",x"baf2",x"0000",x"3a7d",x"3b08",x"b721",x"35da",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10"),
(x"b34f",x"357c",x"3710",x"3448",x"bbb5",x"0000",x"3b06",x"39ae",x"b34f",x"357c",x"36da",x"3913",x"ba2f",x"0000",x"3afb",x"39ae",x"b351",x"3574",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af"),
(x"b1c1",x"35d1",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e",x"b1c1",x"35d1",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1a1",x"35cc",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61"),
(x"b7a4",x"351f",x"3710",x"b64b",x"bb5a",x"0000",x"3a95",x"3a34",x"b7a4",x"351f",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7c7",x"352e",x"3710",x"b744",x"bb20",x"8a8d",x"3a95",x"3a3b"),
(x"b721",x"35da",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10",x"b721",x"35da",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b72e",x"35d1",x"3710",x"39a7",x"b9a8",x"0000",x"3a87",x"3b13"),
(x"b326",x"357e",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae",x"b326",x"357e",x"36da",x"a5e3",x"bbff",x"0000",x"3a6e",x"3bae",x"b34f",x"357c",x"3710",x"3448",x"bbb5",x"0000",x"3a79",x"3bb2"),
(x"b1a1",x"35cc",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61",x"b1a1",x"35cc",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b161",x"35ca",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67"),
(x"b783",x"3511",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d",x"b783",x"3511",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b7a4",x"351f",x"3710",x"b64b",x"bb5a",x"0000",x"3a95",x"3a34"),
(x"b72e",x"35d1",x"3710",x"39a7",x"b9a8",x"0000",x"3aa1",x"39c6",x"b72e",x"35d1",x"36da",x"3b4f",x"b67e",x"0000",x"3a97",x"39c6",x"b72d",x"35c9",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8"),
(x"b2d6",x"3579",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6",x"b2d6",x"3579",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b326",x"357e",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae"),
(x"b161",x"35ca",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67",x"b161",x"35ca",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b135",x"35c1",x"3710",x"3822",x"3ad9",x"0000",x"3a79",x"3b6c"),
(x"b73e",x"350e",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20",x"b73e",x"350e",x"36da",x"27ae",x"bbfe",x"0000",x"3a8a",x"3a20",x"b783",x"3511",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d"),
(x"b72d",x"35c9",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8",x"b72d",x"35c9",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b721",x"35c6",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca"),
(x"b2aa",x"356e",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2",x"b2aa",x"356e",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2d6",x"3579",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6"),
(x"b135",x"35c1",x"3710",x"3822",x"3ad9",x"0000",x"3a79",x"3b6c",x"b135",x"35c1",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b116",x"35af",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70"),
(x"b705",x"351a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15",x"b705",x"351a",x"36da",x"34b8",x"bba4",x"0000",x"3a8a",x"3a15",x"b73e",x"350e",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20"),
(x"b575",x"3615",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28",x"b575",x"3615",x"36da",x"bab5",x"385c",x"0000",x"3a97",x"3a28",x"b568",x"3623",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b"),
(x"b938",x"3576",x"3710",x"bbc9",x"a82f",x"3347",x"3bf8",x"39db",x"b938",x"3576",x"36da",x"bbfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"b93a",x"35c9",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3be8",x"39da"),
(x"b261",x"3559",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a",x"b261",x"3559",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b2aa",x"356e",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2"),
(x"b931",x"3629",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63",x"b931",x"3629",x"36da",x"23ae",x"3bff",x"0000",x"3be3",x"3a63",x"b8ff",x"3627",x"3710",x"257a",x"3bff",x"15bc",x"3bd9",x"3a4f"),
(x"b6f1",x"352c",x"3710",x"3b73",x"b5d3",x"868d",x"3a95",x"3a10",x"b6f1",x"352c",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b705",x"351a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15"),
(x"b721",x"35c6",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca",x"b721",x"35c6",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b669",x"35c7",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed"),
(x"b22d",x"3552",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94",x"b22d",x"3552",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b261",x"3559",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a"),
(x"b6ef",x"3541",x"3710",x"3b57",x"3658",x"868d",x"3a95",x"3a0c",x"b6ef",x"3541",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6f1",x"352c",x"3710",x"3b73",x"b5d3",x"868d",x"3a95",x"3a10"),
(x"b669",x"35c7",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed",x"b669",x"35c7",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b63d",x"35cf",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5"),
(x"b930",x"356e",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c",x"b930",x"356e",x"36da",x"b67a",x"bb50",x"0000",x"3bc0",x"3984",x"b938",x"3576",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a"),
(x"b930",x"356e",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0",x"b92a",x"356e",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b92b",x"3513",x"3732",x"bb64",x"243f",x"361b",x"39f3",x"33aa"),
(x"b92a",x"356e",x"3733",x"bb1e",x"2518",x"3748",x"3a06",x"339f",x"b922",x"356e",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b924",x"3514",x"3749",x"ba3b",x"2680",x"3902",x"39f3",x"3392"),
(x"b922",x"356e",x"3748",x"b86c",x"29d9",x"3aa7",x"3a06",x"3388",x"b91b",x"356e",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b91f",x"3513",x"374e",x"ac96",x"29b2",x"3bf8",x"39f2",x"3387"),
(x"b91b",x"356e",x"3749",x"3594",x"2b76",x"3b7b",x"3a06",x"337b",x"b913",x"356e",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b918",x"3514",x"374b",x"38f0",x"29d6",x"3a48",x"39f2",x"337b"),
(x"b913",x"356e",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b913",x"3575",x"373a",x"3ae3",x"2b4b",x"380a",x"3bb9",x"399f",x"b90e",x"3574",x"370e",x"3754",x"3ae5",x"32eb",x"3bbd",x"39a7"),
(x"b913",x"3575",x"373a",x"3ae3",x"2b4b",x"380a",x"3bb9",x"399f",x"b913",x"356e",x"373b",x"381d",x"3a67",x"34eb",x"3bba",x"399e",x"b91b",x"356e",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b"),
(x"b913",x"3575",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1",x"b913",x"35c8",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b90f",x"35c9",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7"),
(x"b90f",x"35c9",x"3727",x"3bc1",x"a907",x"33bf",x"3be8",x"39f7",x"b90e",x"3574",x"370e",x"3bcb",x"a949",x"330f",x"3bf9",x"39fa",x"b913",x"3575",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1"),
(x"b913",x"35c8",x"373e",x"3a92",x"a9a8",x"388c",x"3be8",x"39f2",x"b913",x"3575",x"373a",x"3b64",x"a9cf",x"3612",x"3bf8",x"39f1",x"b91b",x"3577",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed"),
(x"b91a",x"35c8",x"374d",x"36b8",x"aa9e",x"3b3f",x"3be8",x"39ee",x"b91b",x"3577",x"374a",x"38ae",x"aa28",x"3a79",x"3bf7",x"39ed",x"b924",x"3577",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b928",x"35c8",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b922",x"35c8",x"3751",x"a11e",x"aa52",x"3bfd",x"3be8",x"39eb",x"b924",x"3577",x"374d",x"af62",x"aa90",x"3bef",x"3bf7",x"39ea"),
(x"b92f",x"35c8",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b928",x"35c8",x"374d",x"b867",x"a907",x"3aab",x"3be8",x"39e8",x"b92b",x"3577",x"3744",x"b96c",x"a921",x"39df",x"3bf7",x"39e6"),
(x"b935",x"35c8",x"3725",x"bb50",x"a638",x"3678",x"3be8",x"39de",x"b92f",x"35c8",x"373f",x"baad",x"a687",x"3865",x"3be8",x"39e4",x"b930",x"3577",x"3738",x"bb36",x"a61e",x"36e8",x"3bf7",x"39e3"),
(x"b930",x"3577",x"3738",x"b75b",x"bae5",x"32d3",x"3bb5",x"3992",x"b92a",x"356e",x"3733",x"b800",x"ba99",x"3437",x"3bb7",x"3993",x"b930",x"356e",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bba",x"398c"),
(x"b913",x"356e",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b90c",x"3513",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352",x"b912",x"3513",x"373c",x"3aea",x"2832",x"3802",x"39f2",x"336a"),
(x"b913",x"356e",x"373b",x"3aa1",x"2559",x"3879",x"3a05",x"3369",x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e",x"b90c",x"3513",x"3724",x"3af5",x"1a59",x"37e2",x"39f2",x"3352"),
(x"b91b",x"3577",x"374a",x"3544",x"b37d",x"3b51",x"3bb7",x"399b",x"b91b",x"356e",x"3749",x"382b",x"a432",x"3ad3",x"3bb8",x"399b",x"b922",x"356e",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998"),
(x"b922",x"356e",x"3748",x"b511",x"b92e",x"398b",x"3bb7",x"3998",x"b92a",x"356e",x"3733",x"b800",x"ba99",x"3437",x"3bb7",x"3993",x"b92b",x"3577",x"3744",x"b778",x"ba1b",x"3725",x"3bb4",x"3995"),
(x"b935",x"35c8",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b93a",x"35c9",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"3861",x"b931",x"35cd",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b92f",x"35c8",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b935",x"35c8",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3865",x"b92a",x"35ce",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"386b"),
(x"b928",x"35c8",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"386e",x"b92f",x"35c8",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"386a",x"b925",x"35ce",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"386e"),
(x"b91a",x"35c8",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b922",x"35c8",x"3751",x"9a8d",x"39ac",x"39a3",x"3b24",x"3871",x"b920",x"35ce",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"3871"),
(x"b913",x"35c8",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b91a",x"35c8",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3873",x"b919",x"35cf",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3873"),
(x"b90f",x"35c9",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3879",x"b913",x"35c8",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3876",x"b913",x"35cf",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3875"),
(x"b90d",x"35c9",x"3711",x"b36d",x"a40b",x"3bc7",x"3a19",x"3349",x"b906",x"35cc",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d",x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b92f",x"3629",x"372b",x"bbac",x"a891",x"347c",x"3a2d",x"33b1",x"b92a",x"35ce",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b931",x"35cd",x"3710",x"bbea",x"a7ae",x"307d",x"3a19",x"33c4"),
(x"b92a",x"35ce",x"3739",x"bb13",x"a8dd",x"3771",x"3a1a",x"339e",x"b92c",x"3629",x"373a",x"baa5",x"a5fd",x"3872",x"3a2d",x"33a3",x"b925",x"3628",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b920",x"35ce",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b925",x"35ce",x"3746",x"b918",x"a84d",x"3a28",x"3a1a",x"338e",x"b925",x"3628",x"3749",x"b926",x"a7c8",x"3a1d",x"3a2d",x"3391"),
(x"b919",x"35cf",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b920",x"35ce",x"374b",x"b451",x"a960",x"3bb2",x"3a1a",x"3385",x"b91f",x"3628",x"374f",x"a812",x"a959",x"3bfd",x"3a2d",x"3385"),
(x"b913",x"35cf",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b919",x"35cf",x"3749",x"3647",x"a97a",x"3b59",x"3a1a",x"3379",x"b918",x"3627",x"374b",x"38ec",x"a7f6",x"3a4c",x"3a2d",x"3378"),
(x"b913",x"35cf",x"373e",x"3ac8",x"a7bb",x"383c",x"3a1a",x"336a",x"b911",x"3628",x"373c",x"3ac9",x"a6b5",x"383a",x"3a2d",x"3366",x"b90b",x"3627",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c"),
(x"b90b",x"35ce",x"371c",x"3aa9",x"a818",x"386b",x"3a1a",x"334a",x"b90b",x"3627",x"3722",x"3b0f",x"a82c",x"3781",x"3a2d",x"334c",x"b907",x"3627",x"3718",x"38f7",x"a86d",x"3a44",x"3a2d",x"3340"),
(x"b116",x"35af",x"3710",x"8000",x"0000",x"3c00",x"3a13",x"2451",x"b116",x"358c",x"3710",x"8000",x"0000",x"3c00",x"3a0c",x"2451",x"b135",x"357a",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1"),
(x"b135",x"35c1",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"24c1",x"b135",x"357a",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"24c1",x"b161",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f"),
(x"b161",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"255f",x"b161",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"255f",x"b1a1",x"356f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643"),
(x"b1a1",x"356f",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2643",x"b1c1",x"356b",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"26b3",x"b1c1",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3"),
(x"b1c1",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"26b3",x"b1c1",x"356b",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"26b3",x"b1fd",x"3558",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b"),
(x"b1fd",x"3558",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"278b",x"b22d",x"3552",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"281a",x"b22d",x"35e9",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a"),
(x"b22d",x"35e9",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"281a",x"b22d",x"3552",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"281a",x"b261",x"3559",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878"),
(x"b261",x"35e2",x"3710",x"8000",x"0000",x"3c00",x"3a1e",x"2878",x"b261",x"3559",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2878",x"b2aa",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb"),
(x"b2aa",x"35cd",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"28fb",x"b2aa",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"28fb",x"b2d6",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949"),
(x"b2d6",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2949",x"b2d6",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2949",x"b326",x"357e",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7"),
(x"b326",x"35bd",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"29d7",x"b326",x"357e",x"3710",x"8000",x"0000",x"3c00",x"3a09",x"29d7",x"b34f",x"357c",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20"),
(x"b451",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b50c",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2d8d",x"b50c",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d"),
(x"b451",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2c3f",x"b451",x"35c5",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2c3f",x"b441",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23"),
(x"b441",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2c23",x"b441",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2c23",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b34f",x"35bf",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20"),
(x"b40b",x"3613",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b84",x"b3f4",x"3612",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b413",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2ba0"),
(x"b3f4",x"3612",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2b48",x"b3d2",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b409",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2b7d"),
(x"b3d2",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2b0a",x"b3a5",x"3610",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b407",x"35f1",x"3710",x"8000",x"0000",x"3c00",x"3a21",x"2b76"),
(x"b40b",x"3528",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b84",x"b413",x"352d",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2ba0",x"b413",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0"),
(x"b3f4",x"352a",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2b48",x"b413",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2ba0",x"b409",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d"),
(x"b3d2",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2b0a",x"b409",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2b7d",x"b407",x"354a",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76"),
(x"b3a5",x"352b",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"2aba",x"b407",x"354a",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2b76",x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b3a5",x"3610",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"2aba",x"b368",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b"),
(x"b50c",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2d8d",x"b50c",x"3576",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2d8d",x"b526",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb"),
(x"b62a",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b",x"b62a",x"35cd",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2f8b",x"b5ce",x"35c0",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7"),
(x"b5ce",x"35c0",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ee7",x"b5bd",x"35c3",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ec9",x"b5bd",x"3578",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9"),
(x"b5bd",x"3578",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"2ec9",x"b5bd",x"35c3",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"2ec9",x"b5a1",x"35d3",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97"),
(x"b5a1",x"3568",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2e97",x"b5a1",x"35d3",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2e97",x"b581",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e"),
(x"b581",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"2e5e",x"b568",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b568",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b50d",x"3638",x"3710",x"8000",x"0000",x"3c00",x"3a30",x"2d8e",x"b4f9",x"362f",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"2d6a",x"b4f5",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63"),
(x"b52b",x"3634",x"3710",x"8000",x"0000",x"3c00",x"3a2f",x"2dc4",x"b4f5",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"2d63",x"b4f2",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b4f5",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b4f9",x"350c",x"3710",x"8000",x"0000",x"3c00",x"39f0",x"2d6a",x"b50d",x"3503",x"3710",x"8000",x"0000",x"3c00",x"39ee",x"2d8e"),
(x"b4f2",x"3527",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e",x"b4f5",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2d63",x"b52b",x"3507",x"3710",x"8000",x"0000",x"3c00",x"39ef",x"2dc4"),
(x"b568",x"3518",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"2e32",x"b575",x"3526",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2e49",x"b575",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47"),
(x"b558",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2e14",x"b575",x"3530",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"2e47",x"b569",x"353b",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33"),
(x"b568",x"3623",x"3710",x"8000",x"0000",x"3c00",x"3a2c",x"2e32",x"b558",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b575",x"360b",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"2e47"),
(x"b558",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2e14",x"b544",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0",x"b569",x"3600",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33"),
(x"b4e1",x"35e6",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2d40",x"b51a",x"35db",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b4da",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"2d33"),
(x"b4e1",x"3555",x"3710",x"8000",x"0000",x"3c00",x"3a00",x"2d40",x"b4d8",x"354d",x"3710",x"8000",x"0000",x"3c00",x"39fe",x"2d2f",x"b4da",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33"),
(x"b51a",x"3560",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"2da6",x"b4da",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"2d33",x"b4f2",x"3527",x"3710",x"8000",x"0000",x"3c00",x"39f6",x"2d5e"),
(x"b51a",x"35db",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"2da6",x"b528",x"35d4",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b4f2",x"3615",x"3710",x"8000",x"0000",x"3c00",x"3a29",x"2d5e"),
(x"b528",x"35d4",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b569",x"3600",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"2e33",x"b544",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"2df0"),
(x"b544",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"2df0",x"b569",x"353b",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33",x"b528",x"3567",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf"),
(x"b528",x"35d4",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"2dbf",x"b52c",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5",x"b568",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30"),
(x"b528",x"3567",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"2dbf",x"b569",x"353b",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"2e33",x"b568",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"2e30"),
(x"b526",x"3571",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2dbb",x"b52c",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5",x"b52c",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5"),
(x"b568",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"2e30",x"b52c",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2dc5",x"b52c",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2dc5"),
(x"b63d",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b62a",x"35cd",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"2f8b",x"b62a",x"356e",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2f8b"),
(x"b669",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b63d",x"35cf",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"2fac",x"b63d",x"356c",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2fac"),
(x"b669",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2ffc",x"b669",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"2ffc",x"b721",x"3575",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b72d",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b721",x"35c6",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30a2",x"b721",x"3575",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"30a2"),
(x"b794",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b7c0",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130",x"b7c0",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130"),
(x"b794",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"3109",x"b794",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"3109",x"b77a",x"35d6",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1"),
(x"b77a",x"3565",x"3710",x"8000",x"0000",x"3c00",x"3a03",x"30f1",x"b77a",x"35d6",x"3710",x"8000",x"0000",x"3c00",x"3a1b",x"30f1",x"b776",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b776",x"355b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed",x"b776",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed",x"b72d",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad"),
(x"b6fb",x"3550",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b6ef",x"3541",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3075",x"b6f1",x"352c",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3076"),
(x"b721",x"3562",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b6fb",x"3550",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3080",x"b705",x"351a",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3088"),
(x"b6f1",x"3610",x"3710",x"8000",x"0000",x"3c00",x"3a28",x"3076",x"b6ef",x"35fa",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3075",x"b6fb",x"35eb",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080"),
(x"b705",x"3621",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3088",x"b6fb",x"35eb",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3080",x"b721",x"35da",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2"),
(x"b73e",x"362d",x"3710",x"8000",x"0000",x"3c00",x"3a2e",x"30bc",x"b721",x"35da",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"30a2",x"b72e",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae"),
(x"b72e",x"356a",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b721",x"3562",x"3710",x"8000",x"0000",x"3c00",x"3a02",x"30a2",x"b73e",x"350e",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30bc"),
(x"b7c7",x"352e",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"3135",x"b7c7",x"3533",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"3136",x"b7bd",x"353c",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d"),
(x"b7c7",x"360d",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3135",x"b7a4",x"361c",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b7bd",x"35ff",x"3710",x"8000",x"0000",x"3c00",x"3a24",x"312d"),
(x"b7a4",x"361c",x"3710",x"8000",x"0000",x"3c00",x"3a2a",x"3117",x"b783",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b7a8",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a"),
(x"b7a4",x"351f",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"3117",x"b7bd",x"353c",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"312d",x"b7a8",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a"),
(x"b72e",x"356a",x"3710",x"8000",x"0000",x"3c00",x"3a04",x"30ae",x"b77b",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b776",x"355b",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"30ed"),
(x"b72e",x"35d1",x"3710",x"8000",x"0000",x"3c00",x"3a1a",x"30ae",x"b72d",x"35c9",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"30ad",x"b776",x"35e0",x"3710",x"8000",x"0000",x"3c00",x"3a1d",x"30ed"),
(x"b77b",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"30f2",x"b783",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b790",x"3548",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3107"),
(x"b801",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b7c0",x"35c2",x"3710",x"8000",x"0000",x"3c00",x"3a17",x"3130",x"b7c0",x"3579",x"3710",x"8000",x"0000",x"3c00",x"3a07",x"3130"),
(x"b820",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b801",x"35ca",x"3710",x"8000",x"0000",x"3c00",x"3a19",x"316b",x"b801",x"3572",x"3710",x"8000",x"0000",x"3c00",x"3a06",x"316b"),
(x"b820",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"31a2",x"b820",x"3554",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"31a2",x"b83a",x"351e",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b84a",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b83a",x"361d",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"31d0",x"b83a",x"351e",x"3710",x"8000",x"0000",x"3c00",x"39f4",x"31d0"),
(x"b85e",x"3620",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b84a",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"31ed",x"b84a",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"31ed"),
(x"b865",x"360e",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b85e",x"3620",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3211",x"b85e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3211"),
(x"b867",x"3602",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b865",x"360e",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"321d",x"b865",x"352d",x"3710",x"8000",x"0000",x"3c00",x"39f7",x"321d"),
(x"b867",x"3602",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"3222",x"b867",x"3539",x"3710",x"8000",x"0000",x"3c00",x"39fa",x"3222",x"b86e",x"3541",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b87d",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b86e",x"35fa",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"322d",x"b86e",x"3541",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"322d"),
(x"b88f",x"360c",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b87d",x"35fb",x"3710",x"8000",x"0000",x"3c00",x"3a23",x"3248",x"b87d",x"3540",x"3710",x"8000",x"0000",x"3c00",x"39fb",x"3248"),
(x"b88f",x"360c",x"3710",x"8000",x"0000",x"3c00",x"3a27",x"3269",x"b88f",x"352f",x"3710",x"8000",x"0000",x"3c00",x"39f8",x"3269",x"b89e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b8a3",x"3622",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b89e",x"3620",x"3710",x"8000",x"0000",x"3c00",x"3a2b",x"3284",x"b89e",x"351b",x"3710",x"8000",x"0000",x"3c00",x"39f3",x"3284"),
(x"b8a3",x"3622",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b8a3",x"3519",x"3710",x"2081",x"9ea7",x"3bff",x"39f3",x"328d",x"b907",x"3571",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a06",x"333e"),
(x"b8ff",x"3627",x"3710",x"2904",x"26d5",x"3bfd",x"3a2d",x"3331",x"b8a3",x"3622",x"3710",x"2160",x"1cd0",x"3bff",x"3a2c",x"328d",x"b906",x"35cc",x"3713",x"29ab",x"208e",x"3bfd",x"3a19",x"333d"),
(x"b918",x"3627",x"374b",x"270a",x"3bfd",x"287a",x"3bce",x"3a59",x"b91f",x"3628",x"374f",x"28f4",x"3bfa",x"ac2a",x"3bcd",x"3a5c",x"b925",x"3628",x"3749",x"257a",x"3bfd",x"28f7",x"3bcf",x"3a5e"),
(x"b911",x"3628",x"373c",x"2504",x"3bff",x"2111",x"3bd1",x"3a56",x"b925",x"3628",x"3749",x"257a",x"3bfd",x"28f7",x"3bcf",x"3a5e",x"b92c",x"3629",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60"),
(x"b90b",x"3627",x"3722",x"2773",x"3bfe",x"22dc",x"3bd6",x"3a54",x"b92c",x"3629",x"373a",x"25e9",x"3bff",x"17c8",x"3bd1",x"3a60",x"b92f",x"3629",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62"),
(x"b907",x"3627",x"3718",x"25bc",x"3bfe",x"2673",x"3bd8",x"3a52",x"b92f",x"3629",x"372b",x"26c2",x"3bfe",x"24a2",x"3bd4",x"3a62",x"b931",x"3629",x"3710",x"2418",x"3bff",x"1a24",x"3bd9",x"3a63"),
(x"b924",x"3514",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b91f",x"3513",x"374e",x"281b",x"bbe6",x"b0f4",x"3a92",x"3a5c",x"b918",x"3514",x"374b",x"2511",x"bbff",x"2259",x"3a91",x"3a59"),
(x"b92b",x"3513",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b924",x"3514",x"3749",x"1ef6",x"bbff",x"23ef",x"3a90",x"3a5e",x"b912",x"3513",x"373c",x"184d",x"bbff",x"26c8",x"3a8e",x"3a57"),
(x"b931",x"3514",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63",x"b92b",x"3513",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a8c",x"3a60",x"b90c",x"3513",x"3724",x"9e3f",x"bbff",x"a018",x"3a89",x"3a55"),
(x"b1fd",x"3558",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b22d",x"3552",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b22d",x"3552",x"3710",x"2c28",x"bbfb",x"0000",x"3a79",x"3b94"),
(x"b6fb",x"3550",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6ef",x"3541",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6ef",x"3541",x"3710",x"3b57",x"3658",x"868d",x"3a95",x"3a0c"),
(x"b63d",x"35cf",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b62a",x"35cd",x"36da",x"303a",x"3bed",x"8000",x"3a97",x"39f9",x"b62a",x"35cd",x"3710",x"2fb9",x"3bf1",x"0000",x"3aa1",x"39f9"),
(x"b1c1",x"356b",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1fd",x"3558",x"36da",x"35da",x"bb72",x"0000",x"3a6e",x"3b90",x"b1fd",x"3558",x"3710",x"375d",x"bb1a",x"0000",x"3a79",x"3b90"),
(x"b906",x"3513",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b931",x"3514",x"36da",x"9e3f",x"bc00",x"0000",x"3a7b",x"3a63",x"b931",x"3514",x"3710",x"9edc",x"bc00",x"9dbc",x"3a85",x"3a63"),
(x"b721",x"3562",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b6fb",x"3550",x"36da",x"38e1",x"3a57",x"0000",x"3a8a",x"3a08",x"b6fb",x"3550",x"3710",x"37ed",x"3af2",x"0000",x"3a95",x"3a08"),
(x"b575",x"360b",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"3615",x"36da",x"bab5",x"385c",x"0000",x"3a97",x"3a28",x"b575",x"3615",x"3710",x"bb97",x"350d",x"0000",x"3aa1",x"3a28"),
(x"b1a1",x"356f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1c1",x"356b",x"36da",x"37bd",x"bb00",x"0000",x"3a6e",x"3b89",x"b1c1",x"356b",x"3710",x"3680",x"bb4f",x"0000",x"3a79",x"3b89"),
(x"b72e",x"356a",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b721",x"3562",x"36da",x"3711",x"3b2d",x"0000",x"3a8a",x"3a00",x"b721",x"3562",x"3710",x"37a6",x"3b06",x"0000",x"3a95",x"3a00"),
(x"b62a",x"35cd",x"36da",x"303a",x"3bed",x"8000",x"3a97",x"39f9",x"b5ce",x"35c0",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5ce",x"35c0",x"3710",x"2f27",x"3bf3",x"0000",x"3aa1",x"3a0b"),
(x"b161",x"3571",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b1a1",x"356f",x"36da",x"314e",x"bbe3",x"0000",x"3a6e",x"3b86",x"b1a1",x"356f",x"3710",x"2ede",x"bbf4",x"0000",x"3a79",x"3b86"),
(x"b72d",x"3572",x"36da",x"3a45",x"b8f8",x"0000",x"3a8a",x"39fb",x"b72e",x"356a",x"36da",x"39a7",x"39a8",x"0000",x"3a8a",x"39fd",x"b72e",x"356a",x"3710",x"3b4f",x"367e",x"0000",x"3a95",x"39fd"),
(x"b5ce",x"35c0",x"36da",x"2aec",x"3bfc",x"0000",x"3a97",x"3a0b",x"b5bd",x"35c3",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5bd",x"35c3",x"3710",x"b559",x"3b8a",x"0000",x"3aa1",x"3a0e"),
(x"b135",x"357a",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b161",x"3571",x"36da",x"30d8",x"bbe8",x"8000",x"3a6e",x"3b80",x"b161",x"3571",x"3710",x"3408",x"bbbd",x"0000",x"3a79",x"3b80"),
(x"b721",x"3575",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b72d",x"3572",x"36da",x"3a45",x"b8f8",x"0000",x"3a7c",x"3bb2",x"b72d",x"3572",x"3710",x"3778",x"bb13",x"0000",x"3a87",x"3bb2"),
(x"b5bd",x"35c3",x"36da",x"b6e1",x"3b38",x"0000",x"3a97",x"3a0e",x"b5a1",x"35d3",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b5a1",x"35d3",x"3710",x"b72d",x"3b26",x"0000",x"3aa1",x"3a14"),
(x"b93a",x"35c9",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"385a",x"b931",x"35cd",x"36da",x"b311",x"3bcd",x"0000",x"3b16",x"385d",x"b931",x"35cd",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3864"),
(x"b116",x"358c",x"36da",x"3b51",x"b675",x"8000",x"3a6e",x"3b77",x"b135",x"357a",x"36da",x"3822",x"bad9",x"8000",x"3a6e",x"3b7b",x"b135",x"357a",x"3710",x"3934",x"ba13",x"0000",x"3a79",x"3b7b"),
(x"b568",x"3518",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b575",x"3526",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3526",x"3710",x"bab5",x"b85c",x"0000",x"3a87",x"3b52"),
(x"b5a1",x"35d3",x"36da",x"b67b",x"3b50",x"0000",x"3a97",x"3a14",x"b581",x"35e0",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b581",x"35e0",x"3710",x"b794",x"3b0b",x"0000",x"3aa1",x"3a1a"),
(x"b669",x"3574",x"36da",x"a666",x"bbff",x"0000",x"3a7c",x"3b8d",x"b721",x"3575",x"36da",x"2560",x"bbff",x"0000",x"3a7c",x"3baf",x"b721",x"3575",x"3710",x"0cea",x"bc00",x"0000",x"3a87",x"3baf"),
(x"b581",x"35e0",x"36da",x"b89f",x"3a87",x"0000",x"3a97",x"3a1a",x"b568",x"35f7",x"36da",x"bb03",x"37b2",x"0000",x"3a97",x"3a21",x"b568",x"35f7",x"3710",x"b9f3",x"3958",x"0000",x"3aa1",x"3a21"),
(x"b8a3",x"3519",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b906",x"3513",x"36da",x"2273",x"bbff",x"0000",x"3a7b",x"3a53",x"b906",x"3513",x"3710",x"2546",x"bbff",x"9624",x"3a85",x"3a53"),
(x"b63d",x"356c",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b669",x"3574",x"36da",x"a666",x"bbff",x"0000",x"3a7c",x"3b8d",x"b669",x"3574",x"3710",x"abae",x"bbfc",x"8000",x"3a87",x"3b8d"),
(x"b568",x"3623",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b558",x"362a",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b558",x"362a",x"3710",x"b3cc",x"3bc2",x"8000",x"3aa1",x"3a2f"),
(x"b62a",x"356e",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b63d",x"356c",x"36da",x"affc",x"bbf0",x"8000",x"3a7c",x"3b84",x"b63d",x"356c",x"3710",x"ab45",x"bbfc",x"0000",x"3a87",x"3b84"),
(x"b558",x"362a",x"36da",x"b02d",x"3bee",x"0000",x"3a97",x"3a2f",x"b544",x"362a",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b544",x"362a",x"3710",x"b138",x"3be4",x"0000",x"3aa1",x"3a32"),
(x"b575",x"3526",x"36da",x"bb97",x"b50d",x"0000",x"3a7c",x"3b52",x"b575",x"3530",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b575",x"3530",x"3710",x"bb59",x"3650",x"0000",x"3a87",x"3b54"),
(x"b544",x"362a",x"36da",x"b46b",x"3bb0",x"0000",x"3a97",x"3a32",x"b52b",x"3634",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b52b",x"3634",x"3710",x"b472",x"3baf",x"0000",x"3aa1",x"3a37"),
(x"b5ce",x"357b",x"36da",x"2f27",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b62a",x"356e",x"36da",x"2fbb",x"bbf1",x"0000",x"3a7c",x"3b81",x"b62a",x"356e",x"3710",x"303a",x"bbed",x"0000",x"3a87",x"3b81"),
(x"b52b",x"3634",x"36da",x"b237",x"3bd8",x"8000",x"3a97",x"3a37",x"b50d",x"3638",x"36da",x"324b",x"3bd8",x"0000",x"3a97",x"3a3d",x"b50d",x"3638",x"3710",x"2546",x"3bff",x"068d",x"3aa1",x"3a3d"),
(x"b5bd",x"3578",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5ce",x"357b",x"36da",x"2f27",x"bbf3",x"0000",x"3a7c",x"3b6f",x"b5ce",x"357b",x"3710",x"2aec",x"bbfc",x"0000",x"3a87",x"3b6f"),
(x"b50d",x"3638",x"36da",x"324b",x"3bd8",x"0000",x"3a97",x"3a3d",x"b4f9",x"362f",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f9",x"362f",x"3710",x"38a5",x"3a82",x"0000",x"3aa1",x"3a41"),
(x"b5a1",x"3568",x"36da",x"b72d",x"bb26",x"0000",x"3a7c",x"3b66",x"b5bd",x"3578",x"36da",x"b559",x"bb8a",x"0000",x"3a7c",x"3b6c",x"b5bd",x"3578",x"3710",x"b6e1",x"bb38",x"0000",x"3a87",x"3b6c"),
(x"b4f9",x"362f",x"36da",x"3a57",x"38e0",x"8000",x"3a97",x"3a41",x"b4f5",x"3621",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f5",x"3621",x"3710",x"3bbb",x"341b",x"8000",x"3aa1",x"3a44"),
(x"b581",x"355c",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b5a1",x"3568",x"36da",x"b72d",x"bb26",x"0000",x"3a7c",x"3b66",x"b5a1",x"3568",x"3710",x"b67b",x"bb50",x"8000",x"3a87",x"3b66"),
(x"b4f5",x"3621",x"36da",x"3bc4",x"33a2",x"0000",x"3a97",x"3a44",x"b4f2",x"3615",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4f2",x"3615",x"3710",x"3aea",x"3805",x"0000",x"3aa1",x"3a47"),
(x"b931",x"35cd",x"36da",x"bbff",x"a4d0",x"0000",x"3a18",x"33f3",x"b931",x"3629",x"36da",x"bbff",x"a4d0",x"0000",x"3a2c",x"33f9",x"b931",x"3629",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a2c",x"33c9"),
(x"b8ff",x"3627",x"36da",x"26a7",x"3bff",x"8000",x"3be3",x"3a4f",x"b8a3",x"3622",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b8a3",x"3622",x"3710",x"286a",x"3bfe",x"868d",x"3bd9",x"3a2b"),
(x"b568",x"3544",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b581",x"355c",x"36da",x"b794",x"bb0b",x"0000",x"3a7c",x"3b5f",x"b581",x"355c",x"3710",x"b89f",x"ba87",x"0000",x"3a87",x"3b5f"),
(x"b4f2",x"3615",x"36da",x"3a46",x"38f6",x"0000",x"3a97",x"3a47",x"b4da",x"35fb",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4da",x"35fb",x"3710",x"3a4b",x"38ef",x"0000",x"3aa1",x"3a4d"),
(x"b8a3",x"3622",x"36da",x"2a59",x"3bfd",x"0000",x"3be3",x"3a2b",x"b89e",x"3620",x"36da",x"380f",x"3ae4",x"8000",x"3be3",x"3a29",x"b89e",x"3620",x"3710",x"36ef",x"3b35",x"0000",x"3bd9",x"3a29"),
(x"b558",x"3511",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b568",x"3518",x"36da",x"b919",x"ba29",x"8000",x"3a7c",x"3b4e",x"b568",x"3518",x"3710",x"b810",x"bae4",x"8000",x"3a87",x"3b4e"),
(x"b4da",x"35fb",x"36da",x"3afc",x"37cc",x"0000",x"3a97",x"3a4d",x"b4d8",x"35ef",x"36da",x"3af9",x"b7d7",x"8000",x"3a97",x"3a50",x"b4d8",x"35ef",x"3710",x"3be5",x"b11d",x"0000",x"3aa1",x"3a50"),
(x"b89e",x"3620",x"36da",x"380f",x"3ae4",x"8000",x"3be3",x"3a29",x"b88f",x"360c",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b88f",x"360c",x"3710",x"380a",x"3ae7",x"0000",x"3bd9",x"3a22"),
(x"b544",x"3511",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b558",x"3511",x"36da",x"b3cc",x"bbc2",x"8000",x"3a7c",x"3b4b",x"b558",x"3511",x"3710",x"b02d",x"bbee",x"0000",x"3a87",x"3b4b"),
(x"b4d8",x"35ef",x"36da",x"3af9",x"b7d7",x"8000",x"3a97",x"3a50",x"b4e1",x"35e6",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b4e1",x"35e6",x"3710",x"3599",x"bb7e",x"0000",x"3aa1",x"3a52"),
(x"b88f",x"360c",x"36da",x"377a",x"3b12",x"0000",x"3be3",x"3a22",x"b87d",x"35fb",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b87d",x"35fb",x"3710",x"3541",x"3b8e",x"0000",x"3bd9",x"3a1a"),
(x"b52b",x"3507",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b544",x"3511",x"36da",x"b138",x"bbe4",x"0000",x"3a7c",x"3b47",x"b544",x"3511",x"3710",x"b46b",x"bbb0",x"0000",x"3a87",x"3b47"),
(x"b4e1",x"35e6",x"36da",x"33d2",x"bbc1",x"868d",x"3a97",x"3a52",x"b51a",x"35db",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b51a",x"35db",x"3710",x"332b",x"bbcb",x"0000",x"3aa1",x"3a5d"),
(x"b87d",x"35fb",x"36da",x"3244",x"3bd8",x"0000",x"3be3",x"3a1a",x"b86e",x"35fa",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b86e",x"35fa",x"3710",x"ad01",x"3bf9",x"0000",x"3bd9",x"3a14"),
(x"b50d",x"3503",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b52b",x"3507",x"36da",x"b472",x"bbaf",x"8000",x"3a7c",x"3b42",x"b52b",x"3507",x"3710",x"b238",x"bbd8",x"0000",x"3a87",x"3b42"),
(x"b51a",x"35db",x"36da",x"347c",x"bbad",x"8000",x"3a97",x"3a5d",x"b528",x"35d4",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b528",x"35d4",x"3710",x"37fe",x"baed",x"0000",x"3aa1",x"3a60"),
(x"b86e",x"35fa",x"36da",x"b406",x"3bbe",x"8000",x"3be3",x"3a14",x"b867",x"3602",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b867",x"3602",x"3710",x"b975",x"39d9",x"0000",x"3bd9",x"3a11"),
(x"b4f9",x"350c",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b50d",x"3503",x"36da",x"253f",x"bbff",x"0000",x"3a7c",x"3b3c",x"b50d",x"3503",x"3710",x"324a",x"bbd8",x"0000",x"3a87",x"3b3c"),
(x"b528",x"35d4",x"36da",x"38ed",x"ba4d",x"0000",x"3a97",x"3a60",x"b52c",x"35cf",x"36da",x"3b0d",x"378c",x"0000",x"3a97",x"3a61",x"b52c",x"35cf",x"3710",x"3bfc",x"ab6c",x"0000",x"3aa1",x"3a61"),
(x"b867",x"3602",x"36da",x"baa2",x"3877",x"0000",x"3be3",x"3a11",x"b865",x"360e",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b865",x"360e",x"3710",x"bb0e",x"378a",x"8000",x"3bd9",x"3a0e"),
(x"b4f5",x"351a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f9",x"350c",x"36da",x"38a5",x"ba82",x"868d",x"3a7c",x"3b38",x"b4f9",x"350c",x"3710",x"3a57",x"b8e0",x"0000",x"3a87",x"3b38"),
(x"b52c",x"35cf",x"36da",x"3b0d",x"378c",x"0000",x"3a54",x"39ec",x"b526",x"35ca",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b526",x"35ca",x"3710",x"35f8",x"3b6b",x"0000",x"3a5f",x"39ee"),
(x"b865",x"360e",x"36da",x"baaf",x"3865",x"8000",x"3be3",x"3a0e",x"b85e",x"3620",x"36da",x"b5f3",x"3b6d",x"0a8d",x"3be3",x"3a09",x"b85e",x"3620",x"3710",x"b878",x"3aa2",x"0000",x"3bd9",x"3a09"),
(x"b4f2",x"3527",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f5",x"351a",x"36da",x"3bbb",x"b41b",x"0000",x"3a7c",x"3b35",x"b4f5",x"351a",x"3710",x"3bc4",x"b3a2",x"8000",x"3a87",x"3b35"),
(x"b526",x"35ca",x"36da",x"33bc",x"3bc3",x"0000",x"3a54",x"39ee",x"b50c",x"35c6",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b50c",x"35c6",x"3710",x"292b",x"3bfe",x"8000",x"3a5f",x"39f3"),
(x"b116",x"35af",x"36da",x"3bdf",x"31b0",x"8000",x"3a6e",x"3b70",x"b116",x"358c",x"36da",x"3b51",x"b675",x"8000",x"3a6e",x"3b77",x"b116",x"358c",x"3710",x"3bdf",x"b1b0",x"0000",x"3a79",x"3b77"),
(x"b85e",x"3620",x"36da",x"b5f3",x"3b6d",x"0a8d",x"3be3",x"3a09",x"b84a",x"362a",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b84a",x"362a",x"3710",x"ac15",x"3bfb",x"0000",x"3bd9",x"3a01"),
(x"b4da",x"3540",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4f2",x"3527",x"36da",x"3aea",x"b805",x"0000",x"3a7c",x"3b33",x"b4f2",x"3527",x"3710",x"3a46",x"b8f6",x"0000",x"3a87",x"3b33"),
(x"b451",x"35c5",x"36da",x"a987",x"3bfe",x"068d",x"3a54",x"3a16",x"b441",x"35ca",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b441",x"35ca",x"3710",x"b6f3",x"3b34",x"0000",x"3a5f",x"3a19"),
(x"b89e",x"351b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b8a3",x"3519",x"36da",x"284d",x"bbfe",x"8000",x"3a7b",x"3a2d",x"b8a3",x"3519",x"3710",x"2a1e",x"bbfd",x"0000",x"3a85",x"3a2d"),
(x"b84a",x"362a",x"36da",x"30e0",x"3be8",x"0000",x"3be3",x"3a01",x"b83a",x"361d",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b83a",x"361d",x"3710",x"3890",x"3a92",x"0000",x"3bd9",x"39fa"),
(x"b4d8",x"354d",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4da",x"3540",x"36da",x"3a4b",x"b8ef",x"068d",x"3a7c",x"3b2c",x"b4da",x"3540",x"3710",x"3afc",x"b7cc",x"0000",x"3a87",x"3b2c"),
(x"b50c",x"35c6",x"36da",x"236c",x"3bff",x"0000",x"3a54",x"39f3",x"b451",x"35c5",x"36da",x"a987",x"3bfe",x"068d",x"3a54",x"3a16",x"b451",x"35c5",x"3710",x"a0dd",x"3c00",x"0000",x"3a5f",x"3a16"),
(x"b88f",x"352f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b89e",x"351b",x"36da",x"36f0",x"bb35",x"0000",x"3a7b",x"3a2b",x"b89e",x"351b",x"3710",x"380f",x"bae4",x"0000",x"3a85",x"3a2b"),
(x"b568",x"35f7",x"36da",x"bb03",x"37b2",x"0000",x"3a97",x"3a21",x"b569",x"3600",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b569",x"3600",x"3710",x"bb2d",x"b70f",x"0000",x"3aa1",x"3a23"),
(x"b4e1",x"3555",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4d8",x"354d",x"36da",x"3be5",x"311d",x"8000",x"3a7c",x"3b2a",x"b4d8",x"354d",x"3710",x"3af9",x"37d8",x"8000",x"3a87",x"3b2a"),
(x"b441",x"35ca",x"36da",x"b7a3",x"3b07",x"0000",x"3a54",x"3a19",x"b40d",x"35e8",x"36da",x"b8bf",x"3a70",x"868d",x"3a54",x"3a25",x"b40d",x"35e8",x"3710",x"b83a",x"3aca",x"0000",x"3a5f",x"3a25"),
(x"b87d",x"3540",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b88f",x"352f",x"36da",x"380a",x"bae7",x"0000",x"3a7b",x"3a25",x"b88f",x"352f",x"3710",x"377a",x"bb12",x"0000",x"3a85",x"3a25"),
(x"b83a",x"361d",x"36da",x"3953",x"39f7",x"8000",x"3be3",x"39fa",x"b820",x"35e8",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b820",x"35e8",x"3710",x"391f",x"3a25",x"0000",x"3bd9",x"39ec"),
(x"b51a",x"3560",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b4e1",x"3555",x"36da",x"3599",x"3b7e",x"0000",x"3a7c",x"3b28",x"b4e1",x"3555",x"3710",x"33d2",x"3bc1",x"868d",x"3a87",x"3b28"),
(x"b40d",x"35e8",x"36da",x"b8bf",x"3a70",x"868d",x"3a54",x"3a25",x"b407",x"35f1",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b407",x"35f1",x"3710",x"bb61",x"3629",x"0000",x"3a5f",x"3a27"),
(x"b86e",x"3541",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b87d",x"3540",x"36da",x"3541",x"bb8e",x"0000",x"3a7b",x"3a1d",x"b87d",x"3540",x"3710",x"3244",x"bbd8",x"0000",x"3a85",x"3a1d"),
(x"b569",x"3600",x"36da",x"ba4b",x"b8f0",x"0000",x"3a97",x"3a23",x"b575",x"360b",x"36da",x"bb59",x"b650",x"8000",x"3a97",x"3a26",x"b575",x"360b",x"3710",x"ba67",x"b8cb",x"868d",x"3aa1",x"3a26"),
(x"b528",x"3567",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b51a",x"3560",x"36da",x"332b",x"3bcb",x"0000",x"3a7c",x"3b1d",x"b51a",x"3560",x"3710",x"347c",x"3bad",x"0000",x"3a87",x"3b1d"),
(x"b407",x"35f1",x"36da",x"bbf7",x"2ddb",x"0000",x"3a54",x"3a27",x"b409",x"35f7",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b409",x"35f7",x"3710",x"bb1a",x"b75d",x"8000",x"3a5f",x"3a28"),
(x"b867",x"3539",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b86e",x"3541",x"36da",x"ad01",x"bbf9",x"0000",x"3a7b",x"3a17",x"b86e",x"3541",x"3710",x"b406",x"bbbe",x"0000",x"3a85",x"3a17"),
(x"b820",x"35e8",x"36da",x"385c",x"3ab4",x"0000",x"3be3",x"39ec",x"b801",x"35ca",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b801",x"35ca",x"3710",x"3561",x"3b88",x"0000",x"3bd9",x"39de"),
(x"b52c",x"356c",x"36da",x"3bfc",x"2b6c",x"0000",x"3a7c",x"3b19",x"b528",x"3567",x"36da",x"37fe",x"3aed",x"0000",x"3a7c",x"3b1a",x"b528",x"3567",x"3710",x"38ed",x"3a4d",x"0000",x"3a87",x"3b1a"),
(x"b409",x"35f7",x"36da",x"bab5",x"b85b",x"0000",x"3a54",x"3a28",x"b413",x"3605",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"3605",x"3710",x"bb08",x"b7a1",x"0000",x"3a5f",x"3a2b"),
(x"b865",x"352d",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b867",x"3539",x"36da",x"b975",x"b9d8",x"0000",x"3a7b",x"3a14",x"b867",x"3539",x"3710",x"baa2",x"b877",x"0000",x"3a85",x"3a14"),
(x"b801",x"35ca",x"36da",x"3346",x"3bca",x"0000",x"3be3",x"39de",x"b7c0",x"35c2",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b7c0",x"35c2",x"3710",x"29e3",x"3bfd",x"0000",x"3bd9",x"39d1"),
(x"b526",x"3571",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b52c",x"356c",x"36da",x"3bfc",x"2b6c",x"0000",x"3afb",x"3a11",x"b52c",x"356c",x"3710",x"3b0d",x"b78c",x"0000",x"3b06",x"3a11"),
(x"b413",x"3605",x"36da",x"bba9",x"b498",x"8000",x"3a54",x"3a2b",x"b413",x"360e",x"36da",x"ba12",x"3935",x"068d",x"3a54",x"3a2d",x"b413",x"360e",x"3710",x"bb8c",x"354a",x"0000",x"3a5f",x"3a2d"),
(x"b85e",x"351b",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b865",x"352d",x"36da",x"bb0e",x"b78a",x"0000",x"3a7b",x"3a12",x"b865",x"352d",x"3710",x"baaf",x"b865",x"8000",x"3a85",x"3a12"),
(x"b7c0",x"35c2",x"36da",x"a984",x"3bfe",x"0000",x"3be3",x"39d1",x"b794",x"35c9",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b794",x"35c9",x"3710",x"b357",x"3bc9",x"0000",x"3bd9",x"39c8"),
(x"b50c",x"3576",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b526",x"3571",x"36da",x"35f8",x"bb6b",x"8000",x"3afb",x"3a0f",x"b526",x"3571",x"3710",x"33bb",x"bbc3",x"0000",x"3b06",x"3a0f"),
(x"b413",x"360e",x"36da",x"ba12",x"3935",x"068d",x"3a54",x"3a2d",x"b40b",x"3613",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b40b",x"3613",x"3710",x"b3aa",x"3bc4",x"8000",x"3a5f",x"3a2e"),
(x"b84a",x"3511",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b85e",x"351b",x"36da",x"b878",x"baa2",x"8000",x"3a7b",x"3a0d",x"b85e",x"351b",x"3710",x"b5f3",x"bb6d",x"0000",x"3a85",x"3a0d"),
(x"b794",x"35c9",x"36da",x"b51c",x"3b94",x"0000",x"3be3",x"39c8",x"b77a",x"35d6",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b77a",x"35d6",x"3710",x"b83f",x"3ac7",x"0000",x"3bd9",x"39c2"),
(x"b441",x"3571",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b451",x"3576",x"36da",x"a0ea",x"bc00",x"0000",x"3afb",x"39e7",x"b451",x"3576",x"3710",x"a987",x"bbfe",x"0000",x"3b06",x"39e7"),
(x"b40b",x"3613",x"36da",x"aabe",x"3bfd",x"8000",x"3a54",x"3a2e",x"b3f4",x"3612",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3f4",x"3612",x"3710",x"3148",x"3be3",x"8000",x"3a5f",x"3a32"),
(x"b83a",x"351e",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b84a",x"3511",x"36da",x"ac15",x"bbfb",x"8000",x"3a7b",x"3a05",x"b84a",x"3511",x"3710",x"30e0",x"bbe8",x"8000",x"3a85",x"3a05"),
(x"b77a",x"35d6",x"36da",x"b97c",x"39d2",x"8000",x"3be3",x"39c2",x"b776",x"35e0",x"36da",x"bbce",x"b2fb",x"0000",x"3be3",x"39c0",x"b776",x"35e0",x"3710",x"bbee",x"3038",x"0000",x"3bd9",x"39c0"),
(x"b451",x"3576",x"36da",x"a0ea",x"bc00",x"0000",x"3afb",x"39e7",x"b50c",x"3576",x"36da",x"292b",x"bbfe",x"8000",x"3afb",x"3a0a",x"b50c",x"3576",x"3710",x"236c",x"bbff",x"0000",x"3b06",x"3a0a"),
(x"b3f4",x"3612",x"36da",x"3408",x"3bbd",x"8000",x"3a54",x"3a32",x"b3d2",x"360b",x"36da",x"abf6",x"3bfc",x"0000",x"3a54",x"3a35",x"b3d2",x"360b",x"3710",x"2ffb",x"3bf0",x"0000",x"3a5f",x"3a35"),
(x"b569",x"353b",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b568",x"3544",x"36da",x"b9f3",x"b958",x"0000",x"3a7c",x"3b59",x"b568",x"3544",x"3710",x"bb03",x"b7b2",x"0000",x"3a87",x"3b59"),
(x"b776",x"35e0",x"36da",x"bbce",x"b2fb",x"0000",x"3be3",x"39c0",x"b77b",x"35e8",x"36da",x"b853",x"baba",x"0000",x"3be3",x"39be",x"b77b",x"35e8",x"3710",x"b937",x"ba10",x"0000",x"3bd9",x"39be"),
(x"b40d",x"3553",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b441",x"3571",x"36da",x"b6f3",x"bb34",x"8000",x"3afb",x"39e4",x"b441",x"3571",x"3710",x"b7a4",x"bb07",x"0000",x"3b06",x"39e4"),
(x"b3d2",x"360b",x"36da",x"abf6",x"3bfc",x"0000",x"3a54",x"3a35",x"b3a5",x"3610",x"36da",x"32b5",x"3bd2",x"8000",x"3a54",x"3a39",x"b3a5",x"3610",x"3710",x"24fd",x"3bff",x"0000",x"3a5f",x"3a39"),
(x"b820",x"3554",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b83a",x"351e",x"36da",x"3890",x"ba92",x"0000",x"3a7b",x"39ff",x"b83a",x"351e",x"3710",x"3953",x"b9f7",x"868d",x"3a85",x"39ff"),
(x"b77b",x"35e8",x"36da",x"b853",x"baba",x"0000",x"3a7d",x"3ac5",x"b790",x"35f3",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b790",x"35f3",x"3710",x"b606",x"bb69",x"0000",x"3a87",x"3ac9"),
(x"b407",x"354a",x"36da",x"bb61",x"b629",x"0000",x"3afb",x"39d6",x"b40d",x"3553",x"36da",x"b83a",x"baca",x"0000",x"3afb",x"39d8",x"b40d",x"3553",x"3710",x"b8bf",x"ba70",x"8000",x"3b06",x"39d8"),
(x"b3a5",x"3610",x"36da",x"32b5",x"3bd2",x"8000",x"3a54",x"3a39",x"b368",x"3605",x"36da",x"3912",x"3a2f",x"8000",x"3a54",x"3a40",x"b368",x"3605",x"3710",x"37ea",x"3af3",x"0000",x"3a5f",x"3a40"),
(x"b575",x"3530",x"36da",x"ba67",x"38cb",x"068d",x"3a7c",x"3b54",x"b569",x"353b",x"36da",x"bb2d",x"370f",x"0000",x"3a7c",x"3b57",x"b569",x"353b",x"3710",x"ba4b",x"38f0",x"0000",x"3a87",x"3b57"),
(x"b790",x"35f3",x"36da",x"b461",x"bbb1",x"0000",x"3a7d",x"3ac9",x"b7a8",x"35f7",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7a8",x"35f7",x"3710",x"b360",x"bbc8",x"0000",x"3a87",x"3ace"),
(x"b409",x"3544",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b407",x"354a",x"36da",x"bb61",x"b629",x"0000",x"3afb",x"39d6",x"b407",x"354a",x"3710",x"bbf7",x"addb",x"0000",x"3b06",x"39d6"),
(x"b368",x"3605",x"36da",x"3912",x"3a2f",x"8000",x"3a54",x"3a40",x"b340",x"35ee",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b340",x"35ee",x"3710",x"3aba",x"3853",x"0000",x"3a5f",x"3a45"),
(x"b801",x"3572",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b820",x"3554",x"36da",x"391f",x"ba25",x"0000",x"3a7b",x"39f1",x"b820",x"3554",x"3710",x"385c",x"bab4",x"0000",x"3a85",x"39f1"),
(x"b7a8",x"35f7",x"36da",x"b4b8",x"bba4",x"8000",x"3a7d",x"3ace",x"b7bd",x"35ff",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7bd",x"35ff",x"3710",x"b6d2",x"bb3c",x"0000",x"3a87",x"3ad2"),
(x"b413",x"3536",x"36da",x"bb08",x"37a1",x"868d",x"3afb",x"39d2",x"b409",x"3544",x"36da",x"bb1a",x"375c",x"8000",x"3afb",x"39d5",x"b409",x"3544",x"3710",x"bab5",x"385b",x"0000",x"3b06",x"39d5"),
(x"b340",x"35ee",x"36da",x"3b6b",x"35fb",x"0000",x"3a54",x"3a45",x"b33a",x"35d9",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b33a",x"35d9",x"3710",x"3bf6",x"ae02",x"0000",x"3a5f",x"3a49"),
(x"b7c0",x"3579",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b801",x"3572",x"36da",x"3561",x"bb88",x"0000",x"3a7b",x"39e4",x"b801",x"3572",x"3710",x"3346",x"bbca",x"0000",x"3a85",x"39e4"),
(x"b7bd",x"35ff",x"36da",x"b821",x"bada",x"8000",x"3a7d",x"3ad2",x"b7c7",x"3608",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"3608",x"3710",x"ba01",x"b948",x"8000",x"3a87",x"3ad5"),
(x"b931",x"3514",x"36da",x"bbff",x"26b5",x"0000",x"39f5",x"33fa",x"b930",x"356e",x"36da",x"bbff",x"26b5",x"0000",x"3a09",x"33f0",x"b930",x"356e",x"3710",x"bbeb",x"2604",x"3075",x"3a07",x"33c0"),
(x"b413",x"352d",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"3536",x"36da",x"bb08",x"37a1",x"868d",x"3afb",x"39d2",x"b413",x"3536",x"3710",x"bba9",x"3499",x"8000",x"3b06",x"39d2"),
(x"b33a",x"35d9",x"36da",x"3b88",x"b564",x"8000",x"3a54",x"3a49",x"b351",x"35c7",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b351",x"35c7",x"3710",x"3b23",x"b738",x"0000",x"3a5f",x"3a4d"),
(x"b794",x"3572",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b7c0",x"3579",x"36da",x"29e3",x"bbfd",x"0000",x"3a7b",x"39d7",x"b7c0",x"3579",x"3710",x"a984",x"bbfe",x"0000",x"3a85",x"39d7"),
(x"b7c7",x"3608",x"36da",x"bb43",x"b6b4",x"0000",x"3a7d",x"3ad5",x"b7c7",x"360d",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7c7",x"360d",x"3710",x"b8b7",x"3a76",x"0000",x"3a87",x"3ad6"),
(x"b40b",x"3528",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b413",x"352d",x"36da",x"bb8c",x"b54a",x"868d",x"3afb",x"39d0",x"b413",x"352d",x"3710",x"ba12",x"b935",x"868d",x"3b06",x"39d0"),
(x"b351",x"35c7",x"36da",x"3bb2",x"b458",x"0000",x"3a54",x"3a4d",x"b34f",x"35bf",x"36da",x"3448",x"3bb5",x"0000",x"3a54",x"3a4f",x"b34f",x"35bf",x"3710",x"3913",x"3a2f",x"0000",x"3a5f",x"3a4f"),
(x"b77a",x"3565",x"36da",x"b83f",x"bac7",x"0000",x"3a7b",x"39c9",x"b794",x"3572",x"36da",x"b358",x"bbc9",x"0000",x"3a7b",x"39cf",x"b794",x"3572",x"3710",x"b51c",x"bb94",x"0000",x"3a85",x"39cf"),
(x"b7c7",x"360d",x"36da",x"b744",x"3b20",x"8a8d",x"3a7d",x"3ad6",x"b7a4",x"361c",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b7a4",x"361c",x"3710",x"b655",x"3b58",x"8000",x"3a87",x"3add"),
(x"b3f4",x"352a",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b40b",x"3528",x"36da",x"b3aa",x"bbc4",x"8000",x"3afb",x"39ce",x"b40b",x"3528",x"3710",x"aabe",x"bbfd",x"0000",x"3b06",x"39ce"),
(x"b34f",x"35bf",x"36da",x"3448",x"3bb5",x"0000",x"3a6e",x"3b35",x"b326",x"35bd",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b326",x"35bd",x"3710",x"a5e3",x"3bff",x"0000",x"3a79",x"3b39"),
(x"b776",x"355b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b77a",x"3565",x"36da",x"b83f",x"bac7",x"0000",x"3a8a",x"3a50",x"b77a",x"3565",x"3710",x"b97c",x"b9d2",x"0000",x"3a95",x"3a50"),
(x"b7a4",x"361c",x"36da",x"b64a",x"3b5a",x"8000",x"3a7d",x"3add",x"b783",x"362a",x"36da",x"afa0",x"3bf1",x"068d",x"3a7d",x"3ae4",x"b783",x"362a",x"3710",x"b33d",x"3bca",x"0000",x"3a87",x"3ae4"),
(x"b3d2",x"3530",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3f4",x"352a",x"36da",x"3148",x"bbe3",x"8000",x"3afb",x"39cb",x"b3f4",x"352a",x"3710",x"3408",x"bbbd",x"0000",x"3b06",x"39cb"),
(x"b326",x"35bd",x"36da",x"ad8e",x"3bf8",x"0000",x"3a6e",x"3b39",x"b2d6",x"35c2",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2d6",x"35c2",x"3710",x"b287",x"3bd4",x"0000",x"3a79",x"3b41"),
(x"b77b",x"3553",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b776",x"355b",x"36da",x"bbee",x"b037",x"0000",x"3a8a",x"3a4d",x"b776",x"355b",x"3710",x"bbce",x"32fc",x"0000",x"3a95",x"3a4d"),
(x"b783",x"362a",x"36da",x"afa0",x"3bf1",x"068d",x"3a7d",x"3ae4",x"b73e",x"362d",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b73e",x"362d",x"3710",x"27ae",x"3bfe",x"0000",x"3a87",x"3af1"),
(x"b3a5",x"352b",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3d2",x"3530",x"36da",x"2ffb",x"bbf0",x"0000",x"3afb",x"39c8",x"b3d2",x"3530",x"3710",x"abf6",x"bbfc",x"0000",x"3b06",x"39c8"),
(x"b2d6",x"35c2",x"36da",x"b4dc",x"3b9f",x"0000",x"3a6e",x"3b41",x"b2aa",x"35cd",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b2aa",x"35cd",x"3710",x"b78b",x"3b0e",x"0000",x"3a79",x"3b46"),
(x"b790",x"3548",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b77b",x"3553",x"36da",x"b937",x"3a10",x"8000",x"3a8a",x"3a4c",x"b77b",x"3553",x"3710",x"b853",x"3aba",x"0000",x"3a95",x"3a4c"),
(x"b73e",x"362d",x"36da",x"2f57",x"3bf2",x"8000",x"3a7d",x"3af1",x"b705",x"3621",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b705",x"3621",x"3710",x"34b8",x"3ba4",x"868d",x"3a87",x"3afc"),
(x"b368",x"3536",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b3a5",x"352b",x"36da",x"2504",x"bbff",x"0000",x"3afb",x"39c3",x"b3a5",x"352b",x"3710",x"32b5",x"bbd2",x"068d",x"3b06",x"39c3"),
(x"b2aa",x"35cd",x"36da",x"b7e2",x"3af5",x"0000",x"3a6e",x"3b46",x"b261",x"35e2",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b261",x"35e2",x"3710",x"b72e",x"3b26",x"0000",x"3a79",x"3b4e"),
(x"b7a8",x"3544",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b790",x"3548",x"36da",x"b606",x"3b69",x"0000",x"3a8a",x"3a47",x"b790",x"3548",x"3710",x"b461",x"3bb1",x"0000",x"3a95",x"3a47"),
(x"b705",x"3621",x"36da",x"36ee",x"3b35",x"0000",x"3a7d",x"3afc",x"b6f1",x"3610",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6f1",x"3610",x"3710",x"3a69",x"38c9",x"0000",x"3a87",x"3b01"),
(x"b340",x"354d",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b368",x"3536",x"36da",x"37ea",x"baf3",x"8000",x"3afb",x"39bd",x"b368",x"3536",x"3710",x"3912",x"ba2f",x"8000",x"3b06",x"39bd"),
(x"b261",x"35e2",x"36da",x"b5e0",x"3b70",x"8000",x"3a6e",x"3b4e",x"b22d",x"35e9",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b22d",x"35e9",x"3710",x"ae88",x"3bf5",x"8000",x"3a79",x"3b53"),
(x"b7bd",x"353c",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7a8",x"3544",x"36da",x"b360",x"3bc8",x"8000",x"3a8a",x"3a43",x"b7a8",x"3544",x"3710",x"b4b8",x"3ba4",x"0000",x"3a95",x"3a43"),
(x"b6f1",x"3610",x"36da",x"3b73",x"35d3",x"8000",x"3a7d",x"3b01",x"b6ef",x"35fa",x"36da",x"3b57",x"b658",x"068d",x"3a7d",x"3b05",x"b6ef",x"35fa",x"3710",x"3be9",x"b0b7",x"0000",x"3a87",x"3b05"),
(x"b33a",x"3562",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b340",x"354d",x"36da",x"3aba",x"b853",x"0000",x"3afb",x"39b7",x"b340",x"354d",x"3710",x"3b6b",x"b5fb",x"8000",x"3b06",x"39b7"),
(x"b22d",x"35e9",x"36da",x"2c28",x"3bfb",x"8000",x"3a6e",x"3b53",x"b1fd",x"35e3",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1fd",x"35e3",x"3710",x"35da",x"3b72",x"0000",x"3a79",x"3b57"),
(x"b7c7",x"3533",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7bd",x"353c",x"36da",x"b6d2",x"3b3c",x"8000",x"3a8a",x"3a3e",x"b7bd",x"353c",x"3710",x"b821",x"3ad9",x"8000",x"3a95",x"3a3e"),
(x"b6ef",x"35fa",x"36da",x"3b57",x"b658",x"068d",x"3a7d",x"3b05",x"b6fb",x"35eb",x"36da",x"37ed",x"baf2",x"0000",x"3a7d",x"3b08",x"b6fb",x"35eb",x"3710",x"38e1",x"ba57",x"0000",x"3a87",x"3b08"),
(x"b351",x"3574",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b33a",x"3562",x"36da",x"3bf6",x"2e02",x"8000",x"3afb",x"39b3",x"b33a",x"3562",x"3710",x"3b88",x"3564",x"068d",x"3b06",x"39b3"),
(x"b1fd",x"35e3",x"36da",x"375d",x"3b1a",x"8000",x"3a6e",x"3b57",x"b1c1",x"35d1",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1c1",x"35d1",x"3710",x"37bd",x"3b00",x"0000",x"3a79",x"3b5e"),
(x"b7c7",x"352e",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"3533",x"36da",x"ba01",x"3948",x"0000",x"3a8a",x"3a3c",x"b7c7",x"3533",x"3710",x"bb43",x"36b3",x"0000",x"3a95",x"3a3c"),
(x"b6fb",x"35eb",x"36da",x"37ed",x"baf2",x"0000",x"3a7d",x"3b08",x"b721",x"35da",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b721",x"35da",x"3710",x"3711",x"bb2d",x"0000",x"3a87",x"3b10"),
(x"b34f",x"357c",x"36da",x"3913",x"ba2f",x"0000",x"3afb",x"39ae",x"b351",x"3574",x"36da",x"3b23",x"3738",x"0000",x"3afb",x"39af",x"b351",x"3574",x"3710",x"3bb2",x"3458",x"0000",x"3b06",x"39af"),
(x"b1c1",x"35d1",x"36da",x"3680",x"3b4f",x"8000",x"3a6e",x"3b5e",x"b1a1",x"35cc",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b1a1",x"35cc",x"3710",x"314e",x"3be3",x"0000",x"3a79",x"3b61"),
(x"b7a4",x"351f",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7c7",x"352e",x"36da",x"b8b7",x"ba76",x"0000",x"3a8a",x"3a3b",x"b7c7",x"352e",x"3710",x"b744",x"bb20",x"8a8d",x"3a95",x"3a3b"),
(x"b721",x"35da",x"36da",x"37a6",x"bb06",x"0000",x"3a7d",x"3b10",x"b72e",x"35d1",x"36da",x"3b4f",x"b67e",x"0000",x"3a7d",x"3b13",x"b72e",x"35d1",x"3710",x"39a7",x"b9a8",x"0000",x"3a87",x"3b13"),
(x"b326",x"357e",x"36da",x"a5e3",x"bbff",x"0000",x"3a6e",x"3bae",x"b34f",x"357c",x"36da",x"3913",x"ba2f",x"0000",x"3a6e",x"3bb2",x"b34f",x"357c",x"3710",x"3448",x"bbb5",x"0000",x"3a79",x"3bb2"),
(x"b1a1",x"35cc",x"36da",x"2ede",x"3bf4",x"0000",x"3a6e",x"3b61",x"b161",x"35ca",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b161",x"35ca",x"3710",x"30d8",x"3be8",x"0000",x"3a79",x"3b67"),
(x"b783",x"3511",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b7a4",x"351f",x"36da",x"b654",x"bb58",x"8000",x"3a8a",x"3a34",x"b7a4",x"351f",x"3710",x"b64b",x"bb5a",x"0000",x"3a95",x"3a34"),
(x"b72e",x"35d1",x"36da",x"3b4f",x"b67e",x"0000",x"3a97",x"39c6",x"b72d",x"35c9",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b72d",x"35c9",x"3710",x"3a45",x"38f8",x"0000",x"3aa1",x"39c8"),
(x"b2d6",x"3579",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b326",x"357e",x"36da",x"a5e3",x"bbff",x"0000",x"3a6e",x"3bae",x"b326",x"357e",x"3710",x"ad8e",x"bbf8",x"0000",x"3a79",x"3bae"),
(x"b161",x"35ca",x"36da",x"3408",x"3bbd",x"8000",x"3a6e",x"3b67",x"b135",x"35c1",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b135",x"35c1",x"3710",x"3822",x"3ad9",x"0000",x"3a79",x"3b6c"),
(x"b73e",x"350e",x"36da",x"27ae",x"bbfe",x"0000",x"3a8a",x"3a20",x"b783",x"3511",x"36da",x"b33d",x"bbca",x"0000",x"3a8a",x"3a2d",x"b783",x"3511",x"3710",x"afa0",x"bbf1",x"0000",x"3a95",x"3a2d"),
(x"b72d",x"35c9",x"36da",x"3778",x"3b13",x"0000",x"3a97",x"39c8",x"b721",x"35c6",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b721",x"35c6",x"3710",x"2560",x"3bff",x"0000",x"3aa1",x"39ca"),
(x"b2aa",x"356e",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2d6",x"3579",x"36da",x"b287",x"bbd4",x"0000",x"3a6e",x"3ba6",x"b2d6",x"3579",x"3710",x"b4dc",x"bb9f",x"0000",x"3a79",x"3ba6"),
(x"b135",x"35c1",x"36da",x"3934",x"3a13",x"0000",x"3a6e",x"3b6c",x"b116",x"35af",x"36da",x"3bdf",x"31b0",x"8000",x"3a6e",x"3b70",x"b116",x"35af",x"3710",x"3b51",x"3675",x"0000",x"3a79",x"3b70"),
(x"b705",x"351a",x"36da",x"34b8",x"bba4",x"0000",x"3a8a",x"3a15",x"b73e",x"350e",x"36da",x"27ae",x"bbfe",x"0000",x"3a8a",x"3a20",x"b73e",x"350e",x"3710",x"2f57",x"bbf2",x"0000",x"3a95",x"3a20"),
(x"b575",x"3615",x"36da",x"bab5",x"385c",x"0000",x"3a97",x"3a28",x"b568",x"3623",x"36da",x"b810",x"3ae4",x"8000",x"3a97",x"3a2b",x"b568",x"3623",x"3710",x"b919",x"3a29",x"8000",x"3aa1",x"3a2b"),
(x"b938",x"3576",x"36da",x"bbfe",x"a8f0",x"0000",x"3bf8",x"39d0",x"b93a",x"35c9",x"36da",x"bbfe",x"a8f0",x"0000",x"3be9",x"39cf",x"b93a",x"35c9",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3be8",x"39da"),
(x"b261",x"3559",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b2aa",x"356e",x"36da",x"b78b",x"bb0e",x"0000",x"3a6e",x"3ba2",x"b2aa",x"356e",x"3710",x"b7e2",x"baf5",x"0000",x"3a79",x"3ba2"),
(x"b931",x"3629",x"36da",x"23ae",x"3bff",x"0000",x"3be3",x"3a63",x"b8ff",x"3627",x"36da",x"26a7",x"3bff",x"8000",x"3be3",x"3a4f",x"b8ff",x"3627",x"3710",x"2581",x"3bff",x"1553",x"3bd9",x"3a4f"),
(x"b6f1",x"352c",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b705",x"351a",x"36da",x"34b8",x"bba4",x"0000",x"3a8a",x"3a15",x"b705",x"351a",x"3710",x"36ee",x"bb35",x"0000",x"3a95",x"3a15"),
(x"b721",x"35c6",x"36da",x"0cea",x"3c00",x"0000",x"3a97",x"39ca",x"b669",x"35c7",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b669",x"35c7",x"3710",x"a666",x"3bff",x"0000",x"3aa1",x"39ed"),
(x"b22d",x"3552",x"36da",x"ae88",x"bbf5",x"0000",x"3a6e",x"3b94",x"b261",x"3559",x"36da",x"b72e",x"bb26",x"0000",x"3a6e",x"3b9a",x"b261",x"3559",x"3710",x"b5e0",x"bb70",x"8000",x"3a79",x"3b9a"),
(x"b6ef",x"3541",x"36da",x"3be9",x"30b7",x"8000",x"3a8a",x"3a0c",x"b6f1",x"352c",x"36da",x"3a69",x"b8c9",x"068d",x"3a8a",x"3a10",x"b6f1",x"352c",x"3710",x"3b73",x"b5d3",x"868d",x"3a95",x"3a10"),
(x"b669",x"35c7",x"36da",x"abae",x"3bfc",x"0000",x"3a97",x"39ed",x"b63d",x"35cf",x"36da",x"ab45",x"3bfc",x"0000",x"3a97",x"39f5",x"b63d",x"35cf",x"3710",x"affc",x"3bf0",x"0000",x"3aa1",x"39f5"),
(x"b930",x"356e",x"36da",x"b67a",x"bb50",x"0000",x"3bc0",x"3984",x"b938",x"3576",x"36da",x"b67a",x"bb50",x"0000",x"3bbd",x"3982",x"b938",x"3576",x"3710",x"b678",x"bb4d",x"2af3",x"3bb7",x"398a"),
(x"b7a8",x"35f7",x"3710",x"8000",x"0000",x"3c00",x"3a22",x"311a",x"b783",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b790",x"35f3",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3107"),
(x"b34f",x"35bf",x"3710",x"8000",x"0000",x"3c00",x"3a16",x"2a20",x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b351",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b368",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b351",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b340",x"354d",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2a0e"),
(x"b34f",x"357c",x"3710",x"8000",x"0000",x"3c00",x"3a08",x"2a20",x"b351",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b340",x"3c9f",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"2a04",x"b33a",x"3c9a",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"29f9",x"b351",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b783",x"3c68",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b7a8",x"3c75",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a",x"b790",x"3c76",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3107"),
(x"b783",x"3cae",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b77b",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b790",x"3ca0",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3107"),
(x"b40d",x"3c9e",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b368",x"3ca5",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b351",x"3c95",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b351",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b33a",x"3c7c",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2a04",x"b340",x"3c77",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2a0e"),
(x"b351",x"3c81",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b368",x"3c71",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b40d",x"3c78",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"b340",x"35ee",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"2a04",x"b33a",x"35d9",x"3710",x"8000",x"0000",x"3c00",x"3a1c",x"29f9",x"b351",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b783",x"3511",x"3710",x"8000",x"0000",x"3c00",x"39f1",x"30f9",x"b7a8",x"3544",x"3710",x"8000",x"0000",x"3c00",x"39fc",x"311a",x"b790",x"3548",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"3107"),
(x"b783",x"362a",x"3710",x"8000",x"0000",x"3c00",x"3a2d",x"30f9",x"b77b",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"30f2",x"b790",x"35f3",x"3710",x"8000",x"0000",x"3c00",x"3a20",x"3107"),
(x"b40d",x"35e8",x"3710",x"8000",x"0000",x"3c00",x"3a1f",x"2b8b",x"b368",x"3605",x"3710",x"8000",x"0000",x"3c00",x"3a25",x"2a4d",x"b351",x"35c7",x"3710",x"8000",x"0000",x"3c00",x"3a18",x"2a22"),
(x"b351",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b33a",x"3562",x"3710",x"8000",x"0000",x"3c00",x"3a01",x"2a04",x"b340",x"354d",x"3710",x"8000",x"0000",x"3c00",x"39fd",x"2a0e"),
(x"b351",x"3574",x"3710",x"8000",x"0000",x"3c00",x"3a05",x"2a27",x"b368",x"3536",x"3710",x"8000",x"0000",x"3c00",x"39f9",x"2a4d",x"b40d",x"3553",x"3710",x"8000",x"0000",x"3c00",x"39ff",x"2b8b"),
(x"3a2c",x"3d32",x"36fb",x"3c00",x"0000",x"0000",x"3b04",x"3ac8",x"3a2c",x"4062",x"36fb",x"3c00",x"0000",x"0000",x"3b04",x"3b93",x"3a2c",x"3d32",x"368e",x"3c00",x"0000",x"0000",x"3b0c",x"3ac8"),
(x"2c34",x"3d32",x"368e",x"bc00",x"8000",x"0000",x"3782",x"1d2d",x"2c34",x"4062",x"368e",x"bc00",x"8000",x"0000",x"3782",x"3512",x"2c34",x"3d32",x"36fb",x"bc00",x"8000",x"0000",x"37b6",x"1d2d"),
(x"3193",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3bc7",x"382d",x"394e",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3bc7",x"3920",x"3193",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3bcd",x"382d"),
(x"3a2c",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3bf2",x"282d",x"2c34",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3b1b",x"282d",x"3a2c",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3bf2",x"288d"),
(x"2c34",x"4062",x"368e",x"0000",x"3c00",x"0000",x"3b1b",x"26d5",x"3a2c",x"4062",x"368e",x"0000",x"3c00",x"0000",x"3bf2",x"26d5",x"2c34",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"3b1b",x"2613"),
(x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d",x"3a2c",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3973",x"3962",x"3dde",x"36fb",x"0000",x"0000",x"3c00",x"3b93",x"39a8"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"3009",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3adf",x"39fb",x"3004",x"3eee",x"36fb",x"868d",x"0000",x"3c00",x"3adf",x"39fc"),
(x"394e",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"399a",x"3a2c",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3973",x"3193",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"399a"),
(x"394e",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"3a66",x"3193",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"3a66",x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d"),
(x"3193",x"3dae",x"36d0",x"0000",x"0000",x"3c00",x"386d",x"3bf9",x"3193",x"4024",x"36d0",x"0000",x"0000",x"3c00",x"386d",x"3adb",x"394e",x"3dae",x"36d0",x"0000",x"0000",x"3c00",x"374c",x"3bf9"),
(x"3193",x"3dbd",x"36fb",x"3c00",x"0000",x"0000",x"3b68",x"3aca",x"3193",x"3dc7",x"36e5",x"3c00",x"0000",x"0000",x"3b5e",x"3acf",x"3193",x"3dae",x"36d0",x"3c00",x"0000",x"0000",x"3b78",x"3ad4"),
(x"394e",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3b76",x"3542",x"3193",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3aed",x"3542",x"394e",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3b76",x"3556"),
(x"3141",x"4015",x"36fb",x"396d",x"9af6",x"39e0",x"354c",x"3742",x"316f",x"401e",x"36fb",x"39bc",x"b304",x"394a",x"3548",x"372f",x"3193",x"4016",x"36d7",x"394c",x"a074",x"39fd",x"353f",x"373f"),
(x"3193",x"3dbd",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"399e",x"3193",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"399a",x"3160",x"3dc9",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"39a2"),
(x"3193",x"401e",x"36e4",x"3a1e",x"b321",x"38d5",x"3541",x"3730",x"316f",x"401e",x"36fb",x"39bc",x"b304",x"394a",x"3548",x"372f",x"3193",x"4022",x"36fb",x"39d6",x"b5ae",x"38ac",x"3545",x"3725"),
(x"3193",x"3dae",x"36d0",x"3c00",x"0000",x"0000",x"3b78",x"3ad4",x"3193",x"3dd5",x"36d4",x"3c00",x"0000",x"0000",x"3b4f",x"3ad3",x"3193",x"4024",x"36d0",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4"),
(x"3193",x"401e",x"36e4",x"3c00",x"0000",x"0000",x"3b3f",x"3ad4",x"3193",x"4022",x"36fb",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4",x"3193",x"4024",x"36d0",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4"),
(x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973",x"3143",x"3dd7",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"39a6",x"3160",x"3dc9",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"39a2"),
(x"3143",x"3dd7",x"36fb",x"3993",x"1c9b",x"39bd",x"354c",x"38c9",x"3141",x"4015",x"36fb",x"396d",x"9af6",x"39e0",x"354c",x"3742",x"3193",x"3dd5",x"36d4",x"396e",x"1b2b",x"39df",x"353f",x"38ca"),
(x"3143",x"3dd7",x"36fb",x"3993",x"1c9b",x"39bd",x"354c",x"38c9",x"3193",x"3dd5",x"36d4",x"396e",x"1b2b",x"39df",x"353f",x"38ca",x"3160",x"3dc9",x"36fb",x"3988",x"33a8",x"3973",x"354a",x"38cf"),
(x"3193",x"3dc7",x"36e5",x"396c",x"347c",x"396f",x"3542",x"38d1",x"3193",x"3dbd",x"36fb",x"3969",x"359e",x"392e",x"3546",x"38d6",x"3160",x"3dc9",x"36fb",x"3988",x"33a8",x"3973",x"354a",x"38cf"),
(x"394e",x"4024",x"36d0",x"ba68",x"217a",x"b8c9",x"3a93",x"34bd",x"394e",x"4024",x"36fb",x"bbf4",x"2eb8",x"0000",x"3a92",x"34d1",x"394d",x"4023",x"36fb",x"bbfe",x"276c",x"a4f7",x"3a95",x"34d1"),
(x"394d",x"3dc6",x"36dd",x"bbff",x"a074",x"a611",x"3b18",x"34c0",x"394d",x"3dbb",x"36fb",x"bbff",x"a3a0",x"a0d0",x"3b1b",x"34c2",x"394e",x"3dae",x"36d0",x"3b8d",x"a187",x"b543",x"3b1d",x"34bd"),
(x"394d",x"3dc6",x"36dd",x"ba1a",x"3321",x"38da",x"3594",x"372e",x"3959",x"3dc6",x"36fb",x"ba1d",x"31d2",x"38f2",x"359c",x"372e",x"394d",x"3dbb",x"36fb",x"b9d1",x"35ef",x"389f",x"3599",x"3722"),
(x"394d",x"4016",x"36d8",x"bbf1",x"1553",x"afa7",x"3aaf",x"34c2",x"394d",x"3ddc",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b13",x"34c1",x"394e",x"4024",x"36d0",x"ba68",x"217a",x"b8c9",x"3a93",x"34bd"),
(x"3962",x"3dde",x"36fb",x"b9b6",x"128d",x"3999",x"359f",x"3747",x"3959",x"3dc6",x"36fb",x"ba1d",x"31d2",x"38f2",x"359c",x"372e",x"394d",x"3ddc",x"36ca",x"ba14",x"1cd0",x"3932",x"3590",x"3744"),
(x"3961",x"4016",x"36fb",x"b935",x"9d6d",x"3a12",x"359c",x"38c9",x"3962",x"3dde",x"36fb",x"b9b6",x"128d",x"3999",x"359f",x"3747",x"394d",x"4016",x"36d8",x"b9b2",x"9dbc",x"399d",x"3590",x"38c9"),
(x"3961",x"4016",x"36fb",x"b935",x"9d6d",x"3a12",x"359c",x"38c9",x"394d",x"4016",x"36d8",x"b9b2",x"9dbc",x"399d",x"3590",x"38c9",x"3958",x"401d",x"36fb",x"b94f",x"b2e4",x"39ba",x"3599",x"38d0"),
(x"394d",x"401d",x"36e5",x"b97d",x"b372",x"3982",x"3592",x"38d0",x"394d",x"4023",x"36fb",x"b958",x"b562",x"394e",x"3595",x"38d6",x"3958",x"401d",x"36fb",x"b94f",x"b2e4",x"39ba",x"3599",x"38d0"),
(x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973",x"2ee6",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3ad9",x"39fb",x"2f02",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39ef"),
(x"2c34",x"3d32",x"368e",x"0000",x"8000",x"bc00",x"3bf4",x"30be",x"3a2c",x"3d32",x"368e",x"0000",x"8000",x"bc00",x"3b38",x"30be",x"2c34",x"4062",x"368e",x"0000",x"8000",x"bc00",x"3bf4",x"3418"),
(x"2fe5",x"3ee4",x"36fb",x"bb7d",x"359e",x"0000",x"3b44",x"3a1d",x"2fe5",x"3ee4",x"36b4",x"bb3f",x"36c6",x"8000",x"3b44",x"3a14",x"3009",x"3eea",x"36fb",x"bb8f",x"3538",x"0000",x"3b41",x"3a1d"),
(x"2f02",x"3ec3",x"36fb",x"a460",x"3bff",x"0000",x"3b77",x"3a2c",x"2f02",x"3ec3",x"36b4",x"a460",x"3bff",x"0000",x"3b6d",x"3a2c",x"3025",x"3ec3",x"36fb",x"a460",x"3bff",x"0000",x"3b77",x"3a36"),
(x"2f19",x"3eef",x"36fb",x"3727",x"bb27",x"0000",x"3b36",x"3a1d",x"2f19",x"3eef",x"36b4",x"393c",x"ba0c",x"0000",x"3b36",x"3a14",x"2ee6",x"3eea",x"36fb",x"3bcf",x"b2e7",x"0000",x"3b33",x"3a1d"),
(x"3009",x"3eea",x"36fb",x"bb8f",x"3538",x"0000",x"3b41",x"3a1d",x"3009",x"3eea",x"36b4",x"bbef",x"3012",x"0000",x"3b41",x"3a14",x"3004",x"3eee",x"36fb",x"baa8",x"b870",x"0000",x"3b3e",x"3a1d"),
(x"3025",x"3ec3",x"36fb",x"bbcb",x"b335",x"0000",x"3b56",x"3a1d",x"3025",x"3ec3",x"36b4",x"bbcb",x"b335",x"0000",x"3b56",x"3a14",x"2fda",x"3ee2",x"36fb",x"bbd4",x"b28e",x"868d",x"3b45",x"3a1d"),
(x"2ee6",x"3eea",x"36fb",x"3bcf",x"b2e7",x"0000",x"3b33",x"3a1d",x"2ee6",x"3eea",x"36b4",x"3bf2",x"2f67",x"0000",x"3b33",x"3a14",x"2f10",x"3ee4",x"36fb",x"3bf6",x"2e14",x"0000",x"3b2f",x"3a1d"),
(x"3004",x"3eee",x"36fb",x"baa8",x"b870",x"0000",x"3b3e",x"3a1d",x"3004",x"3eee",x"36b4",x"b8fa",x"ba42",x"0000",x"3b3e",x"3a14",x"2f99",x"3ef2",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a1d"),
(x"2fda",x"3ee2",x"36fb",x"bbd4",x"b28e",x"868d",x"3b45",x"3a1d",x"2fda",x"3ee2",x"36b4",x"bbe8",x"b0e2",x"0000",x"3b45",x"3a14",x"2fe5",x"3ee4",x"36fb",x"bb7d",x"359e",x"0000",x"3b44",x"3a1d"),
(x"2f10",x"3ee4",x"36fb",x"3bf6",x"2e14",x"0000",x"3b2f",x"3a1d",x"2f10",x"3ee4",x"36b4",x"3bff",x"2231",x"068d",x"3b2f",x"3a14",x"2f02",x"3ec3",x"36fb",x"3bff",x"a6cf",x"0000",x"3b1e",x"3a1d"),
(x"2f99",x"3ef2",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a1d",x"2f99",x"3ef2",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a14",x"2f19",x"3eef",x"36fb",x"3727",x"bb27",x"0000",x"3b36",x"3a1d"),
(x"3a2c",x"4062",x"36fb",x"3c00",x"0000",x"0000",x"3b04",x"3b93",x"3a2c",x"4062",x"368e",x"3c00",x"0000",x"0000",x"3b0c",x"3b93",x"3a2c",x"3d32",x"368e",x"3c00",x"0000",x"0000",x"3b0c",x"3ac8"),
(x"2c34",x"4062",x"368e",x"bc00",x"8000",x"0000",x"3782",x"3512",x"2c34",x"4062",x"36fb",x"bc00",x"8000",x"0000",x"37b6",x"3512",x"2c34",x"3d32",x"36fb",x"bc00",x"8000",x"0000",x"37b6",x"1d2d"),
(x"394e",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3bc7",x"3920",x"394e",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3bcd",x"3920",x"3193",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3bcd",x"382d"),
(x"2c34",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3b1b",x"282d",x"2c34",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3b1b",x"288d",x"3a2c",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3bf2",x"288d"),
(x"3a2c",x"4062",x"368e",x"0000",x"3c00",x"0000",x"3bf2",x"26d5",x"3a2c",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"3bf2",x"2613",x"2c34",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"3b1b",x"2613"),
(x"3959",x"3dc6",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"39a1",x"394e",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"399a",x"394d",x"3dbb",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"399d"),
(x"3959",x"3dc6",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"39a1",x"3a2c",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3973",x"394e",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"399a"),
(x"3958",x"401d",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"3a62",x"394e",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"3a66",x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d"),
(x"3958",x"401d",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"3a62",x"394d",x"4023",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"3a66",x"394e",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3b90",x"3a66"),
(x"3a2c",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3973",x"3959",x"3dc6",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"39a1",x"3962",x"3dde",x"36fb",x"0000",x"0000",x"3c00",x"3b93",x"39a8"),
(x"3961",x"4016",x"36fb",x"0000",x"0000",x"3c00",x"3b93",x"3a5e",x"3958",x"401d",x"36fb",x"0000",x"0000",x"3c00",x"3b92",x"3a62",x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d"),
(x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d",x"3962",x"3dde",x"36fb",x"0000",x"0000",x"3c00",x"3b93",x"39a8",x"3961",x"4016",x"36fb",x"0000",x"0000",x"3c00",x"3b93",x"3a5e"),
(x"316f",x"401e",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"3a62",x"3193",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"3a66",x"3193",x"4022",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"3a65"),
(x"316f",x"401e",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"3a62",x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d",x"3193",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"3a66"),
(x"2ee6",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3ad9",x"39fb",x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973",x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d"),
(x"2f19",x"3eef",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39fc",x"2ee6",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3ad9",x"39fb",x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"3143",x"3dd7",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"39a6",x"3025",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ae0",x"39ef"),
(x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d",x"316f",x"401e",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"3a62",x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"2f19",x"3eef",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39fc",x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"2f99",x"3ef2",x"36fb",x"0000",x"0000",x"3c00",x"3add",x"39fd",x"2f19",x"3eef",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39fc"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"3004",x"3eee",x"36fb",x"868d",x"0000",x"3c00",x"3adf",x"39fc",x"2f99",x"3ef2",x"36fb",x"0000",x"0000",x"3c00",x"3add",x"39fd"),
(x"3009",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3adf",x"39fb",x"2fda",x"3ee2",x"36fb",x"0000",x"0000",x"3c00",x"3ade",x"39f8",x"2fe5",x"3ee4",x"36fb",x"068d",x"0000",x"3c00",x"3ade",x"39f9"),
(x"3009",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3adf",x"39fb",x"3025",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ae0",x"39ef",x"2fda",x"3ee2",x"36fb",x"0000",x"0000",x"3c00",x"3ade",x"39f8"),
(x"3141",x"4015",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"3a5d",x"3025",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ae0",x"39ef",x"3009",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3adf",x"39fb"),
(x"3a2c",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3973",x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973",x"3193",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"399a"),
(x"3193",x"4024",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"3a66",x"2c34",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3a8d",x"3a2c",x"4062",x"36fb",x"0000",x"0000",x"3c00",x"3bb4",x"3a8d"),
(x"3193",x"4024",x"36d0",x"0000",x"0000",x"3c00",x"386d",x"3adb",x"394e",x"4024",x"36d0",x"0000",x"0000",x"3c00",x"374c",x"3adb",x"394e",x"3dae",x"36d0",x"0000",x"0000",x"3c00",x"374c",x"3bf9"),
(x"3193",x"3dae",x"36d0",x"3c00",x"0000",x"0000",x"3b78",x"3ad4",x"3193",x"3dae",x"36fb",x"3c00",x"0000",x"0000",x"3b78",x"3aca",x"3193",x"3dbd",x"36fb",x"3c00",x"0000",x"0000",x"3b68",x"3aca"),
(x"3193",x"3dc7",x"36e5",x"3c00",x"0000",x"0000",x"3b5e",x"3acf",x"3193",x"3dd5",x"36d4",x"3c00",x"0000",x"0000",x"3b4f",x"3ad3",x"3193",x"3dae",x"36d0",x"3c00",x"0000",x"0000",x"3b78",x"3ad4"),
(x"3193",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3aed",x"3542",x"3193",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3aed",x"3556",x"394e",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3b76",x"3556"),
(x"316f",x"401e",x"36fb",x"39bc",x"b304",x"394a",x"3548",x"372f",x"3193",x"401e",x"36e4",x"3a1e",x"b321",x"38d5",x"3541",x"3730",x"3193",x"4016",x"36d7",x"394c",x"a074",x"39fd",x"353f",x"373f"),
(x"3193",x"3dae",x"36fb",x"0000",x"0000",x"3c00",x"3aef",x"399a",x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973",x"3160",x"3dc9",x"36fb",x"0000",x"0000",x"3c00",x"3aed",x"39a2"),
(x"3193",x"3dd5",x"36d4",x"3c00",x"0000",x"0000",x"3b4f",x"3ad3",x"3193",x"4016",x"36d7",x"3c00",x"0000",x"0000",x"3b3f",x"3ad4",x"3193",x"4024",x"36d0",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4"),
(x"3193",x"4022",x"36fb",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4",x"3193",x"4024",x"36fb",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4",x"3193",x"4024",x"36d0",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4"),
(x"3193",x"4024",x"36d0",x"3c00",x"0000",x"0000",x"3b3e",x"3ad4",x"3193",x"4016",x"36d7",x"3c00",x"0000",x"0000",x"3b3f",x"3ad4",x"3193",x"401e",x"36e4",x"3c00",x"0000",x"0000",x"3b3f",x"3ad4"),
(x"3141",x"4015",x"36fb",x"396d",x"9af6",x"39e0",x"354c",x"3742",x"3193",x"4016",x"36d7",x"394c",x"a074",x"39fd",x"353f",x"373f",x"3193",x"3dd5",x"36d4",x"396e",x"1b2b",x"39df",x"353f",x"38ca"),
(x"3193",x"3dd5",x"36d4",x"396e",x"1b2b",x"39df",x"353f",x"38ca",x"3193",x"3dc7",x"36e5",x"396c",x"347c",x"396f",x"3542",x"38d1",x"3160",x"3dc9",x"36fb",x"3988",x"33a8",x"3973",x"354a",x"38cf"),
(x"394d",x"401d",x"36e5",x"bbfe",x"2104",x"a780",x"3aa0",x"34c7",x"394d",x"4016",x"36d8",x"bbf1",x"1553",x"afa7",x"3aaf",x"34c2",x"394e",x"4024",x"36d0",x"ba68",x"217a",x"b8c9",x"3a93",x"34bd"),
(x"394e",x"4024",x"36d0",x"ba68",x"217a",x"b8c9",x"3a93",x"34bd",x"394d",x"4023",x"36fb",x"bbfe",x"276c",x"a4f7",x"3a95",x"34d1",x"394d",x"401d",x"36e5",x"bbfe",x"2104",x"a780",x"3aa0",x"34c7"),
(x"394d",x"3dbb",x"36fb",x"bbff",x"a3a0",x"a0d0",x"3b1b",x"34c2",x"394e",x"3dae",x"36fb",x"bbff",x"a5e9",x"0000",x"3b1d",x"34c1",x"394e",x"3dae",x"36d0",x"3b8d",x"a187",x"b543",x"3b1d",x"34bd"),
(x"394e",x"3dae",x"36d0",x"3b8d",x"a187",x"b543",x"3b1d",x"34bd",x"394d",x"3ddc",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b13",x"34c1",x"394d",x"3dc6",x"36dd",x"bbff",x"a074",x"a611",x"3b18",x"34c0"),
(x"394d",x"3ddc",x"36ca",x"b9ed",x"90ea",x"b95f",x"3b13",x"34c1",x"394e",x"3dae",x"36d0",x"3b8d",x"a187",x"b543",x"3b1d",x"34bd",x"394e",x"4024",x"36d0",x"ba68",x"217a",x"b8c9",x"3a93",x"34bd"),
(x"3959",x"3dc6",x"36fb",x"ba1d",x"31d2",x"38f2",x"359c",x"372e",x"394d",x"3dc6",x"36dd",x"ba1a",x"3321",x"38da",x"3594",x"372e",x"394d",x"3ddc",x"36ca",x"ba14",x"1cd0",x"3932",x"3590",x"3744"),
(x"3962",x"3dde",x"36fb",x"b9b6",x"128d",x"3999",x"359f",x"3747",x"394d",x"3ddc",x"36ca",x"ba14",x"1cd0",x"3932",x"3590",x"3744",x"394d",x"4016",x"36d8",x"b9b2",x"9dbc",x"399d",x"3590",x"38c9"),
(x"394d",x"4016",x"36d8",x"b9b2",x"9dbc",x"399d",x"3590",x"38c9",x"394d",x"401d",x"36e5",x"b97d",x"b372",x"3982",x"3592",x"38d0",x"3958",x"401d",x"36fb",x"b94f",x"b2e4",x"39ba",x"3599",x"38d0"),
(x"2f02",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39ef",x"3143",x"3dd7",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"39a6",x"2c34",x"3d32",x"36fb",x"0000",x"0000",x"3c00",x"3acb",x"3973"),
(x"2f02",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39ef",x"3025",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ae0",x"39ef",x"3143",x"3dd7",x"36fb",x"0000",x"0000",x"3c00",x"3aec",x"39a6"),
(x"2ee6",x"3eea",x"36fb",x"0000",x"0000",x"3c00",x"3ad9",x"39fb",x"2f10",x"3ee4",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39f9",x"2f02",x"3ec3",x"36fb",x"0000",x"0000",x"3c00",x"3ada",x"39ef"),
(x"3a2c",x"3d32",x"368e",x"0000",x"8000",x"bc00",x"3b38",x"30be",x"3a2c",x"4062",x"368e",x"0000",x"8000",x"bc00",x"3b38",x"3418",x"2c34",x"4062",x"368e",x"0000",x"8000",x"bc00",x"3bf4",x"3418"),
(x"2fe5",x"3ee4",x"36b4",x"bb3f",x"36c6",x"8000",x"3b44",x"3a14",x"3009",x"3eea",x"36b4",x"bbef",x"3012",x"0000",x"3b41",x"3a14",x"3009",x"3eea",x"36fb",x"bb8f",x"3538",x"0000",x"3b41",x"3a1d"),
(x"2f02",x"3ec3",x"36b4",x"a460",x"3bff",x"0000",x"3b6d",x"3a2c",x"3025",x"3ec3",x"36b4",x"a460",x"3bff",x"0000",x"3b6d",x"3a36",x"3025",x"3ec3",x"36fb",x"a460",x"3bff",x"0000",x"3b77",x"3a36"),
(x"2f19",x"3eef",x"36b4",x"393c",x"ba0c",x"0000",x"3b36",x"3a14",x"2ee6",x"3eea",x"36b4",x"3bf2",x"2f67",x"0000",x"3b33",x"3a14",x"2ee6",x"3eea",x"36fb",x"3bcf",x"b2e7",x"0000",x"3b33",x"3a1d"),
(x"3009",x"3eea",x"36b4",x"bbef",x"3012",x"0000",x"3b41",x"3a14",x"3004",x"3eee",x"36b4",x"b8fa",x"ba42",x"0000",x"3b3e",x"3a14",x"3004",x"3eee",x"36fb",x"baa8",x"b870",x"0000",x"3b3e",x"3a1d"),
(x"3025",x"3ec3",x"36b4",x"bbcb",x"b335",x"0000",x"3b56",x"3a14",x"2fda",x"3ee2",x"36b4",x"bbe8",x"b0e2",x"0000",x"3b45",x"3a14",x"2fda",x"3ee2",x"36fb",x"bbd4",x"b28e",x"868d",x"3b45",x"3a1d"),
(x"2ee6",x"3eea",x"36b4",x"3bf2",x"2f67",x"0000",x"3b33",x"3a14",x"2f10",x"3ee4",x"36b4",x"3bff",x"2231",x"068d",x"3b2f",x"3a14",x"2f10",x"3ee4",x"36fb",x"3bf6",x"2e14",x"0000",x"3b2f",x"3a1d"),
(x"3004",x"3eee",x"36b4",x"b8fa",x"ba42",x"0000",x"3b3e",x"3a14",x"2f99",x"3ef2",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a14",x"2f99",x"3ef2",x"36fb",x"b32d",x"bbcb",x"0000",x"3b3a",x"3a1d"),
(x"2fda",x"3ee2",x"36b4",x"bbe8",x"b0e2",x"0000",x"3b45",x"3a14",x"2fe5",x"3ee4",x"36b4",x"bb3f",x"36c6",x"8000",x"3b44",x"3a14",x"2fe5",x"3ee4",x"36fb",x"bb7d",x"359e",x"0000",x"3b44",x"3a1d"),
(x"2f10",x"3ee4",x"36b4",x"3bff",x"2231",x"068d",x"3b2f",x"3a14",x"2f02",x"3ec3",x"36b4",x"3bff",x"a6cf",x"0000",x"3b1e",x"3a14",x"2f02",x"3ec3",x"36fb",x"3bff",x"a6cf",x"0000",x"3b1e",x"3a1d"),
(x"2f99",x"3ef2",x"36b4",x"28d9",x"bbfe",x"0000",x"3b3a",x"3a14",x"2f19",x"3eef",x"36b4",x"393c",x"ba0c",x"0000",x"3b36",x"3a14",x"2f19",x"3eef",x"36fb",x"3727",x"bb27",x"0000",x"3b36",x"3a1d"),
(x"2f10",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7d",x"350c",x"2fe5",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7c",x"3519",x"2fda",x"3ee2",x"36b4",x"0000",x"0000",x"3c00",x"3a7e",x"3519"),
(x"303e",x"3ee5",x"3718",x"3bb8",x"b22d",x"31b0",x"38f7",x"303b",x"304f",x"3ee5",x"36eb",x"3ba3",x"b453",x"2fdf",x"3902",x"302b",x"3033",x"3ee0",x"3715",x"3bf4",x"2da3",x"2b3e",x"38f6",x"3025"),
(x"303e",x"3ee5",x"3718",x"3bb8",x"b22d",x"31b0",x"38f7",x"303b",x"3048",x"3eed",x"3715",x"3bda",x"2e4f",x"312f",x"38fa",x"305a",x"304f",x"3ee5",x"36eb",x"3ba3",x"b453",x"2fdf",x"3902",x"302b"),
(x"3048",x"3eed",x"3715",x"3bda",x"2e4f",x"312f",x"38fa",x"305a",x"3027",x"3ef4",x"3714",x"3a0a",x"3915",x"3126",x"38fd",x"307d",x"3054",x"3eed",x"36eb",x"3b7a",x"3531",x"30a8",x"3905",x"304d"),
(x"3027",x"3ef4",x"3714",x"3a0a",x"3915",x"3126",x"38fd",x"307d",x"2fca",x"3ef8",x"3714",x"3235",x"3bc0",x"30e0",x"38fe",x"30a4",x"302b",x"3ef6",x"36eb",x"38c7",x"3a49",x"310b",x"3907",x"3079"),
(x"2fca",x"3ef8",x"3714",x"3235",x"3bc0",x"30e0",x"38fe",x"30a4",x"2ef2",x"3ef7",x"3714",x"b35f",x"3baf",x"30fd",x"38ff",x"30df",x"2fcc",x"3efa",x"36eb",x"23ae",x"3bec",x"306c",x"3908",x"30a1"),
(x"2ef2",x"3ef7",x"3714",x"b35f",x"3baf",x"30fd",x"38ff",x"30df",x"2e86",x"3ef1",x"3715",x"ba37",x"38de",x"311d",x"38fe",x"3104",x"2ed8",x"3ef8",x"36eb",x"b6e0",x"3b1c",x"3118",x"3909",x"30e3"),
(x"2e86",x"3ef1",x"3715",x"ba37",x"38de",x"311d",x"38fe",x"3104",x"2e63",x"3eea",x"3715",x"bbf2",x"2495",x"2f43",x"38fd",x"3126",x"2e6e",x"3ef2",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3909",x"310b"),
(x"2e80",x"3ee3",x"3715",x"bb87",x"b537",x"2d81",x"38fc",x"3144",x"2e6b",x"3ee3",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3906",x"314b",x"2e63",x"3eea",x"3715",x"bbf2",x"2495",x"2f43",x"38fd",x"3126"),
(x"2e96",x"3ede",x"3717",x"bbff",x"2481",x"2487",x"38fa",x"3158",x"2e93",x"3ede",x"36eb",x"bbfd",x"212b",x"29e6",x"3905",x"3161",x"2e80",x"3ee3",x"3715",x"bb87",x"b537",x"2d81",x"38fc",x"3144"),
(x"2e34",x"3ec3",x"36eb",x"bb76",x"3593",x"2dee",x"3900",x"31de",x"2e6c",x"3ec4",x"36eb",x"bb9b",x"34d2",x"2ca5",x"3900",x"31ce",x"2e3f",x"3ec2",x"3714",x"bb74",x"35a6",x"2d5e",x"38f6",x"31d7"),
(x"2f2c",x"3ee5",x"36eb",x"3ba6",x"341e",x"3066",x"38ef",x"2dd9",x"2f22",x"3edf",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38ea",x"2ddb",x"2f16",x"3ee4",x"3716",x"3bb3",x"33ed",x"2eeb",x"38ef",x"2e30"),
(x"2f22",x"3edf",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38ea",x"2ddb",x"2f2a",x"3ec5",x"36eb",x"3a79",x"3840",x"3401",x"38ce",x"2de0",x"2f13",x"3edf",x"3718",x"3bf1",x"95bc",x"2fb6",x"38ea",x"2e35"),
(x"3072",x"3eb8",x"3715",x"33c8",x"bbc2",x"236c",x"38e5",x"2f03",x"306e",x"3ec3",x"3715",x"3bb4",x"33e7",x"2ed7",x"38e9",x"2f58",x"3079",x"3eb9",x"36eb",x"3409",x"bbbc",x"27e2",x"38ee",x"2edd"),
(x"2e32",x"3eb9",x"3714",x"af03",x"bbf3",x"23ef",x"38f4",x"31ff",x"2e24",x"3eb8",x"36eb",x"b6d0",x"bb39",x"2ab1",x"38fd",x"320b",x"2e3f",x"3ec2",x"3714",x"bb74",x"35a6",x"2d5e",x"38f6",x"31d7"),
(x"2fd9",x"3edf",x"3716",x"bbce",x"b2bb",x"2b41",x"391c",x"2e40",x"2fc8",x"3ee0",x"36eb",x"bbd3",x"b208",x"2da6",x"391d",x"2de9",x"2fd7",x"3ee3",x"3715",x"bb88",x"3531",x"2dc2",x"3918",x"2e3b"),
(x"2fc7",x"3ee4",x"36ee",x"bb70",x"358e",x"2fc0",x"3918",x"2ded",x"2ffa",x"3ee8",x"36ee",x"bb20",x"3725",x"2d51",x"3913",x"2ded",x"2fd7",x"3ee3",x"3715",x"bb88",x"3531",x"2dc2",x"3918",x"2e3b"),
(x"2ffa",x"3ee8",x"36ee",x"bb20",x"3725",x"2d51",x"3913",x"2ded",x"2fff",x"3eec",x"36ee",x"bb1d",x"b747",x"2911",x"390e",x"2dec",x"3005",x"3ee9",x"3717",x"bbd6",x"323b",x"2a8a",x"3911",x"2e3e"),
(x"2f3e",x"3ef0",x"36ee",x"314a",x"bbe2",x"a87e",x"38ff",x"2de6",x"2f00",x"3eec",x"36ee",x"3a67",x"b8c6",x"2a76",x"38f9",x"2de4",x"2f3a",x"3ef0",x"3715",x"36a0",x"bb47",x"2074",x"38ff",x"2e34"),
(x"2fc8",x"3ee0",x"36eb",x"bbd3",x"b208",x"2da6",x"391d",x"2de9",x"2fd9",x"3edf",x"3716",x"bbce",x"b2bb",x"2b41",x"391c",x"2e40",x"3016",x"3ec6",x"36eb",x"bbe6",x"2cac",x"3077",x"3939",x"2dfc"),
(x"2e77",x"3ec4",x"3717",x"a984",x"a0c2",x"3bfd",x"3980",x"3272",x"2e32",x"3eb9",x"3714",x"a745",x"ad9b",x"3bf7",x"397d",x"3257",x"2e3f",x"3ec2",x"3714",x"b3e6",x"2587",x"3bc0",x"397e",x"326d"),
(x"3056",x"3ec4",x"3718",x"26a1",x"97c8",x"3bff",x"3994",x"3272",x"306e",x"3ec3",x"3715",x"33f3",x"1d38",x"3bbf",x"3995",x"3270",x"3072",x"3eb8",x"3715",x"2081",x"ad9e",x"3bf8",x"3996",x"3257"),
(x"303e",x"3ee5",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3992",x"32bf",x"3033",x"3ee0",x"3715",x"21a1",x"23fc",x"3bff",x"3991",x"32b4",x"2fd7",x"3ee3",x"3715",x"a8d3",x"a80e",x"3bfd",x"398c",x"32bc"),
(x"3048",x"3eed",x"3715",x"1e8d",x"2bdf",x"3bfc",x"3993",x"32d2",x"303e",x"3ee5",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3992",x"32bf",x"3005",x"3ee9",x"3717",x"a511",x"281b",x"3bfe",x"398e",x"32c8"),
(x"3027",x"3ef4",x"3714",x"a63f",x"27c1",x"3bfe",x"3990",x"32e3",x"3048",x"3eed",x"3715",x"1e8d",x"2bdf",x"3bfc",x"3993",x"32d2",x"2fff",x"3eed",x"3716",x"a52b",x"2c96",x"3bfa",x"398e",x"32d3"),
(x"2fca",x"3ef8",x"3714",x"2187",x"a0ea",x"3bff",x"398c",x"32ed",x"3027",x"3ef4",x"3714",x"a63f",x"27c1",x"3bfe",x"3990",x"32e3",x"2fc2",x"3eef",x"3713",x"991e",x"9cea",x"3c00",x"398b",x"32d8"),
(x"2ef2",x"3ef7",x"3714",x"9dd6",x"248e",x"3bff",x"3984",x"32ea",x"2fca",x"3ef8",x"3714",x"2187",x"a0ea",x"3bff",x"398c",x"32ed",x"2f3a",x"3ef0",x"3715",x"1c81",x"1953",x"3c00",x"3987",x"32d9"),
(x"2e86",x"3ef1",x"3715",x"2793",x"184d",x"3bff",x"3980",x"32dc",x"2ef2",x"3ef7",x"3714",x"9dd6",x"248e",x"3bff",x"3984",x"32ea",x"2ef1",x"3eec",x"3714",x"1da1",x"252b",x"3bff",x"3984",x"32cf"),
(x"2e86",x"3ef1",x"3715",x"2793",x"184d",x"3bff",x"3980",x"32dc",x"2ef1",x"3eec",x"3714",x"1da1",x"252b",x"3bff",x"3984",x"32cf",x"2e63",x"3eea",x"3715",x"1818",x"26bb",x"3bff",x"397f",x"32ca"),
(x"2e63",x"3eea",x"3715",x"1818",x"26bb",x"3bff",x"397f",x"32ca",x"2eed",x"3ee8",x"3716",x"a338",x"267a",x"3bff",x"3984",x"32c7",x"2e80",x"3ee3",x"3715",x"a645",x"29e0",x"3bfd",x"3980",x"32ba"),
(x"2e96",x"3ede",x"3717",x"a7d5",x"236c",x"3bfe",x"3981",x"32af",x"2e80",x"3ee3",x"3715",x"a645",x"29e0",x"3bfd",x"3980",x"32ba",x"2f13",x"3edf",x"3718",x"a793",x"243f",x"3bfe",x"3985",x"32b2"),
(x"2f0c",x"3ec2",x"3718",x"a3ae",x"ac2f",x"3bfb",x"3985",x"326e",x"2e77",x"3ec4",x"3717",x"a984",x"a0c2",x"3bfd",x"3980",x"3272",x"2f13",x"3edf",x"3718",x"a793",x"243f",x"3bfe",x"3985",x"32b2"),
(x"2f00",x"3eec",x"36ee",x"3a67",x"b8c6",x"2a76",x"38f9",x"2de4",x"2efa",x"3ee8",x"36ee",x"3b84",x"3534",x"2e9f",x"38f5",x"2de3",x"2ef1",x"3eec",x"3714",x"3b37",x"b6c3",x"2d61",x"38f8",x"2e30"),
(x"3056",x"3ec4",x"3718",x"3ba4",x"33dc",x"313e",x"38e9",x"2f72",x"3033",x"3ee0",x"3715",x"3bf4",x"2da3",x"2b3e",x"38f6",x"3025",x"3065",x"3ec5",x"36eb",x"3baa",x"3479",x"2b93",x"38f4",x"2f49"),
(x"3077",x"3ec4",x"36eb",x"3bc6",x"328d",x"2f71",x"38f3",x"2f37",x"306e",x"3ec3",x"3715",x"3bb4",x"33e7",x"2ed7",x"38e9",x"2f58",x"3065",x"3ec5",x"36eb",x"3baa",x"3479",x"2b93",x"38f4",x"2f49"),
(x"2f0c",x"3ec2",x"3718",x"a3ae",x"ac2f",x"3bfb",x"3985",x"326e",x"2e32",x"3eb9",x"3714",x"a745",x"ad9b",x"3bf7",x"397d",x"3257",x"2e77",x"3ec4",x"3717",x"a984",x"a0c2",x"3bfd",x"3980",x"3272"),
(x"2e32",x"3eb9",x"3714",x"a745",x"ad9b",x"3bf7",x"397d",x"3257",x"2f0c",x"3ec2",x"3718",x"a3ae",x"ac2f",x"3bfb",x"3985",x"326e",x"3072",x"3eb8",x"3715",x"2081",x"ad9e",x"3bf8",x"3996",x"3257"),
(x"301e",x"3ec3",x"3718",x"224c",x"a36c",x"3bff",x"3990",x"326f",x"3056",x"3ec4",x"3718",x"26a1",x"97c8",x"3bff",x"3994",x"3272",x"3072",x"3eb8",x"3715",x"2081",x"ad9e",x"3bf8",x"3996",x"3257"),
(x"2fff",x"3eed",x"3716",x"baa5",x"b86c",x"2baa",x"390c",x"2e3b",x"2fff",x"3eec",x"36ee",x"bb1d",x"b747",x"2911",x"390e",x"2dec",x"2fc2",x"3eef",x"3713",x"b46c",x"bbaf",x"a5f6",x"3908",x"2e32"),
(x"2e96",x"3ede",x"3717",x"bbff",x"2481",x"2487",x"38fa",x"3158",x"2e77",x"3ec4",x"3717",x"bbe8",x"30a2",x"2973",x"38f6",x"31c5",x"2e93",x"3ede",x"36eb",x"bbfd",x"212b",x"29e6",x"3905",x"3161"),
(x"2fc4",x"3ef0",x"36ee",x"b52c",x"bb8d",x"ac0b",x"3908",x"2de8",x"2f3e",x"3ef0",x"36ee",x"314a",x"bbe2",x"a87e",x"38ff",x"2de6",x"2fc2",x"3eef",x"3713",x"b46c",x"bbaf",x"a5f6",x"3908",x"2e32"),
(x"2f0c",x"3ec2",x"3718",x"3a6d",x"3838",x"3468",x"394f",x"2e2f",x"2f2a",x"3ec5",x"36eb",x"3a79",x"3840",x"3401",x"3949",x"2dd9",x"301e",x"3ec3",x"3718",x"b98b",x"396b",x"33db",x"393b",x"2e58"),
(x"2e24",x"3eb8",x"36eb",x"b6d0",x"bb39",x"2ab1",x"38fd",x"320b",x"2e32",x"3eb9",x"3714",x"af03",x"bbf3",x"23ef",x"38f4",x"31ff",x"3079",x"3eb9",x"36eb",x"3409",x"bbbc",x"27e2",x"38ee",x"32c0"),
(x"2eed",x"3ee8",x"3716",x"3ba1",x"34a7",x"2cd8",x"38f4",x"2e32",x"2efa",x"3ee8",x"36ee",x"3b84",x"3534",x"2e9f",x"38f5",x"2de3",x"2f16",x"3ee4",x"3716",x"3bb3",x"33ed",x"2eeb",x"38ef",x"2e30"),
(x"3007",x"3fc7",x"3715",x"ad56",x"20d0",x"3bf8",x"3b8e",x"3bac",x"2f10",x"3fcc",x"370e",x"afd2",x"2717",x"3bef",x"3b82",x"3baf",x"2fbb",x"3fd4",x"3716",x"b0f9",x"a8af",x"3be5",x"3b89",x"3bb7"),
(x"3007",x"3fc7",x"3715",x"3bc5",x"2b9a",x"3358",x"3b5c",x"3886",x"2fbb",x"3fd4",x"3716",x"3add",x"375a",x"334d",x"3b5c",x"388d",x"301b",x"3fc7",x"36eb",x"3b99",x"3315",x"330d",x"3b61",x"3885"),
(x"301b",x"3f85",x"3713",x"291b",x"2b55",x"3bfb",x"3b94",x"3b76",x"2fb0",x"3f87",x"3714",x"2c39",x"29a5",x"3bf9",x"3b8e",x"3b77",x"3001",x"3f8f",x"3712",x"2a69",x"287e",x"3bfc",x"3b91",x"3b7e"),
(x"303e",x"3f87",x"3712",x"2a73",x"2a97",x"3bfa",x"3b97",x"3b78",x"3017",x"3f91",x"3711",x"2994",x"2977",x"3bfc",x"3b93",x"3b80",x"304c",x"3f8d",x"3711",x"2481",x"254c",x"3bff",x"3b98",x"3b7c"),
(x"3017",x"3f91",x"3711",x"2994",x"2977",x"3bfc",x"3b93",x"3b80",x"303e",x"3f87",x"3712",x"2a73",x"2a97",x"3bfa",x"3b97",x"3b78",x"3001",x"3f8f",x"3712",x"2a69",x"287e",x"3bfc",x"3b91",x"3b7e"),
(x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70",x"2ff2",x"3f82",x"3718",x"2e36",x"a160",x"3bf6",x"3b91",x"3b74",x"302f",x"3f81",x"3711",x"2fec",x"ac2c",x"3beb",x"3b96",x"3b73"),
(x"3040",x"3f6b",x"370f",x"1df0",x"a631",x"3bff",x"3b99",x"3b61",x"301b",x"3f6a",x"3713",x"2e9a",x"3366",x"3bbd",x"3b96",x"3b5f",x"2ff4",x"3f71",x"370e",x"a6d5",x"25c2",x"3bfe",x"3b92",x"3b65"),
(x"2ff4",x"3f71",x"370e",x"a6d5",x"25c2",x"3bfe",x"3b92",x"3b65",x"3013",x"3f76",x"3713",x"2538",x"ac79",x"3bfa",x"3b94",x"3b69",x"3040",x"3f6b",x"370f",x"1df0",x"a631",x"3bff",x"3b99",x"3b61"),
(x"305c",x"3f70",x"370f",x"2cd8",x"a71d",x"3bf9",x"3b9c",x"3b65",x"3013",x"3f76",x"3713",x"2538",x"ac79",x"3bfa",x"3b94",x"3b69",x"3058",x"3f79",x"370f",x"2ec5",x"19f0",x"3bf4",x"3b9b",x"3b6d"),
(x"302f",x"3f81",x"3711",x"2fec",x"ac2c",x"3beb",x"3b96",x"3b73",x"3014",x"3f78",x"3713",x"27e9",x"284d",x"3bfd",x"3b94",x"3b6b",x"3000",x"3f7a",x"3710",x"2c5b",x"b0a4",x"3be5",x"3b92",x"3b6d"),
(x"2fd7",x"3f4b",x"3712",x"2f67",x"a981",x"3bf0",x"3b90",x"3b46",x"2f48",x"3f4b",x"3715",x"26c2",x"ac63",x"3bfa",x"3b89",x"3b45",x"2f7f",x"3f52",x"3717",x"2ff2",x"aa7d",x"3bed",x"3b8c",x"3b4c"),
(x"3044",x"3f51",x"3714",x"9553",x"ab62",x"3bfc",x"3b98",x"3b4b",x"302b",x"3f5b",x"3716",x"2cd8",x"a7e2",x"3bf9",x"3b96",x"3b53",x"3050",x"3f55",x"3712",x"3163",x"a345",x"3be2",x"3b99",x"3b4e"),
(x"302b",x"3f5b",x"3716",x"2cd8",x"a7e2",x"3bf9",x"3b96",x"3b53",x"3044",x"3f51",x"3714",x"9553",x"ab62",x"3bfc",x"3b98",x"3b4b",x"300a",x"3f5a",x"3716",x"a818",x"ad04",x"3bf8",x"3b93",x"3b52"),
(x"3000",x"3f4e",x"3711",x"a40b",x"ad5c",x"3bf8",x"3b92",x"3b48",x"2fd3",x"3f57",x"3714",x"2504",x"ada9",x"3bf7",x"3b90",x"3b50",x"300a",x"3f5a",x"3716",x"a818",x"ad04",x"3bf8",x"3b93",x"3b52"),
(x"2fa9",x"3f54",x"3714",x"3036",x"a73e",x"3bed",x"3b8e",x"3b4d",x"3000",x"3f4e",x"3711",x"a40b",x"ad5c",x"3bf8",x"3b92",x"3b48",x"2fe3",x"3f4c",x"3711",x"327d",x"175f",x"3bd5",x"3b90",x"3b47"),
(x"302e",x"3f34",x"3711",x"3115",x"27d5",x"3be4",x"3b97",x"3b33",x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"2fe6",x"3f45",x"3712",x"3146",x"2c91",x"3bde",x"3b91",x"3b41"),
(x"2ef4",x"3f39",x"3719",x"23bb",x"27ae",x"3bfe",x"3b85",x"3b37",x"2f3d",x"3f39",x"3718",x"a138",x"ae95",x"3bf4",x"3b89",x"3b37",x"2ef3",x"3f38",x"3719",x"290e",x"af00",x"3bf2",x"3b85",x"3b37"),
(x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"2f4b",x"3f34",x"3715",x"a8bf",x"afdb",x"3bef",x"3b8a",x"3b33",x"2f3d",x"3f39",x"3718",x"a138",x"ae95",x"3bf4",x"3b89",x"3b37"),
(x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"2f3d",x"3f39",x"3718",x"a138",x"ae95",x"3bf4",x"3b89",x"3b37",x"2f49",x"3f3a",x"3718",x"ab4f",x"2525",x"3bfc",x"3b89",x"3b38"),
(x"2f1d",x"3f49",x"3717",x"ad2d",x"2ecb",x"3bed",x"3b87",x"3b44",x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2ede",x"3f43",x"3718",x"acf2",x"18ea",x"3bf9",x"3b84",x"3b3f"),
(x"2ede",x"3f43",x"3718",x"acf2",x"18ea",x"3bf9",x"3b84",x"3b3f",x"2ed4",x"3f47",x"3712",x"b59c",x"336a",x"3b42",x"3b83",x"3b42",x"2f1d",x"3f49",x"3717",x"ad2d",x"2ecb",x"3bed",x"3b87",x"3b44"),
(x"2fe6",x"3f45",x"3712",x"3146",x"2c91",x"3bde",x"3b91",x"3b41",x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2f3a",x"3f49",x"3716",x"300a",x"2da8",x"3be7",x"3b89",x"3b44"),
(x"2f48",x"3f4b",x"3715",x"26c2",x"ac63",x"3bfa",x"3b89",x"3b45",x"2fd7",x"3f4b",x"3712",x"2f67",x"a981",x"3bf0",x"3b90",x"3b46",x"2f3a",x"3f49",x"3716",x"300a",x"2da8",x"3be7",x"3b89",x"3b44"),
(x"2f5a",x"3f53",x"3717",x"17c8",x"9f79",x"3c00",x"3b8a",x"3b4d",x"2f48",x"3f4b",x"3715",x"26c2",x"ac63",x"3bfa",x"3b89",x"3b45",x"2f3c",x"3f4d",x"3714",x"257a",x"ae8a",x"3bf4",x"3b89",x"3b47"),
(x"2ece",x"3f60",x"3714",x"adba",x"2266",x"3bf7",x"3b83",x"3b57",x"2f11",x"3f58",x"3715",x"251e",x"2d06",x"3bf9",x"3b86",x"3b51",x"2e9f",x"3f5d",x"3714",x"975f",x"2c2c",x"3bfb",x"3b81",x"3b54"),
(x"2ec2",x"3f6b",x"3715",x"b468",x"247a",x"3bb0",x"3b83",x"3b60",x"2ece",x"3f60",x"3714",x"adba",x"2266",x"3bf7",x"3b83",x"3b57",x"2e7c",x"3f69",x"3712",x"b106",x"273e",x"3be5",x"3b80",x"3b5f"),
(x"2ed8",x"3f73",x"3717",x"b273",x"2f43",x"3bc8",x"3b84",x"3b66",x"2ec2",x"3f6b",x"3715",x"b468",x"247a",x"3bb0",x"3b83",x"3b60",x"2ea0",x"3f75",x"3710",x"b550",x"2e33",x"3b81",x"3b81",x"3b68"),
(x"2f3c",x"3f7a",x"3711",x"2e24",x"2a2b",x"3bf4",x"3b89",x"3b6c",x"2ed8",x"3f73",x"3717",x"b273",x"2f43",x"3bc8",x"3b84",x"3b66",x"2ef8",x"3f7d",x"3712",x"ab5c",x"2345",x"3bfc",x"3b85",x"3b6e"),
(x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70",x"2fc1",x"3f7b",x"3713",x"a5b5",x"b7de",x"3af6",x"3b8f",x"3b6e",x"2f7e",x"3f7b",x"3712",x"add2",x"b04b",x"3be4",x"3b8c",x"3b6d"),
(x"2fc5",x"3f84",x"3716",x"2553",x"32c7",x"3bd1",x"3b8f",x"3b75",x"2ff2",x"3f82",x"3718",x"2e36",x"a160",x"3bf6",x"3b91",x"3b74",x"2fad",x"3f83",x"3716",x"af4b",x"aa5f",x"3bf0",x"3b8e",x"3b74"),
(x"300c",x"3f84",x"3716",x"2f15",x"329c",x"3bc6",x"3b93",x"3b75",x"2ff2",x"3f82",x"3718",x"2e36",x"a160",x"3bf6",x"3b91",x"3b74",x"2fc5",x"3f84",x"3716",x"2553",x"32c7",x"3bd1",x"3b8f",x"3b75"),
(x"2f8e",x"3f93",x"370f",x"2edc",x"2cd0",x"3bee",x"3b8c",x"3b81",x"2fe3",x"3f8f",x"3713",x"2da3",x"2f15",x"3beb",x"3b90",x"3b7e",x"2f3b",x"3f8e",x"3717",x"30e7",x"3057",x"3bd4",x"3b88",x"3b7d"),
(x"2f5a",x"3f9e",x"3716",x"2adf",x"a6b5",x"3bfc",x"3b89",x"3b8a",x"2f8e",x"3f93",x"370f",x"2edc",x"2cd0",x"3bee",x"3b8c",x"3b81",x"2eeb",x"3f9c",x"3713",x"29b8",x"a6e2",x"3bfd",x"3b83",x"3b88"),
(x"2f5a",x"3f9e",x"3716",x"2adf",x"a6b5",x"3bfc",x"3b89",x"3b8a",x"2eeb",x"3f9c",x"3713",x"29b8",x"a6e2",x"3bfd",x"3b83",x"3b88",x"2ee1",x"3faa",x"3717",x"2bf6",x"25ae",x"3bfb",x"3b82",x"3b93"),
(x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1",x"2ee1",x"3faa",x"3717",x"2bf6",x"25ae",x"3bfb",x"3b82",x"3b93",x"2ebe",x"3fb5",x"370f",x"b6c9",x"2fac",x"3b2e",x"3b7f",x"3b9c"),
(x"2ebe",x"3fb5",x"370f",x"b6c9",x"2fac",x"3b2e",x"3b7f",x"3b9c",x"2ecd",x"3fb8",x"370d",x"b809",x"2e09",x"3add",x"3b80",x"3b9f",x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1"),
(x"2f10",x"3fcc",x"370e",x"afd2",x"2717",x"3bef",x"3b82",x"3baf",x"3007",x"3fc7",x"3715",x"ad56",x"20d0",x"3bf8",x"3b8e",x"3bac",x"2efa",x"3fc1",x"3712",x"a9f0",x"2b1d",x"3bfa",x"3b81",x"3ba6"),
(x"2ffb",x"3fba",x"3715",x"3b82",x"b440",x"330f",x"3b5b",x"387f",x"300f",x"3fb9",x"36eb",x"3b89",x"b473",x"31fc",x"3b60",x"387e",x"2f8b",x"3fa8",x"370e",x"3b5f",x"b5f1",x"2f4f",x"3b5a",x"3875"),
(x"302f",x"3f1a",x"3710",x"bbfd",x"a997",x"a09b",x"3b92",x"3a0f",x"302b",x"3f12",x"3714",x"bbeb",x"308b",x"98b5",x"3b92",x"3a0b",x"302e",x"3f14",x"36eb",x"bbf5",x"2e59",x"2467",x"3b8d",x"3a0c"),
(x"2ff3",x"3f30",x"3714",x"bb1c",x"b754",x"223f",x"3b92",x"3a1b",x"3024",x"3f23",x"3713",x"bba5",x"b497",x"ac28",x"3b92",x"3a14",x"3029",x"3f23",x"36eb",x"bba1",x"b4cc",x"1f45",x"3b8d",x"3a14"),
(x"3021",x"3f0e",x"3712",x"bb76",x"35c5",x"204d",x"3b92",x"3a09",x"300e",x"3f0b",x"3714",x"b95a",x"39f1",x"2032",x"3b92",x"3a07",x"301c",x"3f0c",x"36eb",x"bab1",x"3862",x"21f0",x"3b8d",x"3a08"),
(x"2fe4",x"3f08",x"3714",x"b5bf",x"3b76",x"27db",x"3b92",x"3a05",x"2fe9",x"3f08",x"36eb",x"b7e1",x"3af5",x"269a",x"3b8d",x"3a05",x"300e",x"3f0b",x"3714",x"b95a",x"39f1",x"2032",x"3b92",x"3a07"),
(x"2f7e",x"3f06",x"3715",x"2836",x"3bfd",x"294c",x"3b92",x"3a01",x"2f83",x"3f07",x"36eb",x"b03c",x"3beb",x"299e",x"3b8d",x"3a01",x"2fe4",x"3f08",x"3714",x"b5bf",x"3b76",x"27db",x"3b92",x"3a05"),
(x"2f19",x"3f08",x"3716",x"386f",x"3aa7",x"2604",x"3b92",x"39fe",x"2f1b",x"3f08",x"36eb",x"3868",x"3aab",x"296a",x"3b8d",x"39fe",x"2f7e",x"3f06",x"3715",x"2836",x"3bfd",x"294c",x"3b92",x"3a01"),
(x"2f19",x"3f08",x"3716",x"386f",x"3aa7",x"2604",x"3b92",x"39fe",x"2ec8",x"3f0e",x"3714",x"3b01",x"37b5",x"2839",x"3b92",x"39f9",x"2f1b",x"3f08",x"36eb",x"3868",x"3aab",x"296a",x"3b8d",x"39fe"),
(x"2eb5",x"3f13",x"3714",x"3be6",x"b10f",x"9bfc",x"3b92",x"39f6",x"2eb5",x"3f13",x"36eb",x"3bf9",x"2d11",x"2511",x"3b8d",x"39f7",x"2ec8",x"3f0e",x"3714",x"3b01",x"37b5",x"2839",x"3b92",x"39f9"),
(x"2ed5",x"3f18",x"3715",x"3928",x"ba1d",x"1553",x"3b92",x"39f4",x"2ecf",x"3f18",x"36eb",x"390c",x"ba34",x"2532",x"3b8d",x"39f4",x"2eb5",x"3f13",x"3714",x"3be6",x"b10f",x"9bfc",x"3b92",x"39f6"),
(x"2ed5",x"3f18",x"3715",x"3928",x"ba1d",x"1553",x"3b8d",x"364c",x"2f14",x"3f18",x"3714",x"afe2",x"bbee",x"28fd",x"3b8d",x"3650",x"2ecf",x"3f18",x"36eb",x"390c",x"ba34",x"2532",x"3b92",x"364a"),
(x"2f14",x"3f18",x"3714",x"afe2",x"bbee",x"28fd",x"3b8d",x"3650",x"2f4a",x"3f16",x"3711",x"b64f",x"bb52",x"2d1b",x"3b8e",x"3654",x"2f19",x"3f18",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3b92",x"364f"),
(x"2f99",x"3f25",x"3713",x"3bc2",x"33a4",x"298a",x"3b8e",x"366b",x"2f9f",x"3f25",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b93",x"366c",x"2faf",x"3f23",x"3711",x"3a7a",x"38af",x"283c",x"3b8e",x"3669"),
(x"2f4a",x"3f16",x"3711",x"b64f",x"bb52",x"2d1b",x"3b8e",x"3654",x"2f9c",x"3f16",x"3710",x"3416",x"bbad",x"2f8d",x"3b8f",x"365a",x"2f44",x"3f15",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3b93",x"3652"),
(x"301b",x"3f6a",x"3713",x"b583",x"bb63",x"3153",x"3b46",x"384c",x"3013",x"3f68",x"36eb",x"b5e4",x"bb4d",x"31a2",x"3b48",x"3847",x"2ff0",x"3f6f",x"370f",x"ba9c",x"b854",x"30fa",x"3b44",x"384a"),
(x"2ffb",x"3fba",x"3715",x"3b82",x"b440",x"330f",x"3b5b",x"387f",x"3007",x"3fc7",x"3715",x"3bc5",x"2b9a",x"3358",x"3b5c",x"3886",x"300f",x"3fb9",x"36eb",x"3b89",x"b473",x"31fc",x"3b60",x"387e"),
(x"2faf",x"3f23",x"3711",x"340b",x"26c2",x"3bbc",x"3b8f",x"3b25",x"2fd1",x"3f20",x"3710",x"2856",x"a9ab",x"3bfc",x"3b90",x"3b23",x"2f3e",x"3f25",x"3718",x"2b65",x"b528",x"3b8f",x"3b89",x"3b27"),
(x"2f14",x"3fbc",x"3715",x"bbd7",x"b1f9",x"2c2a",x"3b55",x"389b",x"2f10",x"3fba",x"3716",x"b8de",x"3a57",x"297d",x"3b55",x"389c",x"2f0d",x"3fbb",x"36eb",x"bbe3",x"2ce7",x"30c3",x"3b59",x"389f"),
(x"2ef8",x"3f7d",x"3712",x"b84e",x"3ab0",x"2ec7",x"3b26",x"3b1d",x"2ea0",x"3f75",x"3710",x"bb6a",x"35bb",x"2efe",x"3b27",x"3b21",x"2ee2",x"3f7e",x"36eb",x"b958",x"39de",x"2fe4",x"3b2b",x"3b1c"),
(x"2fc4",x"3f19",x"3711",x"3a7e",x"b887",x"3089",x"3b8f",x"365d",x"2fd3",x"3f18",x"36eb",x"3aa4",x"b859",x"2fe5",x"3b93",x"365d",x"2f9c",x"3f16",x"3710",x"3416",x"bbad",x"2f8d",x"3b8f",x"365a"),
(x"2f55",x"3f28",x"3718",x"bbe6",x"309e",x"2baa",x"3b22",x"3b6a",x"2f4a",x"3f28",x"36eb",x"bbe6",x"308f",x"2c41",x"3b28",x"3b68",x"2f5a",x"3f31",x"3715",x"bbfa",x"a710",x"2c48",x"3b21",x"3b65"),
(x"2fc4",x"3f19",x"3711",x"3a7e",x"b887",x"3089",x"3b8f",x"365d",x"2fdc",x"3f1c",x"3710",x"3bcc",x"b228",x"2f2f",x"3b8f",x"3661",x"2fd3",x"3f18",x"36eb",x"3aa4",x"b859",x"2fe5",x"3b93",x"365d"),
(x"2ff0",x"3f6f",x"370f",x"ba9c",x"b854",x"30fa",x"3b44",x"384a",x"2fdc",x"3f6e",x"36eb",x"bb7d",x"b521",x"3095",x"3b45",x"3846",x"2ff4",x"3f71",x"370e",x"bb25",x"370e",x"2d6a",x"3b42",x"384a"),
(x"3044",x"3f51",x"3714",x"3972",x"b9bb",x"30de",x"39f5",x"3b7d",x"3048",x"3f4f",x"36eb",x"36fe",x"bb25",x"2ea4",x"39fa",x"3b7b",x"3000",x"3f4e",x"3711",x"34dc",x"bb97",x"2d61",x"39f4",x"3b78"),
(x"2faf",x"3f23",x"3711",x"3a7a",x"38af",x"283c",x"3b8e",x"3669",x"2fb1",x"3f23",x"36eb",x"39db",x"396c",x"2c1a",x"3b93",x"366a",x"2fd1",x"3f20",x"3710",x"3b2f",x"36d9",x"2e52",x"3b8f",x"3666"),
(x"2fad",x"3f83",x"3716",x"b7e9",x"3af1",x"2aa7",x"3b25",x"3b16",x"2ef8",x"3f7d",x"3712",x"b84e",x"3ab0",x"2ec7",x"3b26",x"3b1d",x"2fb4",x"3f84",x"36eb",x"b776",x"3b0b",x"2d41",x"3b2a",x"3b15"),
(x"2f4b",x"3f34",x"3715",x"b95d",x"b9e3",x"2de3",x"3b21",x"3b64",x"2f5a",x"3f31",x"3715",x"bbfa",x"a710",x"2c48",x"3b21",x"3b65",x"2f48",x"3f33",x"36eb",x"b9df",x"b964",x"2d28",x"3b26",x"3b63"),
(x"3013",x"3f76",x"3713",x"bb5b",x"3634",x"2c08",x"3b40",x"384a",x"2ff4",x"3f71",x"370e",x"bb25",x"370e",x"2d6a",x"3b42",x"384a",x"300f",x"3f76",x"36eb",x"bad3",x"3822",x"2c4d",x"3b41",x"3845"),
(x"2f5a",x"3f9e",x"3716",x"3bff",x"20a8",x"2138",x"3b57",x"3870",x"2f8b",x"3fa8",x"370e",x"3b5f",x"b5f1",x"2f4f",x"3b5a",x"3875",x"2f5b",x"3f9d",x"36eb",x"3bfe",x"1e8d",x"2828",x"3b5c",x"386e"),
(x"2fad",x"3f83",x"3716",x"b7e9",x"3af1",x"2aa7",x"3b25",x"3b16",x"2fb4",x"3f84",x"36eb",x"b776",x"3b0b",x"2d41",x"3b2a",x"3b15",x"2fc5",x"3f84",x"3716",x"bbde",x"31b5",x"2825",x"3b25",x"3b15"),
(x"2ef3",x"3f38",x"3719",x"b9a6",x"b994",x"2faf",x"3b1f",x"3b60",x"2f4b",x"3f34",x"3715",x"b95d",x"b9e3",x"2de3",x"3b21",x"3b64",x"2ed5",x"3f38",x"36eb",x"b9ed",x"b94b",x"2f45",x"3b25",x"3b5e"),
(x"2fe3",x"3f4c",x"3711",x"3b12",x"b762",x"2ca3",x"3b1e",x"3bb2",x"3000",x"3f4e",x"3711",x"34dc",x"bb97",x"2d61",x"3b1e",x"3bb3",x"2ff6",x"3f4d",x"36eb",x"37d8",x"baf6",x"2a35",x"3b23",x"3bb4"),
(x"3014",x"3f78",x"3713",x"bb09",x"b791",x"2ab8",x"3b3f",x"3849",x"3013",x"3f76",x"3713",x"bb5b",x"3634",x"2c08",x"3b40",x"384a",x"3010",x"3f77",x"36eb",x"b9e9",x"b955",x"2e31",x"3b40",x"3844"),
(x"2f5a",x"3f9e",x"3716",x"3bff",x"20a8",x"2138",x"3b57",x"3870",x"2f5b",x"3f9d",x"36eb",x"3bfe",x"1e8d",x"2828",x"3b5c",x"386e",x"2f8e",x"3f93",x"370f",x"3ad7",x"3821",x"29e3",x"3b57",x"386a"),
(x"2fc5",x"3f84",x"3716",x"bbde",x"31b5",x"2825",x"3b3f",x"38b1",x"2fc0",x"3f84",x"36eb",x"bb23",x"b71d",x"2cde",x"3b42",x"38b6",x"2fb0",x"3f87",x"3714",x"b9e8",x"b951",x"2f27",x"3b40",x"38b0"),
(x"2ef3",x"3f38",x"3719",x"b9a6",x"b994",x"2faf",x"3b1f",x"3b60",x"2ed5",x"3f38",x"36eb",x"b9ed",x"b94b",x"2f45",x"3b25",x"3b5e",x"2ef4",x"3f39",x"3719",x"b251",x"3bca",x"2f22",x"3b1f",x"3b60"),
(x"2fd7",x"3f4b",x"3712",x"3bf7",x"283f",x"2d8f",x"3b1e",x"3bb1",x"2fe5",x"3f4a",x"36eb",x"3bf8",x"a379",x"2d44",x"3b23",x"3bb2",x"2fe6",x"3f45",x"3712",x"3b92",x"3509",x"2cb4",x"3b1f",x"3bae"),
(x"3000",x"3f7a",x"3710",x"b833",x"bac7",x"2d1d",x"39f6",x"3bab",x"3014",x"3f78",x"3713",x"bb09",x"b791",x"2ab8",x"39f6",x"3bad",x"3010",x"3f77",x"36eb",x"b9e9",x"b955",x"2e31",x"39fb",x"3bac"),
(x"2fe3",x"3f8f",x"3713",x"37c3",x"3af3",x"2e28",x"3b56",x"3866",x"2f8e",x"3f93",x"370f",x"3ad7",x"3821",x"29e3",x"3b57",x"386a",x"2fee",x"3f8f",x"36eb",x"373f",x"3b1a",x"2d3c",x"3b5b",x"3865"),
(x"2fb0",x"3f87",x"3714",x"b9e8",x"b951",x"2f27",x"3b40",x"38b0",x"2f9f",x"3f86",x"36eb",x"b97a",x"b9b6",x"3099",x"3b43",x"38b5",x"2f3b",x"3f8e",x"3717",x"ba77",x"b889",x"310c",x"3b44",x"38ad"),
(x"2f3d",x"3f39",x"3718",x"b0c5",x"3be6",x"2ad9",x"3b1e",x"3b5e",x"2ef4",x"3f39",x"3719",x"b251",x"3bca",x"2f22",x"3b1f",x"3b60",x"2f48",x"3f3a",x"36eb",x"bb01",x"3745",x"3141",x"3b22",x"3b5a"),
(x"2fe6",x"3f45",x"3712",x"3b92",x"3509",x"2cb4",x"3b1f",x"3bae",x"2fee",x"3f46",x"36eb",x"3b57",x"3625",x"2e99",x"3b24",x"3bb0",x"302e",x"3f34",x"3711",x"3b70",x"3585",x"3014",x"3b22",x"3ba5"),
(x"2f7e",x"3f7b",x"3712",x"32e8",x"bbcb",x"2c10",x"39f5",x"3ba7",x"2fc1",x"3f7b",x"3713",x"b0a8",x"bbea",x"22cf",x"39f5",x"3ba9",x"2fb8",x"3f7b",x"36eb",x"b046",x"bbe8",x"2cb7",x"39fa",x"3ba8"),
(x"2fe3",x"3f8f",x"3713",x"37c3",x"3af3",x"2e28",x"3b56",x"3866",x"2fee",x"3f8f",x"36eb",x"373f",x"3b1a",x"2d3c",x"3b5b",x"3865",x"3001",x"3f8f",x"3712",x"b721",x"3b24",x"2bf2",x"3b56",x"3865"),
(x"2f3b",x"3f8e",x"3717",x"ba77",x"b889",x"310c",x"3b44",x"38ad",x"2f20",x"3f8e",x"36eb",x"baff",x"b73c",x"3197",x"3b47",x"38b2",x"2eeb",x"3f9c",x"3713",x"bbc6",x"b1be",x"30de",x"3b4a",x"38a9"),
(x"302e",x"3f34",x"3711",x"3b70",x"3585",x"3014",x"3b22",x"3ba5",x"303d",x"3f33",x"36eb",x"3b99",x"345f",x"30d6",x"3b27",x"3ba6",x"3046",x"3f24",x"3711",x"3be4",x"2d1d",x"308b",x"3b24",x"3b9d"),
(x"2ed8",x"3f73",x"3717",x"3b6f",x"b5e5",x"261e",x"39f4",x"3ba0",x"2f3c",x"3f7a",x"3711",x"3934",x"ba0d",x"2c18",x"39f5",x"3ba5",x"2ede",x"3f73",x"36eb",x"3aaf",x"b860",x"2a70",x"39fa",x"3ba0"),
(x"3001",x"3f8f",x"3712",x"b721",x"3b24",x"2bf2",x"3b56",x"3865",x"3004",x"3f90",x"36eb",x"b8ae",x"3a73",x"2d47",x"3b5b",x"3864",x"3017",x"3f91",x"3711",x"b5dd",x"3b65",x"2eae",x"3b56",x"3864"),
(x"2ee1",x"3faa",x"3717",x"bbf0",x"af10",x"2aec",x"3b4e",x"38a3",x"2eeb",x"3f9c",x"3713",x"bbc6",x"b1be",x"30de",x"3b4a",x"38a9",x"2ed7",x"3fa9",x"36eb",x"bbea",x"ae0a",x"2f12",x"3b52",x"38a8"),
(x"2f49",x"3f3a",x"3718",x"baf6",x"b7e0",x"2460",x"3b25",x"3b46",x"2f3d",x"3f39",x"3718",x"b0c5",x"3be6",x"2ad9",x"3b25",x"3b47",x"2f48",x"3f3a",x"36eb",x"bb01",x"3745",x"3141",x"3b2a",x"3b47"),
(x"3046",x"3f13",x"3714",x"3bec",x"ad02",x"2f52",x"3b26",x"3b94",x"3046",x"3f24",x"3711",x"3be4",x"2d1d",x"308b",x"3b24",x"3b9d",x"304f",x"3f13",x"36eb",x"3be8",x"ad66",x"3010",x"3b2b",x"3b95"),
(x"2ec2",x"3f6b",x"3715",x"3bfe",x"2412",x"286a",x"39f5",x"3b9b",x"2ed8",x"3f73",x"3717",x"3b6f",x"b5e5",x"261e",x"39f4",x"3ba0",x"2ec6",x"3f6b",x"36eb",x"3bfa",x"ac62",x"2617",x"39fa",x"3b9c"),
(x"3017",x"3f91",x"3711",x"b5dd",x"3b65",x"2eae",x"3b56",x"3864",x"3014",x"3f92",x"36eb",x"ae29",x"3be6",x"3005",x"3b5b",x"3863",x"3038",x"3f91",x"3712",x"35a5",x"3b63",x"30cc",x"3b55",x"3861"),
(x"2ee1",x"3faa",x"3717",x"bbf0",x"af10",x"2aec",x"3b4e",x"38a3",x"2ed7",x"3fa9",x"36eb",x"bbea",x"ae0a",x"2f12",x"3b52",x"38a8",x"2ebe",x"3fb5",x"370f",x"bbdd",x"b0de",x"2e6c",x"3b53",x"38a0"),
(x"2f16",x"3f3e",x"3715",x"b9d1",x"b974",x"2cc6",x"3b26",x"3b44",x"2ef5",x"3f3e",x"36eb",x"ba0e",x"b929",x"2e78",x"3b2b",x"3b44",x"2ede",x"3f43",x"3718",x"bb13",x"b732",x"2fec",x"3b26",x"3b41"),
(x"3046",x"3f13",x"3714",x"3bec",x"ad02",x"2f52",x"3b26",x"3b94",x"304f",x"3f13",x"36eb",x"3be8",x"ad66",x"3010",x"3b2b",x"3b95",x"3036",x"3f0b",x"3712",x"3b45",x"b640",x"30a6",x"3b27",x"3b90"),
(x"2fdc",x"3f1c",x"3710",x"3bcc",x"b228",x"2f2f",x"3b8f",x"3661",x"2fd1",x"3f20",x"3710",x"3b2f",x"36d9",x"2e52",x"3b8f",x"3666",x"2fec",x"3f1c",x"36eb",x"3bf4",x"9edc",x"2eb6",x"3b93",x"3662"),
(x"2ece",x"3f60",x"3714",x"3b81",x"3558",x"2da6",x"39f5",x"3b96",x"2ec2",x"3f6b",x"3715",x"3bfe",x"2412",x"286a",x"39f5",x"3b9b",x"2ed7",x"3f61",x"36eb",x"3bcf",x"32aa",x"2bc8",x"39fa",x"3b96"),
(x"3038",x"3f91",x"3712",x"35a5",x"3b63",x"30cc",x"3b55",x"3861",x"3043",x"3f92",x"36eb",x"3913",x"3a0d",x"310f",x"3b5a",x"3860",x"304c",x"3f8d",x"3711",x"3bb2",x"332f",x"30f4",x"3b55",x"385f"),
(x"2ebe",x"3fb5",x"370f",x"bbdd",x"b0de",x"2e6c",x"3b53",x"38a0",x"2eaa",x"3fb4",x"36eb",x"bbe4",x"aadf",x"30ee",x"3b56",x"38a4",x"2ecd",x"3fb8",x"370d",x"bb0d",x"370c",x"3168",x"3b54",x"389f"),
(x"2ede",x"3f43",x"3718",x"bb13",x"b732",x"2fec",x"3b26",x"3b41",x"2ec6",x"3f43",x"36eb",x"bbbf",x"b333",x"2ed2",x"3b2b",x"3b41",x"2ed4",x"3f47",x"3712",x"bbf0",x"2c20",x"2e95",x"3b27",x"3b3e"),
(x"3036",x"3f0b",x"3712",x"3b45",x"b640",x"30a6",x"3b27",x"3b90",x"303e",x"3f0a",x"36eb",x"3ab2",x"b834",x"30cf",x"3b2c",x"3b91",x"3003",x"3f04",x"3715",x"393c",x"b9e9",x"311d",x"3b27",x"3b8b"),
(x"2f11",x"3f58",x"3715",x"3a65",x"38c0",x"2d9c",x"39f5",x"3b91",x"2ece",x"3f60",x"3714",x"3b81",x"3558",x"2da6",x"39f5",x"3b96",x"2f1f",x"3f59",x"36eb",x"3ac2",x"3833",x"2e85",x"39fa",x"3b91"),
(x"304c",x"3f8d",x"3711",x"3bb2",x"332f",x"30f4",x"3b55",x"385f",x"3057",x"3f8d",x"36eb",x"3be5",x"adbc",x"3036",x"3b59",x"385d",x"303e",x"3f87",x"3712",x"3ae4",x"b7c3",x"30c9",x"3b53",x"385c"),
(x"2ee7",x"3fba",x"3713",x"b451",x"3bac",x"2d81",x"3b54",x"389d",x"2ecd",x"3fb8",x"370d",x"bb0d",x"370c",x"3168",x"3b54",x"389f",x"2ee1",x"3fbb",x"36eb",x"b571",x"3b6d",x"30cc",x"3b59",x"38a0"),
(x"2ed4",x"3f47",x"3712",x"bbf0",x"2c20",x"2e95",x"3b27",x"3b3e",x"2ecb",x"3f48",x"36eb",x"bbbf",x"3371",x"2dad",x"3b2b",x"3b3e",x"2ee4",x"3f49",x"3712",x"b297",x"3bcc",x"2d84",x"3b26",x"3b3d"),
(x"3003",x"3f04",x"3715",x"393c",x"b9e9",x"311d",x"3b27",x"3b8b",x"3007",x"3f02",x"36eb",x"37cb",x"bae6",x"3068",x"3b2c",x"3b8b",x"2f91",x"3f01",x"3715",x"1ef6",x"bbee",x"302a",x"3b27",x"3b87"),
(x"2f5a",x"3f53",x"3717",x"3939",x"3a0b",x"29e0",x"39f5",x"3b8e",x"2f11",x"3f58",x"3715",x"3a65",x"38c0",x"2d9c",x"39f5",x"3b91",x"2f61",x"3f54",x"36eb",x"39cd",x"3979",x"2caa",x"39fa",x"3b8e"),
(x"303e",x"3f87",x"3712",x"3ae4",x"b7c3",x"30c9",x"3b53",x"385c",x"3044",x"3f85",x"36eb",x"3902",x"ba23",x"306a",x"3b57",x"3859",x"301b",x"3f85",x"3713",x"3607",x"bb5e",x"2e4d",x"3b52",x"385a"),
(x"2f10",x"3fba",x"3716",x"b8de",x"3a57",x"297d",x"3b55",x"389c",x"2ee7",x"3fba",x"3713",x"b451",x"3bac",x"2d81",x"3b54",x"389d",x"2f0d",x"3fbb",x"36eb",x"bbe3",x"2ce7",x"30c3",x"3b59",x"389f"),
(x"2f1d",x"3f49",x"3717",x"aa07",x"3bfc",x"284d",x"3b26",x"3b3c",x"2ee4",x"3f49",x"3712",x"b297",x"3bcc",x"2d84",x"3b26",x"3b3d",x"2f24",x"3f49",x"36eb",x"ac56",x"3bf7",x"2bc1",x"3b2b",x"3b3b"),
(x"2f0e",x"3f04",x"3713",x"b82e",x"baba",x"306c",x"3b28",x"3b82",x"2f91",x"3f01",x"3715",x"1ef6",x"bbee",x"302a",x"3b27",x"3b87",x"2f13",x"3f02",x"36eb",x"b66a",x"bb44",x"2f81",x"3b2d",x"3b83"),
(x"2f7f",x"3f52",x"3717",x"ac93",x"3bf9",x"2918",x"39f5",x"3b8c",x"2f5a",x"3f53",x"3717",x"3939",x"3a0b",x"29e0",x"39f5",x"3b8e",x"2f7e",x"3f52",x"36eb",x"b5a6",x"3b74",x"2d53",x"39fa",x"3b8d"),
(x"300c",x"3f84",x"3716",x"3ac7",x"383c",x"283f",x"3b51",x"385a",x"301b",x"3f85",x"3713",x"3607",x"bb5e",x"2e4d",x"3b52",x"385a",x"300f",x"3f84",x"36eb",x"394d",x"39f2",x"2dc5",x"3b55",x"3856"),
(x"2f8b",x"3fa8",x"370e",x"3004",x"a71d",x"3bef",x"3b8a",x"3b93",x"2f5a",x"3f9e",x"3716",x"2adf",x"a6b5",x"3bfc",x"3b89",x"3b8a",x"2ee1",x"3faa",x"3717",x"2bf6",x"25ae",x"3bfb",x"3b82",x"3b93"),
(x"2f1d",x"3f49",x"3717",x"aa07",x"3bfc",x"284d",x"3b26",x"3b3c",x"2f24",x"3f49",x"36eb",x"ac56",x"3bf7",x"2bc1",x"3b2b",x"3b3b",x"2f3a",x"3f49",x"3716",x"b8f4",x"3a42",x"2c09",x"3b26",x"3b3b"),
(x"2e95",x"3f0a",x"3715",x"bae0",x"b7cf",x"30d4",x"3b27",x"3b7d",x"2f0e",x"3f04",x"3713",x"b82e",x"baba",x"306c",x"3b28",x"3b82",x"2e80",x"3f09",x"36eb",x"b9f2",x"b938",x"30b5",x"3b2c",x"3b7d"),
(x"2fa9",x"3f54",x"3714",x"b9a7",x"399f",x"2d1e",x"39f5",x"3b8a",x"2f7f",x"3f52",x"3717",x"ac93",x"3bf9",x"2918",x"39f5",x"3b8c",x"2f7e",x"3f52",x"36eb",x"b5a6",x"3b74",x"2d53",x"39fa",x"3b8d"),
(x"300c",x"3f84",x"3716",x"3ac7",x"383c",x"283f",x"3b51",x"385a",x"300f",x"3f84",x"36eb",x"394d",x"39f2",x"2dc5",x"3b55",x"3856",x"302f",x"3f81",x"3711",x"38c8",x"3a4e",x"30a8",x"3b50",x"3857"),
(x"2f3a",x"3f49",x"3716",x"b8f4",x"3a42",x"2c09",x"3b26",x"3b3b",x"2f37",x"3f4a",x"36eb",x"bb71",x"b58a",x"2fc3",x"3b2b",x"3b3a",x"2f48",x"3f4b",x"3715",x"bac2",x"b812",x"3146",x"3b26",x"3b3a"),
(x"2e5f",x"3f13",x"3715",x"bbec",x"abe2",x"2fce",x"3b27",x"3b78",x"2e95",x"3f0a",x"3715",x"bae0",x"b7cf",x"30d4",x"3b27",x"3b7d",x"2e4e",x"3f12",x"36eb",x"bbc4",x"b27a",x"3012",x"3b2c",x"3b77"),
(x"2fd3",x"3f57",x"3714",x"b97e",x"39c5",x"2dbf",x"39f5",x"3b88",x"2fd6",x"3f58",x"36eb",x"b976",x"39cc",x"2dcc",x"39fb",x"3b88",x"300a",x"3f5a",x"3716",x"b7d5",x"3af0",x"2d8e",x"39f6",x"3b86"),
(x"302f",x"3f81",x"3711",x"38c8",x"3a4e",x"30a8",x"3b50",x"3857",x"303f",x"3f82",x"36eb",x"39ec",x"392b",x"31e4",x"3b54",x"3854",x"3058",x"3f79",x"370f",x"3b4b",x"35cc",x"3223",x"3b4e",x"3853"),
(x"2efa",x"3fc1",x"3712",x"bbcf",x"b081",x"3141",x"3b57",x"3899",x"2edb",x"3fc1",x"36eb",x"bbdb",x"1c67",x"320a",x"3b5b",x"389c",x"2f10",x"3fcc",x"370e",x"bb7b",x"34a9",x"3270",x"3b5a",x"3895"),
(x"2f3c",x"3f4d",x"3714",x"3879",x"347b",x"3a3d",x"3b25",x"3b38",x"2f48",x"3f4b",x"3715",x"bac2",x"b812",x"3146",x"3b26",x"3b3a",x"2f06",x"3f51",x"3718",x"bac6",x"b7dc",x"3286",x"3b26",x"3b36"),
(x"2e70",x"3f1b",x"3717",x"bb55",x"35fd",x"307e",x"3b25",x"3b74",x"2e5f",x"3f13",x"3715",x"bbec",x"abe2",x"2fce",x"3b27",x"3b78",x"2e58",x"3f1c",x"36eb",x"bb6e",x"3575",x"309f",x"3b2b",x"3b73"),
(x"2ff3",x"3f30",x"3714",x"305e",x"21a1",x"3bec",x"3b92",x"3b30",x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"302e",x"3f34",x"3711",x"3115",x"27d5",x"3be4",x"3b97",x"3b33"),
(x"300a",x"3f5a",x"3716",x"b7d5",x"3af0",x"2d8e",x"39f6",x"3b86",x"3008",x"3f5b",x"36eb",x"b53f",x"3b87",x"2d28",x"39fb",x"3b86",x"302b",x"3f5b",x"3716",x"2345",x"3bf7",x"2dcc",x"39f6",x"3b83"),
(x"3058",x"3f79",x"370f",x"3b4b",x"35cc",x"3223",x"3b4e",x"3853",x"3065",x"3f79",x"36eb",x"3bbc",x"3212",x"3175",x"3b51",x"3850",x"305c",x"3f70",x"370f",x"3bd3",x"af46",x"3182",x"3b4b",x"384f"),
(x"2f06",x"3f51",x"3718",x"bac6",x"b7dc",x"3286",x"3b26",x"3b36",x"2ed7",x"3f52",x"36eb",x"badb",x"b7e7",x"30ac",x"3b2b",x"3b35",x"2e9f",x"3f5d",x"3714",x"bb6b",x"b587",x"3096",x"3b26",x"3b2f"),
(x"2e70",x"3f1b",x"3717",x"bb55",x"35fd",x"307e",x"3b25",x"3b74",x"2e58",x"3f1c",x"36eb",x"bb6e",x"3575",x"309f",x"3b2b",x"3b73",x"2ec0",x"3f22",x"3711",x"b8a4",x"3a69",x"309a",x"3b25",x"3b6f"),
(x"302b",x"3f5b",x"3716",x"2345",x"3bf7",x"2dcc",x"39f6",x"3b83",x"302e",x"3f5c",x"36eb",x"33e5",x"3bb4",x"2ec2",x"39fb",x"3b84",x"3045",x"3f59",x"3714",x"3976",x"39c0",x"3024",x"39f6",x"3b81"),
(x"305c",x"3f70",x"370f",x"3bd3",x"af46",x"3182",x"3b4b",x"384f",x"3068",x"3f6f",x"36eb",x"3b61",x"b5a0",x"3119",x"3b4e",x"384c",x"3040",x"3f6b",x"370f",x"3891",x"ba72",x"30f5",x"3b48",x"384d"),
(x"2f10",x"3fcc",x"370e",x"bb7b",x"34a9",x"3270",x"3b5a",x"3895",x"2ef9",x"3fcd",x"36eb",x"bade",x"37ab",x"31d3",x"3b5e",x"3897",x"2f7a",x"3fd4",x"3712",x"b8b5",x"3a3e",x"32bd",x"3b5c",x"388f"),
(x"2e9f",x"3f5d",x"3714",x"bb6b",x"b587",x"3096",x"3b26",x"3b2f",x"2e89",x"3f5d",x"36eb",x"bbba",x"b376",x"2f14",x"3b2c",x"3b2e",x"2e7c",x"3f69",x"3712",x"bbf0",x"aa00",x"2f46",x"3b27",x"3b28"),
(x"2f3e",x"3f25",x"3718",x"b8ae",x"3a78",x"2b7c",x"3b23",x"3b6c",x"2ec0",x"3f22",x"3711",x"b8a4",x"3a69",x"309a",x"3b25",x"3b6f",x"2f34",x"3f26",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3b28",x"3b6a"),
(x"3045",x"3f59",x"3714",x"3976",x"39c0",x"3024",x"39f6",x"3b81",x"3050",x"3f5a",x"36eb",x"3acb",x"3812",x"3065",x"39fb",x"3b81",x"3050",x"3f55",x"3712",x"3be0",x"2e5e",x"30a3",x"39f6",x"3b7f"),
(x"301b",x"3f6a",x"3713",x"b583",x"bb63",x"3153",x"3b46",x"384c",x"3040",x"3f6b",x"370f",x"3891",x"ba72",x"30f5",x"3b48",x"384d",x"3013",x"3f68",x"36eb",x"b5e4",x"bb4d",x"31a2",x"3b48",x"3847"),
(x"2fbb",x"3fd4",x"3716",x"3add",x"375a",x"334d",x"3b5c",x"388d",x"2f7a",x"3fd4",x"3712",x"b8b5",x"3a3e",x"32bd",x"3b5c",x"388f",x"2fd0",x"3fd7",x"36eb",x"3996",x"395e",x"33ec",x"3b61",x"388e"),
(x"2e7c",x"3f69",x"3712",x"bbf0",x"aa00",x"2f46",x"3b27",x"3b28",x"2e6b",x"3f6a",x"36eb",x"bbef",x"2d0b",x"2e69",x"3b2c",x"3b27",x"2ea0",x"3f75",x"3710",x"bb6a",x"35bb",x"2efe",x"3b27",x"3b21"),
(x"2f55",x"3f28",x"3718",x"bbe6",x"309e",x"2baa",x"3b22",x"3b6a",x"2f3e",x"3f25",x"3718",x"b8ae",x"3a78",x"2b7c",x"3b23",x"3b6c",x"2f4a",x"3f28",x"36eb",x"bbe6",x"308f",x"2c41",x"3b28",x"3b68"),
(x"3050",x"3f55",x"3712",x"3be0",x"2e5e",x"30a3",x"39f6",x"3b7f",x"305c",x"3f54",x"36eb",x"3bcf",x"b173",x"3043",x"39fb",x"3b7e",x"3044",x"3f51",x"3714",x"3972",x"b9bb",x"30de",x"39f5",x"3b7d"),
(x"3046",x"3f24",x"3711",x"2cd1",x"250b",x"3bf9",x"3b99",x"3b27",x"3046",x"3f13",x"3714",x"aeb0",x"28fa",x"3bf3",x"3b9a",x"3b19",x"302f",x"3f1a",x"3710",x"a828",x"260a",x"3bfe",x"3b97",x"3b1e"),
(x"3036",x"3f0b",x"3712",x"2587",x"208e",x"3bff",x"3b98",x"3b12",x"300e",x"3f0b",x"3714",x"28bf",x"2c20",x"3bfa",x"3b95",x"3b11",x"3021",x"3f0e",x"3712",x"a953",x"27ae",x"3bfd",x"3b96",x"3b14"),
(x"3036",x"3f0b",x"3712",x"2587",x"208e",x"3bff",x"3b98",x"3b12",x"3003",x"3f04",x"3715",x"20ea",x"2afd",x"3bfc",x"3b94",x"3b0c",x"300e",x"3f0b",x"3714",x"28bf",x"2c20",x"3bfa",x"3b95",x"3b11"),
(x"3003",x"3f04",x"3715",x"20ea",x"2afd",x"3bfc",x"3b94",x"3b0c",x"2f91",x"3f01",x"3715",x"a7e2",x"29b2",x"3bfc",x"3b8e",x"3b09",x"2fe4",x"3f08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3b92",x"3b0f"),
(x"2f91",x"3f01",x"3715",x"a7e2",x"29b2",x"3bfc",x"3b8e",x"3b09",x"2f0e",x"3f04",x"3713",x"ab1d",x"aee4",x"3bf0",x"3b88",x"3b0b",x"2f7e",x"3f06",x"3715",x"a70a",x"a779",x"3bfe",x"3b8d",x"3b0d"),
(x"2f0e",x"3f04",x"3713",x"ab1d",x"aee4",x"3bf0",x"3b88",x"3b0b",x"2e95",x"3f0a",x"3715",x"2266",x"9d87",x"3bff",x"3b82",x"3b10",x"2f19",x"3f08",x"3716",x"a4bc",x"aceb",x"3bf9",x"3b89",x"3b0e"),
(x"2e95",x"3f0a",x"3715",x"2266",x"9d87",x"3bff",x"3b82",x"3b10",x"2e5f",x"3f13",x"3715",x"2891",x"a7ce",x"3bfd",x"3b7f",x"3b17",x"2ec8",x"3f0e",x"3714",x"28e0",x"299e",x"3bfc",x"3b85",x"3b13"),
(x"2eb5",x"3f13",x"3714",x"2538",x"a9ab",x"3bfd",x"3b83",x"3b18",x"2e5f",x"3f13",x"3715",x"2891",x"a7ce",x"3bfd",x"3b7f",x"3b17",x"2ed5",x"3f18",x"3715",x"2c67",x"28a5",x"3bf9",x"3b85",x"3b1b"),
(x"2e70",x"3f1b",x"3717",x"2d06",x"2793",x"3bf8",x"3b80",x"3b1e",x"2ec0",x"3f22",x"3711",x"28d9",x"a52b",x"3bfe",x"3b83",x"3b24",x"2ed5",x"3f18",x"3715",x"2c67",x"28a5",x"3bf9",x"3b85",x"3b1b"),
(x"2f14",x"3f18",x"3714",x"2a45",x"2b10",x"3bfa",x"3b88",x"3b1c",x"2fc4",x"3f19",x"3711",x"2bef",x"a8a8",x"3bfa",x"3b90",x"3b1d",x"2f4a",x"3f16",x"3711",x"2a66",x"b31a",x"3bca",x"3b8a",x"3b1a"),
(x"2f55",x"3f28",x"3718",x"3420",x"1418",x"3bba",x"3b8a",x"3b29",x"2f99",x"3f25",x"3713",x"341f",x"ac3c",x"3bb6",x"3b8d",x"3b26",x"2f3e",x"3f25",x"3718",x"2b65",x"b528",x"3b8f",x"3b89",x"3b27"),
(x"2f5a",x"3f31",x"3715",x"27ae",x"a4ea",x"3bfe",x"3b8a",x"3b31",x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"2f94",x"3f29",x"3714",x"2de0",x"a4c2",x"3bf6",x"3b8d",x"3b2a"),
(x"2fd1",x"3f20",x"3710",x"2856",x"a9ab",x"3bfc",x"3b90",x"3b23",x"2fc4",x"3f19",x"3711",x"2bef",x"a8a8",x"3bfa",x"3b90",x"3b1d",x"2f14",x"3f18",x"3714",x"2a45",x"2b10",x"3bfa",x"3b88",x"3b1c"),
(x"3056",x"3ec4",x"3718",x"26a1",x"97c8",x"3bff",x"3994",x"3272",x"301e",x"3ec3",x"3718",x"224c",x"a36c",x"3bff",x"3990",x"326f",x"3033",x"3ee0",x"3715",x"21a1",x"23fc",x"3bff",x"3991",x"32b4"),
(x"2f5a",x"3f31",x"3715",x"27ae",x"a4ea",x"3bfe",x"3b8a",x"3b31",x"2f4b",x"3f34",x"3715",x"a8bf",x"afdb",x"3bef",x"3b8a",x"3b33",x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34"),
(x"2f94",x"3f29",x"3714",x"3bf3",x"ae23",x"2b27",x"3b8e",x"3670",x"2fb5",x"3f36",x"3718",x"39e5",x"b968",x"0000",x"3b8d",x"367d",x"2fb5",x"3f36",x"36eb",x"346a",x"bb91",x"316a",x"3b92",x"367e"),
(x"2f13",x"3dea",x"3715",x"2d56",x"a0d0",x"3bf8",x"385b",x"38b5",x"3008",x"3de5",x"370e",x"2fd2",x"a717",x"3bef",x"386c",x"38b1",x"2f67",x"3ddc",x"3716",x"30f9",x"28af",x"3be5",x"3862",x"38a6"),
(x"2f13",x"3dea",x"3715",x"bbc5",x"ab9a",x"3358",x"3b13",x"3a3f",x"2f67",x"3ddc",x"3716",x"badd",x"b75a",x"334d",x"3b13",x"3a46",x"2eeb",x"3de9",x"36eb",x"bb99",x"b315",x"330d",x"3b18",x"3a3e"),
(x"2eea",x"3e2b",x"3713",x"a91b",x"ab55",x"3bfb",x"3852",x"38ff",x"2f72",x"3e29",x"3714",x"ac39",x"a9a5",x"3bf9",x"385b",x"38fe",x"2f20",x"3e21",x"3712",x"aa69",x"a87e",x"3bfc",x"3856",x"38f5"),
(x"2ea4",x"3e29",x"3712",x"aa73",x"aa97",x"3bfa",x"384e",x"38fd",x"2ef3",x"3e1f",x"3711",x"a994",x"a977",x"3bfc",x"3853",x"38f2",x"2e89",x"3e24",x"3711",x"a481",x"a546",x"3bff",x"384c",x"38f7"),
(x"2ef3",x"3e1f",x"3711",x"a994",x"a977",x"3bfc",x"3853",x"38f2",x"2ea4",x"3e29",x"3712",x"aa73",x"aa97",x"3bfa",x"384e",x"38fd",x"2f20",x"3e21",x"3712",x"aa69",x"a87e",x"3bfc",x"3856",x"38f5"),
(x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908",x"2f2f",x"3e2e",x"3718",x"ae36",x"2160",x"3bf6",x"3857",x"3903",x"2ec3",x"3e2f",x"3711",x"afec",x"2c2c",x"3beb",x"384f",x"3904"),
(x"2ea1",x"3e45",x"370f",x"9df0",x"2631",x"3bff",x"384b",x"391d",x"2eec",x"3e47",x"3713",x"ae9a",x"b366",x"3bbd",x"3850",x"391f",x"2f2d",x"3e3f",x"370e",x"26d5",x"a5c2",x"3bfe",x"3855",x"3917"),
(x"2f2d",x"3e3f",x"370e",x"26d5",x"a5c2",x"3bfe",x"3855",x"3917",x"2efb",x"3e3b",x"3713",x"a538",x"2c79",x"3bfa",x"3852",x"3912",x"2ea1",x"3e45",x"370f",x"9df0",x"2631",x"3bff",x"384b",x"391d"),
(x"2e69",x"3e40",x"370f",x"acd8",x"271d",x"3bf9",x"3848",x"3917",x"2efb",x"3e3b",x"3713",x"a538",x"2c79",x"3bfa",x"3852",x"3912",x"2e71",x"3e37",x"370f",x"aec5",x"9a24",x"3bf4",x"3849",x"390d"),
(x"2ec3",x"3e2f",x"3711",x"afec",x"2c2c",x"3beb",x"384f",x"3904",x"2efa",x"3e39",x"3713",x"a7e9",x"a849",x"3bfd",x"3852",x"390f",x"2f21",x"3e36",x"3710",x"ac5b",x"30a5",x"3be5",x"3855",x"390d"),
(x"2f4a",x"3e66",x"3712",x"af67",x"2981",x"3bf0",x"3858",x"3943",x"2fda",x"3e66",x"3715",x"a6c2",x"2c63",x"3bfa",x"3861",x"3943",x"2fa2",x"3e5e",x"3717",x"aff2",x"2a7d",x"3bed",x"385e",x"393b"),
(x"2e99",x"3e5f",x"3714",x"1553",x"2b62",x"3bfc",x"384d",x"393c",x"2ecb",x"3e55",x"3716",x"acd8",x"27e2",x"3bf9",x"3850",x"3930",x"2e81",x"3e5b",x"3712",x"b162",x"2345",x"3be2",x"384b",x"3937"),
(x"2ecb",x"3e55",x"3716",x"acd8",x"27e2",x"3bf9",x"3850",x"3930",x"2e99",x"3e5f",x"3714",x"1553",x"2b62",x"3bfc",x"384d",x"393c",x"2f0c",x"3e56",x"3716",x"2818",x"2d04",x"3bf8",x"3854",x"3931"),
(x"2f21",x"3e62",x"3711",x"240b",x"2d5c",x"3bf8",x"3855",x"393f",x"2f4f",x"3e59",x"3714",x"a4fd",x"2dab",x"3bf7",x"3858",x"3935",x"2f0c",x"3e56",x"3716",x"2818",x"2d04",x"3bf8",x"3854",x"3931"),
(x"2f79",x"3e5c",x"3714",x"b036",x"273e",x"3bed",x"385b",x"3939",x"2f21",x"3e62",x"3711",x"240b",x"2d5c",x"3bf8",x"3855",x"393f",x"2f3f",x"3e64",x"3711",x"b27d",x"975f",x"3bd5",x"3857",x"3941"),
(x"2ec5",x"3e7c",x"3711",x"b115",x"a7d5",x"3be4",x"384f",x"395c",x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2f3b",x"3e6b",x"3712",x"b146",x"ac91",x"3bde",x"3857",x"3949"),
(x"3017",x"3e77",x"3719",x"a3bb",x"a7ae",x"3bfe",x"3867",x"3957",x"2fe4",x"3e77",x"3718",x"2138",x"2e95",x"3bf4",x"3862",x"3957",x"3017",x"3e78",x"3719",x"a90e",x"2f00",x"3bf2",x"3867",x"3958"),
(x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2fd6",x"3e7d",x"3715",x"28bf",x"2fdb",x"3bef",x"3861",x"395d",x"2fe4",x"3e77",x"3718",x"2138",x"2e95",x"3bf4",x"3862",x"3957"),
(x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2fe4",x"3e77",x"3718",x"2138",x"2e95",x"3bf4",x"3862",x"3957",x"2fd8",x"3e76",x"3718",x"2b4f",x"a525",x"3bfc",x"3861",x"3956"),
(x"3002",x"3e68",x"3717",x"2d2d",x"aecd",x"3bed",x"3864",x"3946",x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"3022",x"3e6e",x"3718",x"2cf2",x"98ea",x"3bf9",x"3868",x"394c"),
(x"3022",x"3e6e",x"3718",x"2cf2",x"98ea",x"3bf9",x"3868",x"394c",x"3027",x"3e69",x"3712",x"359c",x"b36a",x"3b42",x"3869",x"3947",x"3002",x"3e68",x"3717",x"2d2d",x"aecd",x"3bed",x"3864",x"3946"),
(x"2f3b",x"3e6b",x"3712",x"b146",x"ac91",x"3bde",x"3857",x"3949",x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"2fe7",x"3e67",x"3716",x"b009",x"ada8",x"3be7",x"3862",x"3945"),
(x"2fda",x"3e66",x"3715",x"a6c2",x"2c63",x"3bfa",x"3861",x"3943",x"2f4a",x"3e66",x"3712",x"af67",x"2981",x"3bf0",x"3858",x"3943",x"2fe7",x"3e67",x"3716",x"b009",x"ada8",x"3be7",x"3862",x"3945"),
(x"2fc7",x"3e5d",x"3717",x"97c8",x"1f79",x"3c00",x"3860",x"3939",x"2fda",x"3e66",x"3715",x"a6c2",x"2c63",x"3bfa",x"3861",x"3943",x"2fe5",x"3e63",x"3714",x"a581",x"2e8a",x"3bf4",x"3862",x"3940"),
(x"302a",x"3e50",x"3714",x"2dba",x"a266",x"3bf7",x"386a",x"392b",x"3008",x"3e58",x"3715",x"a518",x"ad04",x"3bf9",x"3865",x"3934",x"3041",x"3e53",x"3714",x"175f",x"ac2c",x"3bfb",x"386d",x"392f"),
(x"302f",x"3e45",x"3715",x"3468",x"a47a",x"3bb0",x"386a",x"391f",x"302a",x"3e50",x"3714",x"2dba",x"a266",x"3bf7",x"386a",x"392b",x"3052",x"3e47",x"3712",x"3106",x"a73e",x"3be5",x"386f",x"3920"),
(x"3025",x"3e3d",x"3717",x"3273",x"af43",x"3bc8",x"3868",x"3915",x"302f",x"3e45",x"3715",x"3468",x"a47a",x"3bb0",x"386a",x"391f",x"3041",x"3e3b",x"3710",x"3550",x"ae33",x"3b81",x"386c",x"3913"),
(x"2fe6",x"3e36",x"3711",x"ae24",x"aa2b",x"3bf4",x"3862",x"390d",x"3025",x"3e3d",x"3717",x"3273",x"af43",x"3bc8",x"3868",x"3915",x"3015",x"3e33",x"3712",x"2b5f",x"a345",x"3bfc",x"3867",x"390a"),
(x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908",x"2f61",x"3e35",x"3713",x"25b5",x"37de",x"3af6",x"385a",x"390b",x"2fa3",x"3e35",x"3712",x"2dd2",x"304b",x"3be4",x"385e",x"390c"),
(x"2f5c",x"3e2c",x"3716",x"a553",x"b2c7",x"3bd1",x"385a",x"3901",x"2f2f",x"3e2e",x"3718",x"ae36",x"2160",x"3bf6",x"3857",x"3903",x"2f75",x"3e2e",x"3716",x"2f4d",x"2a5f",x"3bf0",x"385b",x"3903"),
(x"2f0a",x"3e2d",x"3716",x"af14",x"b29c",x"3bc6",x"3854",x"3902",x"2f2f",x"3e2e",x"3718",x"ae36",x"2160",x"3bf6",x"3857",x"3903",x"2f5c",x"3e2c",x"3716",x"a553",x"b2c7",x"3bd1",x"385a",x"3901"),
(x"2f93",x"3e1d",x"370f",x"aedc",x"acd0",x"3bee",x"385e",x"38f0",x"2f3e",x"3e22",x"3713",x"ada3",x"af14",x"3beb",x"3858",x"38f5",x"2fe6",x"3e22",x"3717",x"b0e7",x"b057",x"3bd4",x"3863",x"38f6"),
(x"2fc8",x"3e13",x"3716",x"aadf",x"26b5",x"3bfc",x"3862",x"38e4",x"2f93",x"3e1d",x"370f",x"aedc",x"acd0",x"3bee",x"385e",x"38f0",x"301b",x"3e14",x"3713",x"a9b8",x"26e9",x"3bfd",x"3869",x"38e7"),
(x"2fc8",x"3e13",x"3716",x"aadf",x"26b5",x"3bfc",x"3862",x"38e4",x"301b",x"3e14",x"3713",x"a9b8",x"26e9",x"3bfd",x"3869",x"38e7",x"3020",x"3e07",x"3717",x"abf6",x"a5ae",x"3bfb",x"386b",x"38d8"),
(x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4",x"3020",x"3e07",x"3717",x"abf6",x"a5ae",x"3bfb",x"386b",x"38d8",x"3031",x"3dfc",x"370f",x"36c9",x"afac",x"3b2e",x"386f",x"38cb"),
(x"3031",x"3dfc",x"370f",x"36c9",x"afac",x"3b2e",x"386f",x"38cb",x"302a",x"3df8",x"370d",x"3809",x"ae09",x"3add",x"386f",x"38c7",x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4"),
(x"3008",x"3de5",x"370e",x"2fd2",x"a717",x"3bef",x"386c",x"38b1",x"2f13",x"3dea",x"3715",x"2d56",x"a0d0",x"3bf8",x"385b",x"38b5",x"3013",x"3def",x"3712",x"29f0",x"ab1d",x"3bfa",x"386c",x"38bd"),
(x"2f27",x"3df7",x"3715",x"bb82",x"3440",x"330f",x"3b12",x"3a38",x"2f02",x"3df7",x"36eb",x"bb89",x"3473",x"31fc",x"3b17",x"3a37",x"2f97",x"3e08",x"370e",x"bb5f",x"35f1",x"2f4d",x"3b10",x"3a2e"),
(x"2ec4",x"3e97",x"3710",x"3bfd",x"2997",x"a09b",x"3a11",x"3a2e",x"2eca",x"3e9e",x"3714",x"3beb",x"b08b",x"98ea",x"3a11",x"3a32",x"2ec5",x"3e9c",x"36eb",x"3bf5",x"ae59",x"2467",x"3a16",x"3a31"),
(x"2f2f",x"3e80",x"3714",x"3b1c",x"3754",x"223f",x"3a10",x"3a22",x"2ed8",x"3e8e",x"3713",x"3ba5",x"3497",x"ac28",x"3a11",x"3a29",x"2ece",x"3e8d",x"36eb",x"3ba1",x"34cc",x"1f45",x"3a16",x"3a29"),
(x"2edf",x"3ea3",x"3712",x"3b76",x"b5c5",x"204d",x"3a11",x"3a34",x"2f06",x"3ea6",x"3714",x"395a",x"b9f1",x"2032",x"3a11",x"3a36",x"2ee8",x"3ea4",x"36eb",x"3ab1",x"b862",x"21f0",x"3a16",x"3a35"),
(x"2f3d",x"3ea8",x"3714",x"35bf",x"bb76",x"27db",x"3a11",x"3a39",x"2f38",x"3ea8",x"36eb",x"37e1",x"baf5",x"269a",x"3a16",x"3a38",x"2f06",x"3ea6",x"3714",x"395a",x"b9f1",x"2032",x"3a11",x"3a36"),
(x"2fa3",x"3eaa",x"3715",x"a836",x"bbfd",x"294c",x"3a11",x"3a3c",x"2f9e",x"3eaa",x"36eb",x"303c",x"bbeb",x"299b",x"3a16",x"3a3c",x"2f3d",x"3ea8",x"3714",x"35bf",x"bb76",x"27db",x"3a11",x"3a39"),
(x"3004",x"3ea9",x"3716",x"b86f",x"baa7",x"2604",x"3a11",x"3a40",x"3003",x"3ea9",x"36eb",x"b868",x"baab",x"296a",x"3a16",x"3a3f",x"2fa3",x"3eaa",x"3715",x"a836",x"bbfd",x"294c",x"3a11",x"3a3c"),
(x"3004",x"3ea9",x"3716",x"b86f",x"baa7",x"2604",x"3a11",x"3a40",x"302c",x"3ea3",x"3714",x"bb01",x"b7b5",x"2839",x"3a12",x"3a44",x"3003",x"3ea9",x"36eb",x"b868",x"baab",x"296a",x"3a16",x"3a3f"),
(x"3036",x"3e9d",x"3714",x"bbe6",x"310f",x"9bfc",x"3a12",x"3a47",x"3036",x"3e9d",x"36eb",x"bbf9",x"ad11",x"2511",x"3a17",x"3a46",x"302c",x"3ea3",x"3714",x"bb01",x"b7b5",x"2839",x"3a12",x"3a44"),
(x"3026",x"3e98",x"3715",x"b928",x"3a1d",x"1553",x"3a12",x"3a49",x"3029",x"3e99",x"36eb",x"b90c",x"3a34",x"2532",x"3a17",x"3a49",x"3036",x"3e9d",x"3714",x"bbe6",x"310f",x"9bfc",x"3a12",x"3a47"),
(x"3026",x"3e98",x"3715",x"b928",x"3a1d",x"1553",x"3a12",x"3a49",x"3006",x"3e98",x"3714",x"2fe2",x"3bee",x"28fd",x"3a12",x"3a4b",x"3029",x"3e99",x"36eb",x"b90c",x"3a34",x"2532",x"3a17",x"3a49"),
(x"3006",x"3e98",x"3714",x"2fe2",x"3bee",x"28fd",x"3a12",x"3a4b",x"2fd7",x"3e9a",x"3711",x"364f",x"3b52",x"2d1b",x"3a13",x"3a4d",x"3004",x"3e98",x"36eb",x"35dd",x"3b6d",x"2be9",x"3a17",x"3a4b"),
(x"2f89",x"3e8c",x"3713",x"bbc2",x"b3a4",x"298a",x"3a12",x"3a59",x"2f82",x"3e8c",x"36eb",x"bbf6",x"aa70",x"2d60",x"3a17",x"3a5a",x"2f73",x"3e8e",x"3711",x"ba7a",x"b8af",x"2839",x"3a12",x"3a58"),
(x"2fd7",x"3e9a",x"3711",x"364f",x"3b52",x"2d1b",x"3a13",x"3a4d",x"2f85",x"3e9a",x"3710",x"b416",x"3bad",x"2f8d",x"3a13",x"3a50",x"2fdd",x"3e9b",x"36eb",x"32b1",x"3bc8",x"2e54",x"3a18",x"3a4d"),
(x"2eec",x"3e47",x"3713",x"3583",x"3b63",x"3153",x"3b1c",x"3b74",x"2efa",x"3e48",x"36eb",x"35e4",x"3b4d",x"31a2",x"3b21",x"3b72",x"2f31",x"3e42",x"370f",x"3a9c",x"3854",x"30fa",x"3b1b",x"3b71"),
(x"2f27",x"3df7",x"3715",x"bb82",x"3440",x"330f",x"3b12",x"3a38",x"2f13",x"3dea",x"3715",x"bbc5",x"ab9a",x"3358",x"3b13",x"3a3f",x"2f02",x"3df7",x"36eb",x"bb89",x"3473",x"31fc",x"3b17",x"3a37"),
(x"2f73",x"3e8e",x"3711",x"b40c",x"a6c2",x"3bbc",x"385a",x"3970",x"2f51",x"3e90",x"3710",x"a856",x"29ab",x"3bfc",x"3858",x"3973",x"2fe3",x"3e8b",x"3718",x"ab65",x"3528",x"3b8f",x"3862",x"396d"),
(x"3006",x"3df4",x"3715",x"3bd7",x"31f9",x"2c2a",x"3b0d",x"3a55",x"3008",x"3df6",x"3716",x"38de",x"ba57",x"297d",x"3b0c",x"3a55",x"300a",x"3df5",x"36eb",x"3be3",x"ace8",x"30c3",x"3b11",x"3a58"),
(x"3015",x"3e33",x"3712",x"384e",x"bab0",x"2ec8",x"3a23",x"3a4d",x"3041",x"3e3b",x"3710",x"3b6a",x"b5bb",x"2efe",x"3a23",x"3a52",x"301f",x"3e33",x"36eb",x"3958",x"b9de",x"2fe4",x"3a27",x"3a4d"),
(x"2f5e",x"3e98",x"3711",x"ba7f",x"3887",x"3089",x"3a13",x"3a52",x"2f4e",x"3e99",x"36eb",x"baa4",x"3859",x"2fe4",x"3a18",x"3a52",x"2f85",x"3e9a",x"3710",x"b416",x"3bad",x"2f8d",x"3a13",x"3a50"),
(x"2fcc",x"3e88",x"3718",x"3be6",x"b09f",x"2baa",x"3b45",x"38d6",x"2fd8",x"3e89",x"36eb",x"3be6",x"b08e",x"2c41",x"3b49",x"38d4",x"2fc7",x"3e7f",x"3715",x"3bfa",x"2710",x"2c48",x"3b44",x"38d3"),
(x"2f5e",x"3e98",x"3711",x"ba7f",x"3887",x"3089",x"3a13",x"3a52",x"2f45",x"3e94",x"3710",x"bbcc",x"3227",x"2f2e",x"3a13",x"3a54",x"2f4e",x"3e99",x"36eb",x"baa4",x"3859",x"2fe4",x"3a18",x"3a52"),
(x"2f31",x"3e42",x"370f",x"3a9c",x"3854",x"30fa",x"3b1b",x"3b71",x"2f46",x"3e42",x"36eb",x"3b7d",x"3521",x"3096",x"3b1f",x"3b6f",x"2f2d",x"3e3f",x"370e",x"3b25",x"b70d",x"2d6a",x"3b1a",x"3b70"),
(x"2e99",x"3e5f",x"3714",x"b972",x"39bb",x"30de",x"3b4b",x"38fe",x"2e90",x"3e61",x"36eb",x"b6fe",x"3b25",x"2ea4",x"3b4e",x"38fe",x"2f21",x"3e62",x"3711",x"b4dc",x"3b97",x"2d61",x"3b4b",x"38fc"),
(x"2f73",x"3e8e",x"3711",x"ba7a",x"b8af",x"2839",x"3a12",x"3a58",x"2f71",x"3e8d",x"36eb",x"b9db",x"b96c",x"2c1a",x"3a17",x"3a59",x"2f51",x"3e90",x"3710",x"bb2f",x"b6d9",x"2e52",x"3a13",x"3a56"),
(x"2f75",x"3e2e",x"3716",x"37e9",x"baf1",x"2aa7",x"3a22",x"3a46",x"3015",x"3e33",x"3712",x"384e",x"bab0",x"2ec8",x"3a23",x"3a4d",x"2f6d",x"3e2d",x"36eb",x"3776",x"bb0b",x"2d41",x"3a27",x"3a45"),
(x"2fd6",x"3e7d",x"3715",x"395d",x"39e3",x"2de3",x"3b44",x"38d3",x"2fc7",x"3e7f",x"3715",x"3bfa",x"2710",x"2c48",x"3b44",x"38d3",x"2fd9",x"3e7e",x"36eb",x"39df",x"3964",x"2d28",x"3b47",x"38d2"),
(x"2efb",x"3e3b",x"3713",x"3b5b",x"b634",x"2c08",x"3b18",x"3b6e",x"2f2d",x"3e3f",x"370e",x"3b25",x"b70d",x"2d6a",x"3b1a",x"3b70",x"2f02",x"3e3a",x"36eb",x"3ad3",x"b822",x"2c4d",x"3b1c",x"3b6b"),
(x"2fc8",x"3e13",x"3716",x"bbff",x"a0c2",x"2138",x"3b0e",x"3a29",x"2f97",x"3e08",x"370e",x"bb5f",x"35f1",x"2f4d",x"3b10",x"3a2e",x"2fc6",x"3e13",x"36eb",x"bbfe",x"9ea7",x"2828",x"3b13",x"3a27"),
(x"2f75",x"3e2e",x"3716",x"37e9",x"baf1",x"2aa7",x"3a22",x"3a46",x"2f6d",x"3e2d",x"36eb",x"3776",x"bb0b",x"2d41",x"3a27",x"3a45",x"2f5c",x"3e2c",x"3716",x"3bde",x"b1b5",x"2825",x"3a22",x"3a45"),
(x"3017",x"3e78",x"3719",x"39a6",x"3994",x"2fb1",x"3b43",x"38d1",x"2fd6",x"3e7d",x"3715",x"395d",x"39e3",x"2de3",x"3b44",x"38d3",x"3026",x"3e78",x"36eb",x"39ed",x"394b",x"2f45",x"3b46",x"38cf"),
(x"2f3f",x"3e64",x"3711",x"bb12",x"3763",x"2ca3",x"3b4b",x"38fb",x"2f21",x"3e62",x"3711",x"b4dc",x"3b97",x"2d61",x"3b4b",x"38fc",x"2f2b",x"3e63",x"36eb",x"b7d8",x"3af6",x"2a35",x"3b4f",x"38fc"),
(x"2efa",x"3e39",x"3713",x"3b09",x"3791",x"2ab8",x"3b41",x"3916",x"2efb",x"3e3b",x"3713",x"3b5b",x"b634",x"2c08",x"3b41",x"3917",x"2f01",x"3e39",x"36eb",x"39e9",x"3955",x"2e31",x"3b45",x"3917"),
(x"2fc8",x"3e13",x"3716",x"bbff",x"a0c2",x"2138",x"3b0e",x"3a29",x"2fc6",x"3e13",x"36eb",x"bbfe",x"9ea7",x"2828",x"3b13",x"3a27",x"2f93",x"3e1d",x"370f",x"bad7",x"b821",x"29e6",x"3b0e",x"3a23"),
(x"2f5c",x"3e2c",x"3716",x"3bde",x"b1b5",x"2825",x"3a22",x"3a45",x"2f62",x"3e2c",x"36eb",x"3b24",x"371c",x"2cde",x"3a27",x"3a45",x"2f72",x"3e29",x"3714",x"39e8",x"3951",x"2f27",x"3a22",x"3a44"),
(x"3017",x"3e78",x"3719",x"39a6",x"3994",x"2fb1",x"3b43",x"38d1",x"3026",x"3e78",x"36eb",x"39ed",x"394b",x"2f45",x"3b46",x"38cf",x"3017",x"3e77",x"3719",x"3250",x"bbca",x"2f22",x"3b42",x"38d1"),
(x"2f4a",x"3e66",x"3712",x"bbf7",x"a83f",x"2d8f",x"3b4b",x"38fb",x"2f3c",x"3e66",x"36eb",x"bbf8",x"2379",x"2d44",x"3b4f",x"38fb",x"2f3b",x"3e6b",x"3712",x"bb92",x"b509",x"2cb4",x"3b4c",x"38f9"),
(x"2f21",x"3e36",x"3710",x"3833",x"3ac7",x"2d1d",x"3b42",x"3915",x"2efa",x"3e39",x"3713",x"3b09",x"3791",x"2ab8",x"3b41",x"3916",x"2f01",x"3e39",x"36eb",x"39e9",x"3955",x"2e31",x"3b45",x"3917"),
(x"2f3e",x"3e22",x"3713",x"b7c3",x"baf3",x"2e28",x"3b0c",x"3a20",x"2f93",x"3e1d",x"370f",x"bad7",x"b821",x"29e6",x"3b0e",x"3a23",x"2f33",x"3e21",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3b11",x"3a1e"),
(x"2f72",x"3e29",x"3714",x"39e8",x"3951",x"2f27",x"3a22",x"3a44",x"2f83",x"3e2a",x"36eb",x"397a",x"39b6",x"3099",x"3a27",x"3a44",x"2fe6",x"3e22",x"3717",x"3a77",x"3889",x"310c",x"3a22",x"3a3e"),
(x"2fe4",x"3e77",x"3718",x"30c5",x"bbe6",x"2ad9",x"3b41",x"38d0",x"3017",x"3e77",x"3719",x"3250",x"bbca",x"2f22",x"3b42",x"38d1",x"2fda",x"3e76",x"36eb",x"3b01",x"b745",x"3141",x"3b44",x"38ce"),
(x"2f3b",x"3e6b",x"3712",x"bb92",x"b509",x"2cb4",x"3b4c",x"38f9",x"2f33",x"3e6a",x"36eb",x"bb57",x"b625",x"2e99",x"3b4f",x"38f9",x"2ec5",x"3e7c",x"3711",x"bb70",x"b585",x"3014",x"3b4c",x"38f4"),
(x"2fa3",x"3e35",x"3712",x"b2e8",x"3bcb",x"2c10",x"3b42",x"3913",x"2f61",x"3e35",x"3713",x"30a8",x"3be9",x"22dc",x"3b42",x"3914",x"2f69",x"3e35",x"36eb",x"3046",x"3be8",x"2cb7",x"3b45",x"3914"),
(x"2f3e",x"3e22",x"3713",x"b7c3",x"baf3",x"2e28",x"3b18",x"3b93",x"2f33",x"3e21",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3b1d",x"3b96",x"2f20",x"3e21",x"3712",x"3721",x"bb24",x"2bf2",x"3b19",x"3b92"),
(x"2fe6",x"3e22",x"3717",x"3a77",x"3889",x"310c",x"3a22",x"3a3e",x"3000",x"3e23",x"36eb",x"3aff",x"373c",x"3197",x"3a27",x"3a3e",x"301b",x"3e14",x"3713",x"3bc6",x"31be",x"30de",x"3a22",x"3a37"),
(x"2ec5",x"3e7c",x"3711",x"bb70",x"b585",x"3014",x"3b4c",x"38f4",x"2ea7",x"3e7d",x"36eb",x"bb99",x"b45f",x"30d6",x"3b50",x"38f4",x"2e95",x"3e8c",x"3711",x"bbe4",x"ad1e",x"308c",x"3b4d",x"38f0"),
(x"3025",x"3e3d",x"3717",x"bb6f",x"35e5",x"261e",x"3b43",x"390f",x"2fe6",x"3e36",x"3711",x"b934",x"3a0e",x"2c16",x"3b43",x"3912",x"3021",x"3e3d",x"36eb",x"baaf",x"3860",x"2a70",x"3b47",x"3910"),
(x"2f20",x"3e21",x"3712",x"3721",x"bb24",x"2bf2",x"3b19",x"3b92",x"2f19",x"3e20",x"36eb",x"38ae",x"ba73",x"2d49",x"3b1d",x"3b95",x"2ef3",x"3e1f",x"3711",x"35dd",x"bb65",x"2eae",x"3b1a",x"3b91"),
(x"3020",x"3e07",x"3717",x"3bf0",x"2f10",x"2aec",x"3a21",x"3a30",x"301b",x"3e14",x"3713",x"3bc6",x"31be",x"30de",x"3a22",x"3a37",x"3025",x"3e07",x"36eb",x"3bea",x"2e09",x"2f12",x"3a26",x"3a2f"),
(x"2fd8",x"3e76",x"3718",x"3af6",x"37e0",x"2460",x"3b7d",x"366f",x"2fe4",x"3e77",x"3718",x"30c5",x"bbe6",x"2ad9",x"3b7d",x"3670",x"2fda",x"3e76",x"36eb",x"3b01",x"b745",x"3141",x"3b83",x"3670"),
(x"2e95",x"3e9d",x"3714",x"bbec",x"2d02",x"2f52",x"3b4d",x"38eb",x"2e95",x"3e8c",x"3711",x"bbe4",x"ad1e",x"308c",x"3b4d",x"38f0",x"2e82",x"3e9d",x"36eb",x"bbe8",x"2d66",x"3010",x"3b50",x"38eb"),
(x"302f",x"3e45",x"3715",x"bbfe",x"a412",x"2867",x"3b44",x"390d",x"3025",x"3e3d",x"3717",x"bb6f",x"35e5",x"261e",x"3b43",x"390f",x"302e",x"3e45",x"36eb",x"bbfa",x"2c62",x"2617",x"3b48",x"390e"),
(x"2ef3",x"3e1f",x"3711",x"35dd",x"bb65",x"2eae",x"3b1a",x"3b91",x"2efa",x"3e1e",x"36eb",x"2e29",x"bbe6",x"3005",x"3b1e",x"3b94",x"2eb1",x"3e20",x"3712",x"b5a6",x"bb63",x"30cc",x"3b1b",x"3b8f"),
(x"3020",x"3e07",x"3717",x"3bf0",x"2f10",x"2aec",x"3a21",x"3a30",x"3025",x"3e07",x"36eb",x"3bea",x"2e09",x"2f12",x"3a26",x"3a2f",x"3031",x"3dfc",x"370f",x"3bdd",x"30de",x"2e6c",x"3a21",x"3a2a"),
(x"3006",x"3e73",x"3715",x"39d1",x"3974",x"2cc6",x"3b7e",x"366a",x"3016",x"3e72",x"36eb",x"3a0e",x"3929",x"2e76",x"3b83",x"3669",x"3022",x"3e6e",x"3718",x"3b13",x"3732",x"2fec",x"3b7d",x"3663"),
(x"2e95",x"3e9d",x"3714",x"bbec",x"2d02",x"2f52",x"3b4d",x"38eb",x"2e82",x"3e9d",x"36eb",x"bbe8",x"2d66",x"3010",x"3b50",x"38eb",x"2eb5",x"3ea5",x"3712",x"bb45",x"3640",x"30a6",x"3b4d",x"38e9"),
(x"2f45",x"3e94",x"3710",x"bbcc",x"3227",x"2f2e",x"3a13",x"3a54",x"2f51",x"3e90",x"3710",x"bb2f",x"b6d9",x"2e52",x"3a13",x"3a56",x"2f36",x"3e94",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3a18",x"3a55"),
(x"302a",x"3e50",x"3714",x"bb81",x"b558",x"2da6",x"3b46",x"390a",x"302f",x"3e45",x"3715",x"bbfe",x"a412",x"2867",x"3b44",x"390d",x"3025",x"3e4f",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"3b49",x"390b"),
(x"2eb1",x"3e20",x"3712",x"b5a6",x"bb63",x"30cc",x"3b1b",x"3b8f",x"2e9b",x"3e1f",x"36eb",x"b913",x"ba0d",x"310f",x"3b20",x"3b91",x"2e89",x"3e24",x"3711",x"bbb2",x"b32f",x"30f4",x"3b1c",x"3b8d"),
(x"3031",x"3dfc",x"370f",x"3bdd",x"30de",x"2e6c",x"3a21",x"3a2a",x"303b",x"3dfc",x"36eb",x"3be4",x"2adf",x"30ee",x"3a26",x"3a29",x"302a",x"3df8",x"370d",x"3b0d",x"b70c",x"3169",x"3a21",x"3a28"),
(x"3022",x"3e6e",x"3718",x"3b13",x"3732",x"2fec",x"3b7d",x"3663",x"302e",x"3e6e",x"36eb",x"3bbf",x"3333",x"2ed0",x"3b83",x"3663",x"3027",x"3e69",x"3712",x"3bf0",x"ac20",x"2e95",x"3b7e",x"365f"),
(x"2eb5",x"3ea5",x"3712",x"bb45",x"3640",x"30a6",x"3b4d",x"38e9",x"2ea5",x"3ea6",x"36eb",x"bab2",x"3834",x"30cf",x"3b50",x"38e8",x"2f1a",x"3eac",x"3715",x"b93c",x"39e9",x"311d",x"3b4d",x"38e6"),
(x"3008",x"3e58",x"3715",x"ba65",x"b8c1",x"2d9e",x"3b47",x"3908",x"302a",x"3e50",x"3714",x"bb81",x"b558",x"2da6",x"3b46",x"390a",x"3001",x"3e57",x"36eb",x"bac2",x"b833",x"2e85",x"3b4a",x"3909"),
(x"2e89",x"3e24",x"3711",x"bbb2",x"b32f",x"30f4",x"3b1c",x"3b8d",x"2e73",x"3e23",x"36eb",x"bbe5",x"2dbc",x"3036",x"3b20",x"3b8e",x"2ea4",x"3e29",x"3712",x"bae4",x"37c3",x"30c9",x"3b1c",x"3b8a"),
(x"301d",x"3df6",x"3713",x"3451",x"bbac",x"2d81",x"3a20",x"3a27",x"302a",x"3df8",x"370d",x"3b0d",x"b70c",x"3169",x"3a21",x"3a28",x"3020",x"3df5",x"36eb",x"3571",x"bb6d",x"30cc",x"3a25",x"3a25"),
(x"3027",x"3e69",x"3712",x"3bf0",x"ac20",x"2e95",x"3b7e",x"365f",x"302b",x"3e68",x"36eb",x"3bbf",x"b371",x"2dad",x"3b83",x"365d",x"301e",x"3e68",x"3712",x"3297",x"bbcc",x"2d84",x"3b7e",x"365d"),
(x"2f1a",x"3eac",x"3715",x"b93c",x"39e9",x"311d",x"3b4d",x"38e6",x"2f13",x"3eae",x"36eb",x"b7cb",x"3ae6",x"3068",x"3b50",x"38e6",x"2f91",x"3eaf",x"3715",x"9ef6",x"3bee",x"302a",x"3b4c",x"38e4"),
(x"2fc7",x"3e5d",x"3717",x"b939",x"ba0b",x"29e0",x"3b47",x"3906",x"3008",x"3e58",x"3715",x"ba65",x"b8c1",x"2d9e",x"3b47",x"3908",x"2fc1",x"3e5c",x"36eb",x"b9cd",x"b979",x"2caa",x"3b4b",x"3907"),
(x"2ea4",x"3e29",x"3712",x"bae4",x"37c3",x"30c9",x"3b1c",x"3b8a",x"2e9a",x"3e2b",x"36eb",x"b902",x"3a23",x"306a",x"3b21",x"3b8a",x"2eea",x"3e2b",x"3713",x"b607",x"3b5e",x"2e4f",x"3b1d",x"3b87"),
(x"3008",x"3df6",x"3716",x"38de",x"ba57",x"297d",x"3a1f",x"3a26",x"301d",x"3df6",x"3713",x"3451",x"bbac",x"2d81",x"3a20",x"3a27",x"300a",x"3df5",x"36eb",x"3be3",x"ace8",x"30c3",x"3a24",x"3a23"),
(x"3002",x"3e68",x"3717",x"2a07",x"bbfc",x"284d",x"3b7d",x"3659",x"301e",x"3e68",x"3712",x"3297",x"bbcc",x"2d84",x"3b7e",x"365d",x"2ffe",x"3e67",x"36eb",x"2c58",x"bbf7",x"2bc5",x"3b82",x"3657"),
(x"300a",x"3ead",x"3713",x"382e",x"3aba",x"306c",x"3b4c",x"38e2",x"2f91",x"3eaf",x"3715",x"9ef6",x"3bee",x"302a",x"3b4c",x"38e4",x"3007",x"3eae",x"36eb",x"366a",x"3b44",x"2f81",x"3b4f",x"38e1"),
(x"2fa2",x"3e5e",x"3717",x"2c95",x"bbf9",x"2914",x"3b48",x"3906",x"2fc7",x"3e5d",x"3717",x"b939",x"ba0b",x"29e0",x"3b47",x"3906",x"2fa3",x"3e5e",x"36eb",x"35a5",x"bb74",x"2d53",x"3b4b",x"3907"),
(x"2f0a",x"3e2d",x"3716",x"bac7",x"b83c",x"283f",x"3b1c",x"3b86",x"2eea",x"3e2b",x"3713",x"b607",x"3b5e",x"2e4f",x"3b1d",x"3b87",x"2f03",x"3e2d",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3b22",x"3b87"),
(x"2f97",x"3e08",x"370e",x"b004",x"271d",x"3bef",x"3860",x"38d8",x"2fc8",x"3e13",x"3716",x"aadf",x"26b5",x"3bfc",x"3862",x"38e4",x"3020",x"3e07",x"3717",x"abf6",x"a5ae",x"3bfb",x"386b",x"38d8"),
(x"3002",x"3e68",x"3717",x"2a07",x"bbfc",x"284d",x"3b7d",x"3659",x"2ffe",x"3e67",x"36eb",x"2c58",x"bbf7",x"2bc5",x"3b82",x"3657",x"2fe7",x"3e67",x"3716",x"38f4",x"ba42",x"2c09",x"3b7d",x"3657"),
(x"3046",x"3ea6",x"3715",x"3ae0",x"37cf",x"30d4",x"3b4b",x"38df",x"300a",x"3ead",x"3713",x"382e",x"3aba",x"306c",x"3b4c",x"38e2",x"3051",x"3ea8",x"36eb",x"39f2",x"3938",x"30b5",x"3b4e",x"38de"),
(x"2f79",x"3e5c",x"3714",x"39a7",x"b99f",x"2d1e",x"3b48",x"3905",x"2fa2",x"3e5e",x"3717",x"2c95",x"bbf9",x"2914",x"3b48",x"3906",x"2fa3",x"3e5e",x"36eb",x"35a5",x"bb74",x"2d53",x"3b4b",x"3907"),
(x"2f0a",x"3e2d",x"3716",x"bac7",x"b83c",x"283f",x"3b1c",x"3b86",x"2f03",x"3e2d",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3b22",x"3b87",x"2ec3",x"3e2f",x"3711",x"b8c8",x"ba4e",x"30a8",x"3b1d",x"3b84"),
(x"2fe7",x"3e67",x"3716",x"38f4",x"ba42",x"2c09",x"3b7d",x"3657",x"2fea",x"3e66",x"36eb",x"3a75",x"b8ad",x"2ccc",x"3b82",x"3655",x"2fda",x"3e66",x"3715",x"3b3f",x"b6b6",x"2b9d",x"3b7d",x"3655"),
(x"3061",x"3e9d",x"3715",x"3bec",x"2be2",x"2fce",x"3b4a",x"38dc",x"3046",x"3ea6",x"3715",x"3ae0",x"37cf",x"30d4",x"3b4b",x"38df",x"306a",x"3e9e",x"36eb",x"3bc4",x"327a",x"3012",x"3b4d",x"38dc"),
(x"2f4f",x"3e59",x"3714",x"397e",x"b9c5",x"2dbf",x"3b49",x"3904",x"2f4c",x"3e58",x"36eb",x"3976",x"b9cc",x"2dcc",x"3b4c",x"3905",x"2f0c",x"3e56",x"3716",x"37d5",x"baf0",x"2d8e",x"3b4a",x"3903"),
(x"2ec3",x"3e2f",x"3711",x"b8c8",x"ba4e",x"30a8",x"3b1d",x"3b84",x"2ea2",x"3e2e",x"36eb",x"b9ec",x"b92b",x"31e4",x"3b22",x"3b83",x"2e71",x"3e37",x"370f",x"bb4b",x"b5cc",x"3223",x"3b1e",x"3b7f"),
(x"3013",x"3def",x"3712",x"3bcf",x"3082",x"3141",x"3b0f",x"3a53",x"3023",x"3def",x"36eb",x"3bdb",x"9c67",x"320a",x"3b13",x"3a55",x"3008",x"3de5",x"370e",x"3b7b",x"b4a9",x"3270",x"3b12",x"3a4e"),
(x"2fe5",x"3e63",x"3714",x"b879",x"b47b",x"3a3d",x"3a1f",x"3a69",x"2fda",x"3e66",x"3715",x"3a5f",x"3873",x"3389",x"3a20",x"3a6a",x"300d",x"3e5f",x"3718",x"3ac6",x"37dc",x"3285",x"3a20",x"3a66"),
(x"3058",x"3e95",x"3717",x"3b55",x"b5fd",x"307e",x"3b49",x"38da",x"3061",x"3e9d",x"3715",x"3bec",x"2be2",x"2fce",x"3b4a",x"38dc",x"3065",x"3e94",x"36eb",x"3b6e",x"b575",x"309e",x"3b4c",x"38d9"),
(x"2f2f",x"3e80",x"3714",x"b05e",x"a194",x"3bec",x"3856",x"3961",x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2ec5",x"3e7c",x"3711",x"b115",x"a7d5",x"3be4",x"384f",x"395c"),
(x"2f0c",x"3e56",x"3716",x"37d5",x"baf0",x"2d8e",x"3b4a",x"3903",x"2f11",x"3e55",x"36eb",x"353f",x"bb87",x"2d28",x"3b4d",x"3904",x"2ecb",x"3e55",x"3716",x"a345",x"bbf7",x"2dcc",x"3b4a",x"3901"),
(x"2e71",x"3e37",x"370f",x"bb4b",x"b5cc",x"3223",x"3b1e",x"3b7f",x"2e56",x"3e37",x"36eb",x"bbbc",x"b212",x"3175",x"3b22",x"3b7e",x"2e69",x"3e40",x"370f",x"bbd3",x"2f46",x"3182",x"3b1d",x"3b7a"),
(x"300d",x"3e5f",x"3718",x"3ac6",x"37dc",x"3286",x"3a20",x"3a66",x"3025",x"3e5f",x"36eb",x"3afe",x"375c",x"30f4",x"3a26",x"3a65",x"3041",x"3e53",x"3714",x"3b6b",x"3587",x"3096",x"3a21",x"3a5f"),
(x"3058",x"3e95",x"3717",x"3b55",x"b5fd",x"307e",x"3b49",x"38da",x"3065",x"3e94",x"36eb",x"3b6e",x"b575",x"309e",x"3b4c",x"38d9",x"3030",x"3e8e",x"3711",x"38a4",x"ba69",x"309a",x"3b48",x"38d8"),
(x"2ecb",x"3e55",x"3716",x"a345",x"bbf7",x"2dcc",x"3b4a",x"3901",x"2ec4",x"3e54",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"3b4d",x"3902",x"2e97",x"3e57",x"3714",x"b976",x"b9c0",x"3023",x"3b4b",x"3901"),
(x"2e69",x"3e40",x"370f",x"bbd3",x"2f46",x"3182",x"3b1d",x"3b7a",x"2e52",x"3e41",x"36eb",x"bb61",x"35a0",x"3119",x"3b22",x"3b79",x"2ea1",x"3e45",x"370f",x"b891",x"3a72",x"30f5",x"3b1d",x"3b77"),
(x"3008",x"3de5",x"370e",x"3b7b",x"b4a9",x"3270",x"3b12",x"3a4e",x"3014",x"3de3",x"36eb",x"3ade",x"b7ab",x"31d3",x"3b16",x"3a50",x"2fa8",x"3ddc",x"3712",x"38b5",x"ba3e",x"32bd",x"3b13",x"3a49"),
(x"3041",x"3e53",x"3714",x"3b6b",x"3587",x"3096",x"3a21",x"3a5f",x"304c",x"3e53",x"36eb",x"3bba",x"3376",x"2f14",x"3a26",x"3a5f",x"3052",x"3e47",x"3712",x"3bf0",x"2a00",x"2f46",x"3a22",x"3a58"),
(x"2fe3",x"3e8b",x"3718",x"38ae",x"ba78",x"2b79",x"3b46",x"38d6",x"3030",x"3e8e",x"3711",x"38a4",x"ba69",x"309a",x"3b48",x"38d8",x"2fed",x"3e8b",x"36eb",x"360d",x"bb5a",x"2ef3",x"3b49",x"38d5"),
(x"2e97",x"3e57",x"3714",x"b976",x"b9c0",x"3023",x"3b4b",x"3901",x"2e81",x"3e56",x"36eb",x"bacb",x"b812",x"3065",x"3b4e",x"3901",x"2e81",x"3e5b",x"3712",x"bbe0",x"ae5e",x"30a3",x"3b4b",x"38ff"),
(x"2eec",x"3e47",x"3713",x"3583",x"3b63",x"3153",x"3b1c",x"3b74",x"2ea1",x"3e45",x"370f",x"b891",x"3a72",x"30f5",x"3b1d",x"3b77",x"2efa",x"3e48",x"36eb",x"35e4",x"3b4d",x"31a2",x"3b21",x"3b72"),
(x"2f67",x"3ddc",x"3716",x"badd",x"b75a",x"334d",x"3b13",x"3a46",x"2fa8",x"3ddc",x"3712",x"38b5",x"ba3e",x"32bd",x"3b13",x"3a49",x"2f52",x"3dd9",x"36eb",x"b996",x"b95e",x"33ec",x"3b19",x"3a47"),
(x"3052",x"3e47",x"3712",x"3bf0",x"2a00",x"2f46",x"3a22",x"3a58",x"305b",x"3e46",x"36eb",x"3bef",x"ad09",x"2e69",x"3a27",x"3a58",x"3041",x"3e3b",x"3710",x"3b6a",x"b5bb",x"2efe",x"3a23",x"3a52"),
(x"2fcc",x"3e88",x"3718",x"3be6",x"b09f",x"2baa",x"3b45",x"38d6",x"2fe3",x"3e8b",x"3718",x"38ae",x"ba78",x"2b79",x"3b46",x"38d6",x"2fd8",x"3e89",x"36eb",x"3be6",x"b08e",x"2c41",x"3b49",x"38d4"),
(x"2e81",x"3e5b",x"3712",x"bbe0",x"ae5e",x"30a3",x"3b4b",x"38ff",x"2e6a",x"3e5c",x"36eb",x"bbcf",x"3174",x"3043",x"3b4e",x"3900",x"2e99",x"3e5f",x"3714",x"b972",x"39bb",x"30de",x"3b4b",x"38fe"),
(x"2e95",x"3e8c",x"3711",x"acd1",x"a504",x"3bf9",x"384b",x"396e",x"2e95",x"3e9d",x"3714",x"2eb0",x"a8fa",x"3bf3",x"384b",x"3981",x"2ec4",x"3e97",x"3710",x"2828",x"a60a",x"3bfe",x"384e",x"397a"),
(x"2eb5",x"3ea5",x"3712",x"a587",x"a08e",x"3bff",x"384c",x"398a",x"2f06",x"3ea6",x"3714",x"a8bf",x"ac22",x"3bfa",x"3852",x"398b",x"2edf",x"3ea3",x"3712",x"2953",x"a7ae",x"3bfd",x"384f",x"3987"),
(x"2eb5",x"3ea5",x"3712",x"a587",x"a08e",x"3bff",x"384c",x"398a",x"2f1a",x"3eac",x"3715",x"a0ea",x"aafd",x"3bfc",x"3853",x"3993",x"2f06",x"3ea6",x"3714",x"a8bf",x"ac22",x"3bfa",x"3852",x"398b"),
(x"2f1a",x"3eac",x"3715",x"a0ea",x"aafd",x"3bfc",x"3853",x"3993",x"2f91",x"3eaf",x"3715",x"27db",x"a9b2",x"3bfc",x"385a",x"3996",x"2f3d",x"3ea8",x"3714",x"231d",x"ab5f",x"3bfc",x"3855",x"398e"),
(x"2f91",x"3eaf",x"3715",x"27db",x"a9b2",x"3bfc",x"385a",x"3996",x"300a",x"3ead",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3863",x"3994",x"2fa3",x"3eaa",x"3715",x"270a",x"2779",x"3bfe",x"385c",x"3991"),
(x"300a",x"3ead",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3863",x"3994",x"3046",x"3ea6",x"3715",x"a266",x"1d87",x"3bff",x"386b",x"398d",x"3004",x"3ea9",x"3716",x"24bc",x"2ceb",x"3bf9",x"3862",x"3990"),
(x"3046",x"3ea6",x"3715",x"a266",x"1d87",x"3bff",x"386b",x"398d",x"3061",x"3e9d",x"3715",x"a891",x"27ce",x"3bfd",x"386f",x"3983",x"302c",x"3ea3",x"3714",x"a8e0",x"a99e",x"3bfc",x"3868",x"3989"),
(x"3036",x"3e9d",x"3714",x"a538",x"29ab",x"3bfd",x"386a",x"3983",x"3061",x"3e9d",x"3715",x"a891",x"27ce",x"3bfd",x"386f",x"3983",x"3026",x"3e98",x"3715",x"ac67",x"a8a5",x"3bf9",x"3868",x"397d"),
(x"3058",x"3e95",x"3717",x"ad06",x"a793",x"3bf8",x"386f",x"397a",x"3030",x"3e8e",x"3711",x"a8d9",x"252b",x"3bfe",x"386a",x"3972",x"3026",x"3e98",x"3715",x"ac67",x"a8a5",x"3bf9",x"3868",x"397d"),
(x"3006",x"3e98",x"3714",x"aa45",x"ab10",x"3bfa",x"3864",x"397c",x"2f5e",x"3e98",x"3711",x"abef",x"28a8",x"3bfa",x"3858",x"397c",x"2fd7",x"3e9a",x"3711",x"aa66",x"331a",x"3bca",x"3860",x"397f"),
(x"2fcc",x"3e88",x"3718",x"b420",x"9418",x"3bba",x"3860",x"396a",x"2f89",x"3e8c",x"3713",x"b41f",x"2c3a",x"3bb6",x"385b",x"396e",x"2fe3",x"3e8b",x"3718",x"ab65",x"3528",x"3b8f",x"3862",x"396d"),
(x"2fc7",x"3e7f",x"3715",x"a7ae",x"24ea",x"3bfe",x"3860",x"395f",x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2f8e",x"3e87",x"3714",x"ade0",x"24c2",x"3bf6",x"385c",x"3969"),
(x"2f51",x"3e90",x"3710",x"a856",x"29ab",x"3bfc",x"3858",x"3973",x"2f5e",x"3e98",x"3711",x"abef",x"28a8",x"3bfa",x"3858",x"397c",x"3006",x"3e98",x"3714",x"aa45",x"ab10",x"3bfa",x"3864",x"397c"),
(x"2fc7",x"3e7f",x"3715",x"a7ae",x"24ea",x"3bfe",x"3860",x"395f",x"2fd6",x"3e7d",x"3715",x"28bf",x"2fdb",x"3bef",x"3861",x"395d",x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b"),
(x"2f8e",x"3e87",x"3714",x"bbf3",x"2e23",x"2b27",x"3a11",x"3a5b",x"2f6c",x"3e7b",x"3718",x"b9e5",x"3968",x"0000",x"3a10",x"3a62",x"2f6c",x"3e7b",x"36eb",x"b46a",x"3b91",x"316a",x"3a15",x"3a63"),
(x"2f37",x"3f4a",x"36eb",x"bb71",x"b58a",x"2fc3",x"3b2b",x"3b3a",x"2ed7",x"3f52",x"36eb",x"badb",x"b7e7",x"30ac",x"3b2b",x"3b35",x"2f48",x"3f4b",x"3715",x"bac2",x"b812",x"3146",x"3b26",x"3b3a"),
(x"304f",x"3ee5",x"36eb",x"3ba3",x"b453",x"2fdf",x"3902",x"302b",x"302e",x"3ee0",x"36eb",x"3bf4",x"2d6d",x"ac2c",x"3900",x"3012",x"3033",x"3ee0",x"3715",x"3bf4",x"2da3",x"2b3e",x"38f6",x"3025"),
(x"3048",x"3eed",x"3715",x"3bda",x"2e4f",x"312f",x"38fa",x"305a",x"3054",x"3eed",x"36eb",x"3b7a",x"3531",x"30a8",x"3905",x"304d",x"304f",x"3ee5",x"36eb",x"3ba3",x"b453",x"2fdf",x"3902",x"302b"),
(x"3027",x"3ef4",x"3714",x"3a0a",x"3915",x"3126",x"38fd",x"307d",x"302b",x"3ef6",x"36eb",x"38c7",x"3a49",x"310b",x"3907",x"3079",x"3054",x"3eed",x"36eb",x"3b7a",x"3531",x"30a8",x"3905",x"304d"),
(x"2fca",x"3ef8",x"3714",x"3235",x"3bc0",x"30e0",x"38fe",x"30a4",x"2fcc",x"3efa",x"36eb",x"23ae",x"3bec",x"306c",x"3908",x"30a1",x"302b",x"3ef6",x"36eb",x"38c7",x"3a49",x"310b",x"3907",x"3079"),
(x"2ef2",x"3ef7",x"3714",x"b35f",x"3baf",x"30fd",x"38ff",x"30df",x"2ed8",x"3ef8",x"36eb",x"b6e0",x"3b1c",x"3118",x"3909",x"30e3",x"2fcc",x"3efa",x"36eb",x"23ae",x"3bec",x"306c",x"3908",x"30a1"),
(x"2e86",x"3ef1",x"3715",x"ba37",x"38de",x"311d",x"38fe",x"3104",x"2e6e",x"3ef2",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3909",x"310b",x"2ed8",x"3ef8",x"36eb",x"b6e0",x"3b1c",x"3118",x"3909",x"30e3"),
(x"2e63",x"3eea",x"3715",x"bbf2",x"2495",x"2f43",x"38fd",x"3126",x"2e54",x"3eea",x"36eb",x"bbf7",x"2138",x"2dce",x"3908",x"312d",x"2e6e",x"3ef2",x"36eb",x"bb2d",x"36c9",x"2ff6",x"3909",x"310b"),
(x"2e6b",x"3ee3",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3906",x"314b",x"2e54",x"3eea",x"36eb",x"bbf7",x"2138",x"2dce",x"3908",x"312d",x"2e63",x"3eea",x"3715",x"bbf2",x"2495",x"2f43",x"38fd",x"3126"),
(x"2e93",x"3ede",x"36eb",x"bbfd",x"212b",x"29e6",x"3905",x"3161",x"2e6b",x"3ee3",x"36eb",x"bb9a",x"b4b0",x"2eae",x"3906",x"314b",x"2e80",x"3ee3",x"3715",x"bb87",x"b537",x"2d81",x"38fc",x"3144"),
(x"2e6c",x"3ec4",x"36eb",x"bb9b",x"34d2",x"2ca5",x"3900",x"31ce",x"2e77",x"3ec4",x"3717",x"bbe8",x"30a2",x"2973",x"38f6",x"31c5",x"2e3f",x"3ec2",x"3714",x"bb74",x"35a6",x"2d5e",x"38f6",x"31d7"),
(x"2f22",x"3edf",x"36eb",x"3bf7",x"9e73",x"2dbc",x"38ea",x"2ddb",x"2f13",x"3edf",x"3718",x"3bf1",x"95bc",x"2fb6",x"38ea",x"2e35",x"2f16",x"3ee4",x"3716",x"3bb3",x"33ed",x"2eeb",x"38ef",x"2e30"),
(x"2f2a",x"3ec5",x"36eb",x"3a79",x"3840",x"3401",x"38ce",x"2de0",x"2f0c",x"3ec2",x"3718",x"3a6d",x"3838",x"3468",x"38cb",x"2e3c",x"2f13",x"3edf",x"3718",x"3bf1",x"95bc",x"2fb6",x"38ea",x"2e35"),
(x"306e",x"3ec3",x"3715",x"3bb4",x"33e7",x"2ed7",x"38e9",x"2f58",x"3077",x"3ec4",x"36eb",x"3bc6",x"328d",x"2f71",x"38f3",x"2f37",x"3079",x"3eb9",x"36eb",x"3409",x"bbbc",x"27e2",x"38ee",x"2edd"),
(x"2e24",x"3eb8",x"36eb",x"b6d0",x"bb39",x"2ab1",x"38fd",x"320b",x"2e34",x"3ec3",x"36eb",x"bb76",x"3593",x"2dee",x"3900",x"31de",x"2e3f",x"3ec2",x"3714",x"bb74",x"35a6",x"2d5e",x"38f6",x"31d7"),
(x"2fc8",x"3ee0",x"36eb",x"bbd3",x"b208",x"2da6",x"391d",x"2de9",x"2fc7",x"3ee4",x"36ee",x"bb70",x"358e",x"2fc0",x"3918",x"2ded",x"2fd7",x"3ee3",x"3715",x"bb88",x"3531",x"2dc2",x"3918",x"2e3b"),
(x"2ffa",x"3ee8",x"36ee",x"bb20",x"3725",x"2d51",x"3913",x"2ded",x"3005",x"3ee9",x"3717",x"bbd6",x"323b",x"2a8a",x"3911",x"2e3e",x"2fd7",x"3ee3",x"3715",x"bb88",x"3531",x"2dc2",x"3918",x"2e3b"),
(x"2fff",x"3eec",x"36ee",x"bb1d",x"b747",x"2911",x"390e",x"2dec",x"2fff",x"3eed",x"3716",x"baa5",x"b86c",x"2baa",x"390c",x"2e3b",x"3005",x"3ee9",x"3717",x"bbd6",x"323b",x"2a8a",x"3911",x"2e3e"),
(x"2f00",x"3eec",x"36ee",x"3a67",x"b8c6",x"2a76",x"38f9",x"2de4",x"2ef1",x"3eec",x"3714",x"3b37",x"b6c3",x"2d61",x"38f8",x"2e30",x"2f3a",x"3ef0",x"3715",x"36a0",x"bb47",x"2074",x"38ff",x"2e34"),
(x"2fd9",x"3edf",x"3716",x"bbce",x"b2bb",x"2b41",x"391c",x"2e40",x"301e",x"3ec3",x"3718",x"b98b",x"396b",x"33db",x"393b",x"2e58",x"3016",x"3ec6",x"36eb",x"bbe6",x"2cac",x"3077",x"3939",x"2dfc"),
(x"3033",x"3ee0",x"3715",x"21a1",x"23fc",x"3bff",x"3991",x"32b4",x"2fd9",x"3edf",x"3716",x"282f",x"2808",x"3bfd",x"398c",x"32b2",x"2fd7",x"3ee3",x"3715",x"a8d3",x"a80e",x"3bfd",x"398c",x"32bc"),
(x"303e",x"3ee5",x"3718",x"a8fa",x"a4f7",x"3bfe",x"3992",x"32bf",x"2fd7",x"3ee3",x"3715",x"a8d3",x"a80e",x"3bfd",x"398c",x"32bc",x"3005",x"3ee9",x"3717",x"a511",x"281b",x"3bfe",x"398e",x"32c8"),
(x"3048",x"3eed",x"3715",x"1e8d",x"2bdf",x"3bfc",x"3993",x"32d2",x"3005",x"3ee9",x"3717",x"a511",x"281b",x"3bfe",x"398e",x"32c8",x"2fff",x"3eed",x"3716",x"a52b",x"2c96",x"3bfa",x"398e",x"32d3"),
(x"3027",x"3ef4",x"3714",x"a63f",x"27c1",x"3bfe",x"3990",x"32e3",x"2fff",x"3eed",x"3716",x"a52b",x"2c96",x"3bfa",x"398e",x"32d3",x"2fc2",x"3eef",x"3713",x"991e",x"9cea",x"3c00",x"398b",x"32d8"),
(x"2fca",x"3ef8",x"3714",x"2187",x"a0ea",x"3bff",x"398c",x"32ed",x"2fc2",x"3eef",x"3713",x"991e",x"9cea",x"3c00",x"398b",x"32d8",x"2f3a",x"3ef0",x"3715",x"1c81",x"1953",x"3c00",x"3987",x"32d9"),
(x"2ef2",x"3ef7",x"3714",x"9dd6",x"248e",x"3bff",x"3984",x"32ea",x"2f3a",x"3ef0",x"3715",x"1c81",x"1953",x"3c00",x"3987",x"32d9",x"2ef1",x"3eec",x"3714",x"1da1",x"252b",x"3bff",x"3984",x"32cf"),
(x"2ef1",x"3eec",x"3714",x"1da1",x"252b",x"3bff",x"3984",x"32cf",x"2eed",x"3ee8",x"3716",x"a338",x"267a",x"3bff",x"3984",x"32c7",x"2e63",x"3eea",x"3715",x"1818",x"26bb",x"3bff",x"397f",x"32ca"),
(x"2eed",x"3ee8",x"3716",x"a338",x"267a",x"3bff",x"3984",x"32c7",x"2f16",x"3ee4",x"3716",x"a4bc",x"2b17",x"3bfc",x"3985",x"32bd",x"2e80",x"3ee3",x"3715",x"a645",x"29e0",x"3bfd",x"3980",x"32ba"),
(x"2e80",x"3ee3",x"3715",x"a645",x"29e0",x"3bfd",x"3980",x"32ba",x"2f16",x"3ee4",x"3716",x"a4bc",x"2b17",x"3bfc",x"3985",x"32bd",x"2f13",x"3edf",x"3718",x"a793",x"243f",x"3bfe",x"3985",x"32b2"),
(x"2e77",x"3ec4",x"3717",x"a984",x"a0c2",x"3bfd",x"3980",x"3272",x"2e96",x"3ede",x"3717",x"a7d5",x"236c",x"3bfe",x"3981",x"32af",x"2f13",x"3edf",x"3718",x"a793",x"243f",x"3bfe",x"3985",x"32b2"),
(x"2efa",x"3ee8",x"36ee",x"3b84",x"3534",x"2e9f",x"38f5",x"2de3",x"2eed",x"3ee8",x"3716",x"3ba1",x"34a7",x"2cd8",x"38f4",x"2e32",x"2ef1",x"3eec",x"3714",x"3b37",x"b6c3",x"2d61",x"38f8",x"2e30"),
(x"3033",x"3ee0",x"3715",x"3bf4",x"2da3",x"2b3e",x"38f6",x"3025",x"302e",x"3ee0",x"36eb",x"3bf4",x"2d6d",x"ac2c",x"3900",x"3012",x"3065",x"3ec5",x"36eb",x"3baa",x"3479",x"2b93",x"38f4",x"2f49"),
(x"306e",x"3ec3",x"3715",x"3bb4",x"33e7",x"2ed7",x"38e9",x"2f58",x"3056",x"3ec4",x"3718",x"3ba4",x"33dc",x"313e",x"38e9",x"2f72",x"3065",x"3ec5",x"36eb",x"3baa",x"3479",x"2b93",x"38f4",x"2f49"),
(x"2f0c",x"3ec2",x"3718",x"a3ae",x"ac2f",x"3bfb",x"3985",x"326e",x"301e",x"3ec3",x"3718",x"224c",x"a36c",x"3bff",x"3990",x"326f",x"3072",x"3eb8",x"3715",x"2081",x"ad9e",x"3bf8",x"3996",x"3257"),
(x"2fff",x"3eec",x"36ee",x"bb1d",x"b747",x"2911",x"390e",x"2dec",x"2fc4",x"3ef0",x"36ee",x"b52c",x"bb8d",x"ac0b",x"3908",x"2de8",x"2fc2",x"3eef",x"3713",x"b46c",x"bbaf",x"a5f6",x"3908",x"2e32"),
(x"2e77",x"3ec4",x"3717",x"bbe8",x"30a2",x"2973",x"38f6",x"31c5",x"2e6c",x"3ec4",x"36eb",x"bb9b",x"34d2",x"2ca5",x"3900",x"31ce",x"2e93",x"3ede",x"36eb",x"bbfd",x"212b",x"29e6",x"3905",x"3161"),
(x"2f3e",x"3ef0",x"36ee",x"314a",x"bbe2",x"a87e",x"38ff",x"2de6",x"2f3a",x"3ef0",x"3715",x"36a0",x"bb47",x"2074",x"38ff",x"2e34",x"2fc2",x"3eef",x"3713",x"b46c",x"bbaf",x"a5f6",x"3908",x"2e32"),
(x"2f2a",x"3ec5",x"36eb",x"3a79",x"3840",x"3401",x"3949",x"2dd9",x"3016",x"3ec6",x"36eb",x"bbe6",x"2cac",x"3077",x"3939",x"2dfc",x"301e",x"3ec3",x"3718",x"b98b",x"396b",x"33db",x"393b",x"2e58"),
(x"2e32",x"3eb9",x"3714",x"af03",x"bbf3",x"23ef",x"38f4",x"31ff",x"3072",x"3eb8",x"3715",x"33c8",x"bbc2",x"236c",x"38e5",x"32ad",x"3079",x"3eb9",x"36eb",x"3409",x"bbbc",x"27e2",x"38ee",x"32c0"),
(x"2efa",x"3ee8",x"36ee",x"3b84",x"3534",x"2e9f",x"38f5",x"2de3",x"2f2c",x"3ee5",x"36eb",x"3ba6",x"341e",x"3066",x"38ef",x"2dd9",x"2f16",x"3ee4",x"3716",x"3bb3",x"33ed",x"2eeb",x"38ef",x"2e30"),
(x"2f10",x"3fcc",x"370e",x"afd2",x"2717",x"3bef",x"3b82",x"3baf",x"2f7a",x"3fd4",x"3712",x"b42b",x"2e69",x"3bae",x"3b86",x"3bb7",x"2fbb",x"3fd4",x"3716",x"b0f9",x"a8af",x"3be5",x"3b89",x"3bb7"),
(x"2fbb",x"3fd4",x"3716",x"3add",x"375a",x"334d",x"3b5c",x"388d",x"2fd0",x"3fd7",x"36eb",x"3996",x"395e",x"33ec",x"3b61",x"388e",x"301b",x"3fc7",x"36eb",x"3b99",x"3315",x"330d",x"3b61",x"3885"),
(x"2fb0",x"3f87",x"3714",x"2c39",x"29a5",x"3bf9",x"3b8e",x"3b77",x"2fe3",x"3f8f",x"3713",x"2da3",x"2f15",x"3beb",x"3b90",x"3b7e",x"3001",x"3f8f",x"3712",x"2a69",x"287e",x"3bfc",x"3b91",x"3b7e"),
(x"3017",x"3f91",x"3711",x"2994",x"2977",x"3bfc",x"3b93",x"3b80",x"3038",x"3f91",x"3712",x"aa38",x"ad35",x"3bf6",x"3b96",x"3b80",x"304c",x"3f8d",x"3711",x"2481",x"254c",x"3bff",x"3b98",x"3b7c"),
(x"303e",x"3f87",x"3712",x"2a73",x"2a97",x"3bfa",x"3b97",x"3b78",x"301b",x"3f85",x"3713",x"291b",x"2b55",x"3bfb",x"3b94",x"3b76",x"3001",x"3f8f",x"3712",x"2a69",x"287e",x"3bfc",x"3b91",x"3b7e"),
(x"2ff2",x"3f82",x"3718",x"2e36",x"a160",x"3bf6",x"3b91",x"3b74",x"300c",x"3f84",x"3716",x"2f15",x"329c",x"3bc6",x"3b93",x"3b75",x"302f",x"3f81",x"3711",x"2fec",x"ac2c",x"3beb",x"3b96",x"3b73"),
(x"301b",x"3f6a",x"3713",x"2e9a",x"3366",x"3bbd",x"3b96",x"3b5f",x"2ff0",x"3f6f",x"370f",x"ab8a",x"30af",x"3be6",x"3b92",x"3b63",x"2ff4",x"3f71",x"370e",x"a6d5",x"25c2",x"3bfe",x"3b92",x"3b65"),
(x"3013",x"3f76",x"3713",x"2538",x"ac79",x"3bfa",x"3b94",x"3b69",x"305c",x"3f70",x"370f",x"2cd8",x"a71d",x"3bf9",x"3b9c",x"3b65",x"3040",x"3f6b",x"370f",x"1df0",x"a631",x"3bff",x"3b99",x"3b61"),
(x"3013",x"3f76",x"3713",x"2538",x"ac79",x"3bfa",x"3b94",x"3b69",x"3014",x"3f78",x"3713",x"27e9",x"284d",x"3bfd",x"3b94",x"3b6b",x"3058",x"3f79",x"370f",x"2ec5",x"19f0",x"3bf4",x"3b9b",x"3b6d"),
(x"302f",x"3f81",x"3711",x"2fec",x"ac2c",x"3beb",x"3b96",x"3b73",x"3058",x"3f79",x"370f",x"2ec5",x"19f0",x"3bf4",x"3b9b",x"3b6d",x"3014",x"3f78",x"3713",x"27e9",x"284d",x"3bfd",x"3b94",x"3b6b"),
(x"3000",x"3f7a",x"3710",x"2c5b",x"b0a4",x"3be5",x"3b92",x"3b6d",x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70",x"302f",x"3f81",x"3711",x"2fec",x"ac2c",x"3beb",x"3b96",x"3b73"),
(x"3000",x"3f7a",x"3710",x"2c5b",x"b0a4",x"3be5",x"3b92",x"3b6d",x"2fc1",x"3f7b",x"3713",x"a5b5",x"b7de",x"3af6",x"3b8f",x"3b6e",x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70"),
(x"2f48",x"3f4b",x"3715",x"26c2",x"ac63",x"3bfa",x"3b89",x"3b45",x"2f5a",x"3f53",x"3717",x"17c8",x"9f79",x"3c00",x"3b8a",x"3b4d",x"2f7f",x"3f52",x"3717",x"2ff2",x"aa7d",x"3bed",x"3b8c",x"3b4c"),
(x"302b",x"3f5b",x"3716",x"2cd8",x"a7e2",x"3bf9",x"3b96",x"3b53",x"3045",x"3f59",x"3714",x"285d",x"af8b",x"3bf0",x"3b98",x"3b51",x"3050",x"3f55",x"3712",x"3163",x"a345",x"3be2",x"3b99",x"3b4e"),
(x"3044",x"3f51",x"3714",x"9553",x"ab62",x"3bfc",x"3b98",x"3b4b",x"3000",x"3f4e",x"3711",x"a40b",x"ad5c",x"3bf8",x"3b92",x"3b48",x"300a",x"3f5a",x"3716",x"a818",x"ad04",x"3bf8",x"3b93",x"3b52"),
(x"2fa9",x"3f54",x"3714",x"3036",x"a73e",x"3bed",x"3b8e",x"3b4d",x"2fd3",x"3f57",x"3714",x"2504",x"ada9",x"3bf7",x"3b90",x"3b50",x"3000",x"3f4e",x"3711",x"a40b",x"ad5c",x"3bf8",x"3b92",x"3b48"),
(x"2fe3",x"3f4c",x"3711",x"327d",x"175f",x"3bd5",x"3b90",x"3b47",x"2f7f",x"3f52",x"3717",x"2ff2",x"aa7d",x"3bed",x"3b8c",x"3b4c",x"2fa9",x"3f54",x"3714",x"3036",x"a73e",x"3bed",x"3b8e",x"3b4d"),
(x"2fe3",x"3f4c",x"3711",x"327d",x"175f",x"3bd5",x"3b90",x"3b47",x"2fd7",x"3f4b",x"3712",x"2f67",x"a981",x"3bf0",x"3b90",x"3b46",x"2f7f",x"3f52",x"3717",x"2ff2",x"aa7d",x"3bed",x"3b8c",x"3b4c"),
(x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34",x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2fe6",x"3f45",x"3712",x"3146",x"2c91",x"3bde",x"3b91",x"3b41"),
(x"2f3d",x"3f39",x"3718",x"a138",x"ae95",x"3bf4",x"3b89",x"3b37",x"2f4b",x"3f34",x"3715",x"a8bf",x"afdb",x"3bef",x"3b8a",x"3b33",x"2ef3",x"3f38",x"3719",x"290e",x"af00",x"3bf2",x"3b85",x"3b37"),
(x"2f49",x"3f3a",x"3718",x"ab4f",x"2525",x"3bfc",x"3b89",x"3b38",x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2fb5",x"3f36",x"3718",x"2e3b",x"1fae",x"3bf6",x"3b8e",x"3b34"),
(x"2f49",x"3f3a",x"3718",x"ab4f",x"2525",x"3bfc",x"3b89",x"3b38",x"2f16",x"3f3e",x"3715",x"ad65",x"ac5a",x"3bf3",x"3b87",x"3b3b",x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e"),
(x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2f16",x"3f3e",x"3715",x"ad65",x"ac5a",x"3bf3",x"3b87",x"3b3b",x"2ede",x"3f43",x"3718",x"acf2",x"18ea",x"3bf9",x"3b84",x"3b3f"),
(x"2ed4",x"3f47",x"3712",x"b59c",x"336a",x"3b42",x"3b83",x"3b42",x"2ee4",x"3f49",x"3712",x"b541",x"30b9",x"3b76",x"3b84",x"3b44",x"2f1d",x"3f49",x"3717",x"ad2d",x"2ecb",x"3bed",x"3b87",x"3b44"),
(x"2f73",x"3f42",x"3718",x"2bb4",x"28d3",x"3bfa",x"3b8b",x"3b3e",x"2f1d",x"3f49",x"3717",x"ad2d",x"2ecb",x"3bed",x"3b87",x"3b44",x"2f3a",x"3f49",x"3716",x"300a",x"2da8",x"3be7",x"3b89",x"3b44"),
(x"2fd7",x"3f4b",x"3712",x"2f67",x"a981",x"3bf0",x"3b90",x"3b46",x"2fe6",x"3f45",x"3712",x"3146",x"2c91",x"3bde",x"3b91",x"3b41",x"2f3a",x"3f49",x"3716",x"300a",x"2da8",x"3be7",x"3b89",x"3b44"),
(x"2f5a",x"3f53",x"3717",x"17c8",x"9f79",x"3c00",x"3b8a",x"3b4d",x"2f06",x"3f51",x"3718",x"2c00",x"290e",x"3bfa",x"3b86",x"3b4a",x"2f11",x"3f58",x"3715",x"251e",x"2d06",x"3bf9",x"3b86",x"3b51"),
(x"2f5a",x"3f53",x"3717",x"17c8",x"9f79",x"3c00",x"3b8a",x"3b4d",x"2f3c",x"3f4d",x"3714",x"257a",x"ae8a",x"3bf4",x"3b89",x"3b47",x"2f06",x"3f51",x"3718",x"2c00",x"290e",x"3bfa",x"3b86",x"3b4a"),
(x"2f11",x"3f58",x"3715",x"251e",x"2d06",x"3bf9",x"3b86",x"3b51",x"2f06",x"3f51",x"3718",x"2c00",x"290e",x"3bfa",x"3b86",x"3b4a",x"2e9f",x"3f5d",x"3714",x"975f",x"2c2c",x"3bfb",x"3b81",x"3b54"),
(x"2ece",x"3f60",x"3714",x"adba",x"2266",x"3bf7",x"3b83",x"3b57",x"2e9f",x"3f5d",x"3714",x"975f",x"2c2c",x"3bfb",x"3b81",x"3b54",x"2e7c",x"3f69",x"3712",x"b106",x"273e",x"3be5",x"3b80",x"3b5f"),
(x"2ec2",x"3f6b",x"3715",x"b468",x"247a",x"3bb0",x"3b83",x"3b60",x"2e7c",x"3f69",x"3712",x"b106",x"273e",x"3be5",x"3b80",x"3b5f",x"2ea0",x"3f75",x"3710",x"b550",x"2e33",x"3b81",x"3b81",x"3b68"),
(x"2ed8",x"3f73",x"3717",x"b273",x"2f43",x"3bc8",x"3b84",x"3b66",x"2ea0",x"3f75",x"3710",x"b550",x"2e33",x"3b81",x"3b81",x"3b68",x"2ef8",x"3f7d",x"3712",x"ab5c",x"2345",x"3bfc",x"3b85",x"3b6e"),
(x"2f7e",x"3f7b",x"3712",x"add2",x"b04b",x"3be4",x"3b8c",x"3b6d",x"2fad",x"3f83",x"3716",x"af4b",x"aa5f",x"3bf0",x"3b8e",x"3b74",x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70"),
(x"2f7e",x"3f7b",x"3712",x"add2",x"b04b",x"3be4",x"3b8c",x"3b6d",x"2ef8",x"3f7d",x"3712",x"ab5c",x"2345",x"3bfc",x"3b85",x"3b6e",x"2fad",x"3f83",x"3716",x"af4b",x"aa5f",x"3bf0",x"3b8e",x"3b74"),
(x"2f7e",x"3f7b",x"3712",x"add2",x"b04b",x"3be4",x"3b8c",x"3b6d",x"2f3c",x"3f7a",x"3711",x"2e24",x"2a2b",x"3bf4",x"3b89",x"3b6c",x"2ef8",x"3f7d",x"3712",x"ab5c",x"2345",x"3bfc",x"3b85",x"3b6e"),
(x"2ff2",x"3f82",x"3718",x"2e36",x"a160",x"3bf6",x"3b91",x"3b74",x"2fbb",x"3f7e",x"3718",x"2c13",x"b1c5",x"3bda",x"3b8f",x"3b70",x"2fad",x"3f83",x"3716",x"af4b",x"aa5f",x"3bf0",x"3b8e",x"3b74"),
(x"300c",x"3f84",x"3716",x"2f15",x"329c",x"3bc6",x"3b93",x"3b75",x"2fb0",x"3f87",x"3714",x"2c39",x"29a5",x"3bf9",x"3b8e",x"3b77",x"301b",x"3f85",x"3713",x"291b",x"2b55",x"3bfb",x"3b94",x"3b76"),
(x"300c",x"3f84",x"3716",x"2f15",x"329c",x"3bc6",x"3b93",x"3b75",x"2fc5",x"3f84",x"3716",x"2553",x"32c7",x"3bd1",x"3b8f",x"3b75",x"2fb0",x"3f87",x"3714",x"2c39",x"29a5",x"3bf9",x"3b8e",x"3b77"),
(x"2fe3",x"3f8f",x"3713",x"2da3",x"2f15",x"3beb",x"3b90",x"3b7e",x"2fb0",x"3f87",x"3714",x"2c39",x"29a5",x"3bf9",x"3b8e",x"3b77",x"2f3b",x"3f8e",x"3717",x"30e7",x"3057",x"3bd4",x"3b88",x"3b7d"),
(x"2f8e",x"3f93",x"370f",x"2edc",x"2cd0",x"3bee",x"3b8c",x"3b81",x"2f3b",x"3f8e",x"3717",x"30e7",x"3057",x"3bd4",x"3b88",x"3b7d",x"2eeb",x"3f9c",x"3713",x"29b8",x"a6e2",x"3bfd",x"3b83",x"3b88"),
(x"2ecd",x"3fb8",x"370d",x"b809",x"2e09",x"3add",x"3b80",x"3b9f",x"2ee7",x"3fba",x"3713",x"af9f",x"b907",x"3a26",x"3b81",x"3ba1",x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1"),
(x"3007",x"3fc7",x"3715",x"ad56",x"20d0",x"3bf8",x"3b8e",x"3bac",x"2ffb",x"3fba",x"3715",x"99f0",x"a6cf",x"3bff",x"3b8e",x"3ba2",x"2efa",x"3fc1",x"3712",x"a9f0",x"2b1d",x"3bfa",x"3b81",x"3ba6"),
(x"300f",x"3fb9",x"36eb",x"3b89",x"b473",x"31fc",x"3b60",x"387e",x"2f92",x"3fa7",x"36eb",x"3b4a",x"b677",x"2cfa",x"3b5e",x"3874",x"2f8b",x"3fa8",x"370e",x"3b5f",x"b5f1",x"2f4f",x"3b5a",x"3875"),
(x"3029",x"3f23",x"36eb",x"bba1",x"b4cc",x"1f45",x"3b8d",x"3a14",x"3024",x"3f23",x"3713",x"bba5",x"b497",x"ac28",x"3b92",x"3a14",x"302f",x"3f1a",x"3710",x"bbfd",x"a997",x"a09b",x"3b92",x"3a0f"),
(x"302f",x"3f1a",x"3710",x"bbfd",x"a997",x"a09b",x"3b92",x"3a0f",x"302e",x"3f14",x"36eb",x"bbf5",x"2e59",x"2467",x"3b8d",x"3a0c",x"3029",x"3f23",x"36eb",x"bba1",x"b4cc",x"1f45",x"3b8d",x"3a14"),
(x"2fb5",x"3f36",x"36eb",x"346a",x"bb91",x"316a",x"3b8d",x"3a1f",x"2fb5",x"3f36",x"3718",x"39e5",x"b968",x"0000",x"3b92",x"3a1f",x"2ff3",x"3f30",x"3714",x"bb1c",x"b754",x"223f",x"3b92",x"3a1b"),
(x"2ff3",x"3f30",x"3714",x"bb1c",x"b754",x"223f",x"3b92",x"3a1b",x"3029",x"3f23",x"36eb",x"bba1",x"b4cc",x"1f45",x"3b8d",x"3a14",x"2fb5",x"3f36",x"36eb",x"346a",x"bb91",x"316a",x"3b8d",x"3a1f"),
(x"302e",x"3f14",x"36eb",x"bbf5",x"2e59",x"2467",x"3b8d",x"3a0c",x"302b",x"3f12",x"3714",x"bbeb",x"308b",x"98b5",x"3b92",x"3a0b",x"3021",x"3f0e",x"3712",x"bb76",x"35c5",x"204d",x"3b92",x"3a09"),
(x"3021",x"3f0e",x"3712",x"bb76",x"35c5",x"204d",x"3b92",x"3a09",x"301c",x"3f0c",x"36eb",x"bab1",x"3862",x"21f0",x"3b8d",x"3a08",x"302e",x"3f14",x"36eb",x"bbf5",x"2e59",x"2467",x"3b8d",x"3a0c"),
(x"2fe9",x"3f08",x"36eb",x"b7e1",x"3af5",x"269a",x"3b8d",x"3a05",x"301c",x"3f0c",x"36eb",x"bab1",x"3862",x"21f0",x"3b8d",x"3a08",x"300e",x"3f0b",x"3714",x"b95a",x"39f1",x"2032",x"3b92",x"3a07"),
(x"2f83",x"3f07",x"36eb",x"b03c",x"3beb",x"299e",x"3b8d",x"3a01",x"2fe9",x"3f08",x"36eb",x"b7e1",x"3af5",x"269a",x"3b8d",x"3a05",x"2fe4",x"3f08",x"3714",x"b5bf",x"3b76",x"27db",x"3b92",x"3a05"),
(x"2f1b",x"3f08",x"36eb",x"3868",x"3aab",x"296a",x"3b8d",x"39fe",x"2f83",x"3f07",x"36eb",x"b03c",x"3beb",x"299e",x"3b8d",x"3a01",x"2f7e",x"3f06",x"3715",x"2836",x"3bfd",x"294c",x"3b92",x"3a01"),
(x"2ec8",x"3f0e",x"3714",x"3b01",x"37b5",x"2839",x"3b92",x"39f9",x"2ecf",x"3f0e",x"36eb",x"3af3",x"37df",x"2b38",x"3b8d",x"39fa",x"2f1b",x"3f08",x"36eb",x"3868",x"3aab",x"296a",x"3b8d",x"39fe"),
(x"2eb5",x"3f13",x"36eb",x"3bf9",x"2d11",x"2511",x"3b8d",x"39f7",x"2ecf",x"3f0e",x"36eb",x"3af3",x"37df",x"2b38",x"3b8d",x"39fa",x"2ec8",x"3f0e",x"3714",x"3b01",x"37b5",x"2839",x"3b92",x"39f9"),
(x"2ecf",x"3f18",x"36eb",x"390c",x"ba34",x"2532",x"3b8d",x"39f4",x"2eb5",x"3f13",x"36eb",x"3bf9",x"2d11",x"2511",x"3b8d",x"39f7",x"2eb5",x"3f13",x"3714",x"3be6",x"b10f",x"9bfc",x"3b92",x"39f6"),
(x"2f14",x"3f18",x"3714",x"afe2",x"bbee",x"28fd",x"3b8d",x"3650",x"2f19",x"3f18",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3b92",x"364f",x"2ecf",x"3f18",x"36eb",x"390c",x"ba34",x"2532",x"3b92",x"364a"),
(x"2f4a",x"3f16",x"3711",x"b64f",x"bb52",x"2d1b",x"3b8e",x"3654",x"2f44",x"3f15",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3b93",x"3652",x"2f19",x"3f18",x"36eb",x"b5dd",x"bb6d",x"2be9",x"3b92",x"364f"),
(x"2f9f",x"3f25",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b93",x"366c",x"2fb1",x"3f23",x"36eb",x"39db",x"396c",x"2c1a",x"3b93",x"366a",x"2faf",x"3f23",x"3711",x"3a7a",x"38af",x"283c",x"3b8e",x"3669"),
(x"2f9c",x"3f16",x"3710",x"3416",x"bbad",x"2f8d",x"3b8f",x"365a",x"2fa8",x"3f15",x"36eb",x"337e",x"bbba",x"2ef6",x"3b93",x"3659",x"2f44",x"3f15",x"36eb",x"b2b2",x"bbc8",x"2e54",x"3b93",x"3652"),
(x"3013",x"3f68",x"36eb",x"b5e4",x"bb4d",x"31a2",x"3b48",x"3847",x"2fdc",x"3f6e",x"36eb",x"bb7d",x"b521",x"3095",x"3b45",x"3846",x"2ff0",x"3f6f",x"370f",x"ba9c",x"b854",x"30fa",x"3b44",x"384a"),
(x"3007",x"3fc7",x"3715",x"3bc5",x"2b9a",x"3358",x"3b5c",x"3886",x"301b",x"3fc7",x"36eb",x"3b99",x"3315",x"330d",x"3b61",x"3885",x"300f",x"3fb9",x"36eb",x"3b89",x"b473",x"31fc",x"3b60",x"387e"),
(x"2fd1",x"3f20",x"3710",x"2856",x"a9ab",x"3bfc",x"3b90",x"3b23",x"2ec0",x"3f22",x"3711",x"28d9",x"a52b",x"3bfe",x"3b83",x"3b24",x"2f3e",x"3f25",x"3718",x"2b65",x"b528",x"3b8f",x"3b89",x"3b27"),
(x"2f0d",x"3fbb",x"36eb",x"bbe3",x"2ce7",x"30c3",x"3b59",x"389f",x"2efa",x"3fc1",x"3712",x"bbcf",x"b081",x"3141",x"3b57",x"3899",x"2f14",x"3fbc",x"3715",x"bbd7",x"b1f9",x"2c2a",x"3b55",x"389b"),
(x"2f0d",x"3fbb",x"36eb",x"bbe3",x"2ce7",x"30c3",x"3b59",x"389f",x"2edb",x"3fc1",x"36eb",x"bbdb",x"1c67",x"320a",x"3b5b",x"389c",x"2efa",x"3fc1",x"3712",x"bbcf",x"b081",x"3141",x"3b57",x"3899"),
(x"2ea0",x"3f75",x"3710",x"bb6a",x"35bb",x"2efe",x"3b27",x"3b21",x"2e95",x"3f76",x"36eb",x"bb75",x"35a2",x"2d46",x"3b2b",x"3b21",x"2ee2",x"3f7e",x"36eb",x"b958",x"39de",x"2fe4",x"3b2b",x"3b1c"),
(x"2fd3",x"3f18",x"36eb",x"3aa4",x"b859",x"2fe5",x"3b93",x"365d",x"2fa8",x"3f15",x"36eb",x"337e",x"bbba",x"2ef6",x"3b93",x"3659",x"2f9c",x"3f16",x"3710",x"3416",x"bbad",x"2f8d",x"3b8f",x"365a"),
(x"2f4a",x"3f28",x"36eb",x"bbe6",x"308f",x"2c41",x"3b28",x"3b68",x"2f4e",x"3f31",x"36eb",x"bbfa",x"a0a8",x"2cba",x"3b26",x"3b64",x"2f5a",x"3f31",x"3715",x"bbfa",x"a710",x"2c48",x"3b21",x"3b65"),
(x"2fdc",x"3f1c",x"3710",x"3bcc",x"b228",x"2f2f",x"3b8f",x"3661",x"2fec",x"3f1c",x"36eb",x"3bf4",x"9edc",x"2eb6",x"3b93",x"3662",x"2fd3",x"3f18",x"36eb",x"3aa4",x"b859",x"2fe5",x"3b93",x"365d"),
(x"2fdc",x"3f6e",x"36eb",x"bb7d",x"b521",x"3095",x"3b45",x"3846",x"2fe5",x"3f71",x"36eb",x"bb19",x"3744",x"2cf7",x"3b44",x"3845",x"2ff4",x"3f71",x"370e",x"bb25",x"370e",x"2d6a",x"3b42",x"384a"),
(x"3048",x"3f4f",x"36eb",x"36fe",x"bb25",x"2ea4",x"39fa",x"3b7b",x"2ff6",x"3f4d",x"36eb",x"37d8",x"baf6",x"2a35",x"39f9",x"3b76",x"3000",x"3f4e",x"3711",x"34dc",x"bb97",x"2d61",x"39f4",x"3b78"),
(x"2fb1",x"3f23",x"36eb",x"39db",x"396c",x"2c1a",x"3b93",x"366a",x"2fe0",x"3f21",x"36eb",x"3b02",x"3776",x"2fc8",x"3b93",x"3666",x"2fd1",x"3f20",x"3710",x"3b2f",x"36d9",x"2e52",x"3b8f",x"3666"),
(x"2ef8",x"3f7d",x"3712",x"b84e",x"3ab0",x"2ec7",x"3b26",x"3b1d",x"2ee2",x"3f7e",x"36eb",x"b958",x"39de",x"2fe4",x"3b2b",x"3b1c",x"2fb4",x"3f84",x"36eb",x"b776",x"3b0b",x"2d41",x"3b2a",x"3b15"),
(x"2f5a",x"3f31",x"3715",x"bbfa",x"a710",x"2c48",x"3b21",x"3b65",x"2f4e",x"3f31",x"36eb",x"bbfa",x"a0a8",x"2cba",x"3b26",x"3b64",x"2f48",x"3f33",x"36eb",x"b9df",x"b964",x"2d28",x"3b26",x"3b63"),
(x"2ff4",x"3f71",x"370e",x"bb25",x"370e",x"2d6a",x"3b42",x"384a",x"2fe5",x"3f71",x"36eb",x"bb19",x"3744",x"2cf7",x"3b44",x"3845",x"300f",x"3f76",x"36eb",x"bad3",x"3822",x"2c4d",x"3b41",x"3845"),
(x"2f8b",x"3fa8",x"370e",x"3b5f",x"b5f1",x"2f4f",x"3b5a",x"3875",x"2f92",x"3fa7",x"36eb",x"3b4a",x"b677",x"2cfa",x"3b5e",x"3874",x"2f5b",x"3f9d",x"36eb",x"3bfe",x"1e8d",x"2828",x"3b5c",x"386e"),
(x"2fb4",x"3f84",x"36eb",x"b776",x"3b0b",x"2d41",x"3b2a",x"3b15",x"2fc0",x"3f84",x"36eb",x"bb23",x"b71d",x"2cde",x"3b2a",x"3b14",x"2fc5",x"3f84",x"3716",x"bbde",x"31b5",x"2825",x"3b25",x"3b15"),
(x"2f4b",x"3f34",x"3715",x"b95d",x"b9e3",x"2de3",x"3b21",x"3b64",x"2f48",x"3f33",x"36eb",x"b9df",x"b964",x"2d28",x"3b26",x"3b63",x"2ed5",x"3f38",x"36eb",x"b9ed",x"b94b",x"2f45",x"3b25",x"3b5e"),
(x"2fe5",x"3f4a",x"36eb",x"3bf8",x"a379",x"2d44",x"3b23",x"3bb2",x"2fd7",x"3f4b",x"3712",x"3bf7",x"283f",x"2d8f",x"3b1e",x"3bb1",x"2fe3",x"3f4c",x"3711",x"3b12",x"b762",x"2ca3",x"3b1e",x"3bb2"),
(x"2fe3",x"3f4c",x"3711",x"3b12",x"b762",x"2ca3",x"3b1e",x"3bb2",x"2ff6",x"3f4d",x"36eb",x"37d8",x"baf6",x"2a35",x"3b23",x"3bb4",x"2fe5",x"3f4a",x"36eb",x"3bf8",x"a379",x"2d44",x"3b23",x"3bb2"),
(x"3013",x"3f76",x"3713",x"bb5b",x"3634",x"2c08",x"3b40",x"384a",x"300f",x"3f76",x"36eb",x"bad3",x"3822",x"2c4d",x"3b41",x"3845",x"3010",x"3f77",x"36eb",x"b9e9",x"b955",x"2e31",x"3b40",x"3844"),
(x"2f5b",x"3f9d",x"36eb",x"3bfe",x"1e8d",x"2828",x"3b5c",x"386e",x"2f92",x"3f94",x"36eb",x"3ab4",x"3859",x"2a59",x"3b5b",x"3869",x"2f8e",x"3f93",x"370f",x"3ad7",x"3821",x"29e3",x"3b57",x"386a"),
(x"2fc0",x"3f84",x"36eb",x"bb23",x"b71d",x"2cde",x"3b42",x"38b6",x"2f9f",x"3f86",x"36eb",x"b97a",x"b9b6",x"3099",x"3b43",x"38b5",x"2fb0",x"3f87",x"3714",x"b9e8",x"b951",x"2f27",x"3b40",x"38b0"),
(x"2ed5",x"3f38",x"36eb",x"b9ed",x"b94b",x"2f45",x"3b25",x"3b5e",x"2edf",x"3f3b",x"36eb",x"b2cb",x"3bc1",x"2fc5",x"3b24",x"3b5d",x"2ef4",x"3f39",x"3719",x"b251",x"3bca",x"2f22",x"3b1f",x"3b60"),
(x"2fe5",x"3f4a",x"36eb",x"3bf8",x"a379",x"2d44",x"3b23",x"3bb2",x"2fee",x"3f46",x"36eb",x"3b57",x"3625",x"2e99",x"3b24",x"3bb0",x"2fe6",x"3f45",x"3712",x"3b92",x"3509",x"2cb4",x"3b1f",x"3bae"),
(x"2fb8",x"3f7b",x"36eb",x"b046",x"bbe8",x"2cb7",x"39fa",x"3ba8",x"2fc1",x"3f7b",x"3713",x"b0a8",x"bbea",x"22cf",x"39f5",x"3ba9",x"3000",x"3f7a",x"3710",x"b833",x"bac7",x"2d1d",x"39f6",x"3bab"),
(x"3000",x"3f7a",x"3710",x"b833",x"bac7",x"2d1d",x"39f6",x"3bab",x"3010",x"3f77",x"36eb",x"b9e9",x"b955",x"2e31",x"39fb",x"3bac",x"2fb8",x"3f7b",x"36eb",x"b046",x"bbe8",x"2cb7",x"39fa",x"3ba8"),
(x"2f8e",x"3f93",x"370f",x"3ad7",x"3821",x"29e3",x"3b57",x"386a",x"2f92",x"3f94",x"36eb",x"3ab4",x"3859",x"2a59",x"3b5b",x"3869",x"2fee",x"3f8f",x"36eb",x"373f",x"3b1a",x"2d3c",x"3b5b",x"3865"),
(x"2f9f",x"3f86",x"36eb",x"b97a",x"b9b6",x"3099",x"3b43",x"38b5",x"2f20",x"3f8e",x"36eb",x"baff",x"b73c",x"3197",x"3b47",x"38b2",x"2f3b",x"3f8e",x"3717",x"ba77",x"b889",x"310c",x"3b44",x"38ad"),
(x"2ef4",x"3f39",x"3719",x"b251",x"3bca",x"2f22",x"3b1f",x"3b60",x"2edf",x"3f3b",x"36eb",x"b2cb",x"3bc1",x"2fc5",x"3b24",x"3b5d",x"2f48",x"3f3a",x"36eb",x"bb01",x"3745",x"3141",x"3b22",x"3b5a"),
(x"2fee",x"3f46",x"36eb",x"3b57",x"3625",x"2e99",x"3b24",x"3bb0",x"303d",x"3f33",x"36eb",x"3b99",x"345f",x"30d6",x"3b27",x"3ba6",x"302e",x"3f34",x"3711",x"3b70",x"3585",x"3014",x"3b22",x"3ba5"),
(x"2f42",x"3f79",x"36eb",x"374a",x"bb15",x"2de4",x"39fa",x"3ba4",x"2f3c",x"3f7a",x"3711",x"3934",x"ba0d",x"2c18",x"39f5",x"3ba5",x"2f7e",x"3f7b",x"3712",x"32e8",x"bbcb",x"2c10",x"39f5",x"3ba7"),
(x"2f7e",x"3f7b",x"3712",x"32e8",x"bbcb",x"2c10",x"39f5",x"3ba7",x"2fb8",x"3f7b",x"36eb",x"b046",x"bbe8",x"2cb7",x"39fa",x"3ba8",x"2f42",x"3f79",x"36eb",x"374a",x"bb15",x"2de4",x"39fa",x"3ba4"),
(x"2fee",x"3f8f",x"36eb",x"373f",x"3b1a",x"2d3c",x"3b5b",x"3865",x"3004",x"3f90",x"36eb",x"b8ae",x"3a73",x"2d47",x"3b5b",x"3864",x"3001",x"3f8f",x"3712",x"b721",x"3b24",x"2bf2",x"3b56",x"3865"),
(x"2f20",x"3f8e",x"36eb",x"baff",x"b73c",x"3197",x"3b47",x"38b2",x"2ecb",x"3f9c",x"36eb",x"bbbf",x"b113",x"322d",x"3b4d",x"38ad",x"2eeb",x"3f9c",x"3713",x"bbc6",x"b1be",x"30de",x"3b4a",x"38a9"),
(x"303d",x"3f33",x"36eb",x"3b99",x"345f",x"30d6",x"3b27",x"3ba6",x"3051",x"3f24",x"36eb",x"3be6",x"2c79",x"308b",x"3b29",x"3b9e",x"3046",x"3f24",x"3711",x"3be4",x"2d1d",x"308b",x"3b24",x"3b9d"),
(x"2f3c",x"3f7a",x"3711",x"3934",x"ba0d",x"2c18",x"39f5",x"3ba5",x"2f42",x"3f79",x"36eb",x"374a",x"bb15",x"2de4",x"39fa",x"3ba4",x"2ede",x"3f73",x"36eb",x"3aaf",x"b860",x"2a70",x"39fa",x"3ba0"),
(x"3004",x"3f90",x"36eb",x"b8ae",x"3a73",x"2d47",x"3b5b",x"3864",x"3014",x"3f92",x"36eb",x"ae29",x"3be6",x"3005",x"3b5b",x"3863",x"3017",x"3f91",x"3711",x"b5dd",x"3b65",x"2eae",x"3b56",x"3864"),
(x"2eeb",x"3f9c",x"3713",x"bbc6",x"b1be",x"30de",x"3b4a",x"38a9",x"2ecb",x"3f9c",x"36eb",x"bbbf",x"b113",x"322d",x"3b4d",x"38ad",x"2ed7",x"3fa9",x"36eb",x"bbea",x"ae0a",x"2f12",x"3b52",x"38a8"),
(x"2f48",x"3f3a",x"36eb",x"bb01",x"3745",x"3141",x"3b2a",x"3b47",x"2f16",x"3f3e",x"3715",x"b9d1",x"b974",x"2cc6",x"3b26",x"3b44",x"2f49",x"3f3a",x"3718",x"baf6",x"b7e0",x"2460",x"3b25",x"3b46"),
(x"2f48",x"3f3a",x"36eb",x"bb01",x"3745",x"3141",x"3b2a",x"3b47",x"2ef5",x"3f3e",x"36eb",x"ba0e",x"b929",x"2e78",x"3b2b",x"3b44",x"2f16",x"3f3e",x"3715",x"b9d1",x"b974",x"2cc6",x"3b26",x"3b44"),
(x"3046",x"3f24",x"3711",x"3be4",x"2d1d",x"308b",x"3b24",x"3b9d",x"3051",x"3f24",x"36eb",x"3be6",x"2c79",x"308b",x"3b29",x"3b9e",x"304f",x"3f13",x"36eb",x"3be8",x"ad66",x"3010",x"3b2b",x"3b95"),
(x"2ed8",x"3f73",x"3717",x"3b6f",x"b5e5",x"261e",x"39f4",x"3ba0",x"2ede",x"3f73",x"36eb",x"3aaf",x"b860",x"2a70",x"39fa",x"3ba0",x"2ec6",x"3f6b",x"36eb",x"3bfa",x"ac62",x"2617",x"39fa",x"3b9c"),
(x"3014",x"3f92",x"36eb",x"ae29",x"3be6",x"3005",x"3b5b",x"3863",x"3043",x"3f92",x"36eb",x"3913",x"3a0d",x"310f",x"3b5a",x"3860",x"3038",x"3f91",x"3712",x"35a5",x"3b63",x"30cc",x"3b55",x"3861"),
(x"2ed7",x"3fa9",x"36eb",x"bbea",x"ae0a",x"2f12",x"3b52",x"38a8",x"2eaa",x"3fb4",x"36eb",x"bbe4",x"aadf",x"30ee",x"3b56",x"38a4",x"2ebe",x"3fb5",x"370f",x"bbdd",x"b0de",x"2e6c",x"3b53",x"38a0"),
(x"2ef5",x"3f3e",x"36eb",x"ba0e",x"b929",x"2e78",x"3b2b",x"3b44",x"2ec6",x"3f43",x"36eb",x"bbbf",x"b333",x"2ed2",x"3b2b",x"3b41",x"2ede",x"3f43",x"3718",x"bb13",x"b732",x"2fec",x"3b26",x"3b41"),
(x"304f",x"3f13",x"36eb",x"3be8",x"ad66",x"3010",x"3b2b",x"3b95",x"303e",x"3f0a",x"36eb",x"3ab2",x"b834",x"30cf",x"3b2c",x"3b91",x"3036",x"3f0b",x"3712",x"3b45",x"b640",x"30a6",x"3b27",x"3b90"),
(x"2fd1",x"3f20",x"3710",x"3b2f",x"36d9",x"2e52",x"3b8f",x"3666",x"2fe0",x"3f21",x"36eb",x"3b02",x"3776",x"2fc8",x"3b93",x"3666",x"2fec",x"3f1c",x"36eb",x"3bf4",x"9edc",x"2eb6",x"3b93",x"3662"),
(x"2ec2",x"3f6b",x"3715",x"3bfe",x"2412",x"286a",x"39f5",x"3b9b",x"2ec6",x"3f6b",x"36eb",x"3bfa",x"ac62",x"2617",x"39fa",x"3b9c",x"2ed7",x"3f61",x"36eb",x"3bcf",x"32aa",x"2bc8",x"39fa",x"3b96"),
(x"3043",x"3f92",x"36eb",x"3913",x"3a0d",x"310f",x"3b5a",x"3860",x"3057",x"3f8d",x"36eb",x"3be5",x"adbc",x"3036",x"3b59",x"385d",x"304c",x"3f8d",x"3711",x"3bb2",x"332f",x"30f4",x"3b55",x"385f"),
(x"2eaa",x"3fb4",x"36eb",x"bbe4",x"aadf",x"30ee",x"3b56",x"38a4",x"2eb7",x"3fba",x"36eb",x"baf6",x"3714",x"32f0",x"3b58",x"38a2",x"2ecd",x"3fb8",x"370d",x"bb0d",x"370c",x"3168",x"3b54",x"389f"),
(x"2ec6",x"3f43",x"36eb",x"bbbf",x"b333",x"2ed2",x"3b2b",x"3b41",x"2ecb",x"3f48",x"36eb",x"bbbf",x"3371",x"2dad",x"3b2b",x"3b3e",x"2ed4",x"3f47",x"3712",x"bbf0",x"2c20",x"2e95",x"3b27",x"3b3e"),
(x"303e",x"3f0a",x"36eb",x"3ab2",x"b834",x"30cf",x"3b2c",x"3b91",x"3007",x"3f02",x"36eb",x"37cb",x"bae6",x"3068",x"3b2c",x"3b8b",x"3003",x"3f04",x"3715",x"393c",x"b9e9",x"311d",x"3b27",x"3b8b"),
(x"2ece",x"3f60",x"3714",x"3b81",x"3558",x"2da6",x"39f5",x"3b96",x"2ed7",x"3f61",x"36eb",x"3bcf",x"32aa",x"2bc8",x"39fa",x"3b96",x"2f1f",x"3f59",x"36eb",x"3ac2",x"3833",x"2e85",x"39fa",x"3b91"),
(x"3057",x"3f8d",x"36eb",x"3be5",x"adbc",x"3036",x"3b59",x"385d",x"3044",x"3f85",x"36eb",x"3902",x"ba23",x"306a",x"3b57",x"3859",x"303e",x"3f87",x"3712",x"3ae4",x"b7c3",x"30c9",x"3b53",x"385c"),
(x"2ecd",x"3fb8",x"370d",x"bb0d",x"370c",x"3168",x"3b54",x"389f",x"2eb7",x"3fba",x"36eb",x"baf6",x"3714",x"32f0",x"3b58",x"38a2",x"2ee1",x"3fbb",x"36eb",x"b571",x"3b6d",x"30cc",x"3b59",x"38a0"),
(x"2ecb",x"3f48",x"36eb",x"bbbf",x"3371",x"2dad",x"3b2b",x"3b3e",x"2ed6",x"3f49",x"36eb",x"aeda",x"3bea",x"2e47",x"3b2b",x"3b3d",x"2ee4",x"3f49",x"3712",x"b297",x"3bcc",x"2d84",x"3b26",x"3b3d"),
(x"3007",x"3f02",x"36eb",x"37cb",x"bae6",x"3068",x"3b2c",x"3b8b",x"2f90",x"3f00",x"36eb",x"168d",x"bbf5",x"2e99",x"3b2d",x"3b87",x"2f91",x"3f01",x"3715",x"1ef6",x"bbee",x"302a",x"3b27",x"3b87"),
(x"2f11",x"3f58",x"3715",x"3a65",x"38c0",x"2d9c",x"39f5",x"3b91",x"2f1f",x"3f59",x"36eb",x"3ac2",x"3833",x"2e85",x"39fa",x"3b91",x"2f61",x"3f54",x"36eb",x"39cd",x"3979",x"2caa",x"39fa",x"3b8e"),
(x"3044",x"3f85",x"36eb",x"3902",x"ba23",x"306a",x"3b57",x"3859",x"3017",x"3f85",x"36eb",x"33f1",x"bbbc",x"2b5c",x"3b56",x"3857",x"301b",x"3f85",x"3713",x"3607",x"bb5e",x"2e4d",x"3b52",x"385a"),
(x"2ee7",x"3fba",x"3713",x"b451",x"3bac",x"2d81",x"3b54",x"389d",x"2ee1",x"3fbb",x"36eb",x"b571",x"3b6d",x"30cc",x"3b59",x"38a0",x"2f0d",x"3fbb",x"36eb",x"bbe3",x"2ce7",x"30c3",x"3b59",x"389f"),
(x"2ee4",x"3f49",x"3712",x"b297",x"3bcc",x"2d84",x"3b26",x"3b3d",x"2ed6",x"3f49",x"36eb",x"aeda",x"3bea",x"2e47",x"3b2b",x"3b3d",x"2f24",x"3f49",x"36eb",x"ac56",x"3bf7",x"2bc1",x"3b2b",x"3b3b"),
(x"2f91",x"3f01",x"3715",x"1ef6",x"bbee",x"302a",x"3b27",x"3b87",x"2f90",x"3f00",x"36eb",x"168d",x"bbf5",x"2e99",x"3b2d",x"3b87",x"2f13",x"3f02",x"36eb",x"b66a",x"bb44",x"2f81",x"3b2d",x"3b83"),
(x"2f5a",x"3f53",x"3717",x"3939",x"3a0b",x"29e0",x"39f5",x"3b8e",x"2f61",x"3f54",x"36eb",x"39cd",x"3979",x"2caa",x"39fa",x"3b8e",x"2f7e",x"3f52",x"36eb",x"b5a6",x"3b74",x"2d53",x"39fa",x"3b8d"),
(x"301b",x"3f85",x"3713",x"3607",x"bb5e",x"2e4d",x"3b52",x"385a",x"3017",x"3f85",x"36eb",x"33f1",x"bbbc",x"2b5c",x"3b56",x"3857",x"300f",x"3f84",x"36eb",x"394d",x"39f2",x"2dc5",x"3b55",x"3856"),
(x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1",x"2ffb",x"3fba",x"3715",x"99f0",x"a6cf",x"3bff",x"3b8e",x"3ba2",x"2f8b",x"3fa8",x"370e",x"3004",x"a71d",x"3bef",x"3b8a",x"3b93"),
(x"2f14",x"3fbc",x"3715",x"258e",x"307a",x"3beb",x"3b83",x"3ba2",x"2efa",x"3fc1",x"3712",x"a9f0",x"2b1d",x"3bfa",x"3b81",x"3ba6",x"2ffb",x"3fba",x"3715",x"99f0",x"a6cf",x"3bff",x"3b8e",x"3ba2"),
(x"2ffb",x"3fba",x"3715",x"99f0",x"a6cf",x"3bff",x"3b8e",x"3ba2",x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1",x"2f14",x"3fbc",x"3715",x"258e",x"307a",x"3beb",x"3b83",x"3ba2"),
(x"2f8b",x"3fa8",x"370e",x"3004",x"a71d",x"3bef",x"3b8a",x"3b93",x"2ee1",x"3faa",x"3717",x"2bf6",x"25ae",x"3bfb",x"3b82",x"3b93",x"2f10",x"3fba",x"3716",x"20ea",x"a780",x"3bfe",x"3b83",x"3ba1"),
(x"2f24",x"3f49",x"36eb",x"ac56",x"3bf7",x"2bc1",x"3b2b",x"3b3b",x"2f37",x"3f4a",x"36eb",x"bb71",x"b58a",x"2fc3",x"3b2b",x"3b3a",x"2f3a",x"3f49",x"3716",x"b8f4",x"3a42",x"2c09",x"3b26",x"3b3b"),
(x"2f0e",x"3f04",x"3713",x"b82e",x"baba",x"306c",x"3b28",x"3b82",x"2f13",x"3f02",x"36eb",x"b66a",x"bb44",x"2f81",x"3b2d",x"3b83",x"2e80",x"3f09",x"36eb",x"b9f2",x"b938",x"30b5",x"3b2c",x"3b7d"),
(x"2fd6",x"3f58",x"36eb",x"b976",x"39cc",x"2dcc",x"39fb",x"3b88",x"2fd3",x"3f57",x"3714",x"b97e",x"39c5",x"2dbf",x"39f5",x"3b88",x"2fa9",x"3f54",x"3714",x"b9a7",x"399f",x"2d1e",x"39f5",x"3b8a"),
(x"2fa9",x"3f54",x"3714",x"b9a7",x"399f",x"2d1e",x"39f5",x"3b8a",x"2f7e",x"3f52",x"36eb",x"b5a6",x"3b74",x"2d53",x"39fa",x"3b8d",x"2fd6",x"3f58",x"36eb",x"b976",x"39cc",x"2dcc",x"39fb",x"3b88"),
(x"300f",x"3f84",x"36eb",x"394d",x"39f2",x"2dc5",x"3b55",x"3856",x"303f",x"3f82",x"36eb",x"39ec",x"392b",x"31e4",x"3b54",x"3854",x"302f",x"3f81",x"3711",x"38c8",x"3a4e",x"30a8",x"3b50",x"3857"),
(x"2e95",x"3f0a",x"3715",x"bae0",x"b7cf",x"30d4",x"3b27",x"3b7d",x"2e80",x"3f09",x"36eb",x"b9f2",x"b938",x"30b5",x"3b2c",x"3b7d",x"2e4e",x"3f12",x"36eb",x"bbc4",x"b27a",x"3012",x"3b2c",x"3b77"),
(x"2fd6",x"3f58",x"36eb",x"b976",x"39cc",x"2dcc",x"39fb",x"3b88",x"3008",x"3f5b",x"36eb",x"b53f",x"3b87",x"2d28",x"39fb",x"3b86",x"300a",x"3f5a",x"3716",x"b7d5",x"3af0",x"2d8e",x"39f6",x"3b86"),
(x"303f",x"3f82",x"36eb",x"39ec",x"392b",x"31e4",x"3b54",x"3854",x"3065",x"3f79",x"36eb",x"3bbc",x"3212",x"3175",x"3b51",x"3850",x"3058",x"3f79",x"370f",x"3b4b",x"35cc",x"3223",x"3b4e",x"3853"),
(x"2edb",x"3fc1",x"36eb",x"bbdb",x"1c67",x"320a",x"3b5b",x"389c",x"2ef9",x"3fcd",x"36eb",x"bade",x"37ab",x"31d3",x"3b5e",x"3897",x"2f10",x"3fcc",x"370e",x"bb7b",x"34a9",x"3270",x"3b5a",x"3895"),
(x"2f48",x"3f4b",x"3715",x"bac2",x"b812",x"3146",x"3b26",x"3b3a",x"2ed7",x"3f52",x"36eb",x"badb",x"b7e7",x"30ac",x"3b2b",x"3b35",x"2f06",x"3f51",x"3718",x"bac6",x"b7dc",x"3286",x"3b26",x"3b36"),
(x"2e5f",x"3f13",x"3715",x"bbec",x"abe2",x"2fce",x"3b27",x"3b78",x"2e4e",x"3f12",x"36eb",x"bbc4",x"b27a",x"3012",x"3b2c",x"3b77",x"2e58",x"3f1c",x"36eb",x"bb6e",x"3575",x"309f",x"3b2b",x"3b73"),
(x"2ff3",x"3f30",x"3714",x"305e",x"21a1",x"3bec",x"3b92",x"3b30",x"3046",x"3f24",x"3711",x"2cd1",x"250b",x"3bf9",x"3b99",x"3b27",x"3024",x"3f23",x"3713",x"30f4",x"19bc",x"3be7",x"3b96",x"3b25"),
(x"2ff3",x"3f30",x"3714",x"305e",x"21a1",x"3bec",x"3b92",x"3b30",x"302e",x"3f34",x"3711",x"3115",x"27d5",x"3be4",x"3b97",x"3b33",x"3046",x"3f24",x"3711",x"2cd1",x"250b",x"3bf9",x"3b99",x"3b27"),
(x"3008",x"3f5b",x"36eb",x"b53f",x"3b87",x"2d28",x"39fb",x"3b86",x"302e",x"3f5c",x"36eb",x"33e5",x"3bb4",x"2ec2",x"39fb",x"3b84",x"302b",x"3f5b",x"3716",x"2345",x"3bf7",x"2dcc",x"39f6",x"3b83"),
(x"3065",x"3f79",x"36eb",x"3bbc",x"3212",x"3175",x"3b51",x"3850",x"3068",x"3f6f",x"36eb",x"3b61",x"b5a0",x"3119",x"3b4e",x"384c",x"305c",x"3f70",x"370f",x"3bd3",x"af46",x"3182",x"3b4b",x"384f"),
(x"2ed7",x"3f52",x"36eb",x"badb",x"b7e7",x"30ac",x"3b2b",x"3b35",x"2e89",x"3f5d",x"36eb",x"bbba",x"b376",x"2f14",x"3b2c",x"3b2e",x"2e9f",x"3f5d",x"3714",x"bb6b",x"b587",x"3096",x"3b26",x"3b2f"),
(x"2e58",x"3f1c",x"36eb",x"bb6e",x"3575",x"309f",x"3b2b",x"3b73",x"2ead",x"3f24",x"36eb",x"b884",x"3a69",x"324a",x"3b2a",x"3b6e",x"2ec0",x"3f22",x"3711",x"b8a4",x"3a69",x"309a",x"3b25",x"3b6f"),
(x"302e",x"3f5c",x"36eb",x"33e5",x"3bb4",x"2ec2",x"39fb",x"3b84",x"3050",x"3f5a",x"36eb",x"3acb",x"3812",x"3065",x"39fb",x"3b81",x"3045",x"3f59",x"3714",x"3976",x"39c0",x"3024",x"39f6",x"3b81"),
(x"3068",x"3f6f",x"36eb",x"3b61",x"b5a0",x"3119",x"3b4e",x"384c",x"3042",x"3f6a",x"36eb",x"386e",x"ba87",x"313e",x"3b4b",x"3849",x"3040",x"3f6b",x"370f",x"3891",x"ba72",x"30f5",x"3b48",x"384d"),
(x"2ef9",x"3fcd",x"36eb",x"bade",x"37ab",x"31d3",x"3b5e",x"3897",x"2f7f",x"3fd7",x"36eb",x"b8a6",x"3a54",x"3207",x"3b61",x"3891",x"2f7a",x"3fd4",x"3712",x"b8b5",x"3a3e",x"32bd",x"3b5c",x"388f"),
(x"2e89",x"3f5d",x"36eb",x"bbba",x"b376",x"2f14",x"3b2c",x"3b2e",x"2e6b",x"3f6a",x"36eb",x"bbef",x"2d0b",x"2e69",x"3b2c",x"3b27",x"2e7c",x"3f69",x"3712",x"bbf0",x"aa00",x"2f46",x"3b27",x"3b28"),
(x"2ec0",x"3f22",x"3711",x"b8a4",x"3a69",x"309a",x"3b25",x"3b6f",x"2ead",x"3f24",x"36eb",x"b884",x"3a69",x"324a",x"3b2a",x"3b6e",x"2f34",x"3f26",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3b28",x"3b6a"),
(x"3050",x"3f5a",x"36eb",x"3acb",x"3812",x"3065",x"39fb",x"3b81",x"305c",x"3f54",x"36eb",x"3bcf",x"b173",x"3043",x"39fb",x"3b7e",x"3050",x"3f55",x"3712",x"3be0",x"2e5e",x"30a3",x"39f6",x"3b7f"),
(x"3040",x"3f6b",x"370f",x"3891",x"ba72",x"30f5",x"3b48",x"384d",x"3042",x"3f6a",x"36eb",x"386e",x"ba87",x"313e",x"3b4b",x"3849",x"3013",x"3f68",x"36eb",x"b5e4",x"bb4d",x"31a2",x"3b48",x"3847"),
(x"2f7a",x"3fd4",x"3712",x"b8b5",x"3a3e",x"32bd",x"3b5c",x"388f",x"2f7f",x"3fd7",x"36eb",x"b8a6",x"3a54",x"3207",x"3b61",x"3891",x"2fd0",x"3fd7",x"36eb",x"3996",x"395e",x"33ec",x"3b61",x"388e"),
(x"2e6b",x"3f6a",x"36eb",x"bbef",x"2d0b",x"2e69",x"3b2c",x"3b27",x"2e95",x"3f76",x"36eb",x"bb75",x"35a2",x"2d46",x"3b2b",x"3b21",x"2ea0",x"3f75",x"3710",x"bb6a",x"35bb",x"2efe",x"3b27",x"3b21"),
(x"2f3e",x"3f25",x"3718",x"b8ae",x"3a78",x"2b7c",x"3b23",x"3b6c",x"2f34",x"3f26",x"36eb",x"b60d",x"3b5a",x"2ef3",x"3b28",x"3b6a",x"2f4a",x"3f28",x"36eb",x"bbe6",x"308f",x"2c41",x"3b28",x"3b68"),
(x"305c",x"3f54",x"36eb",x"3bcf",x"b173",x"3043",x"39fb",x"3b7e",x"3048",x"3f4f",x"36eb",x"36fe",x"bb25",x"2ea4",x"39fa",x"3b7b",x"3044",x"3f51",x"3714",x"3972",x"b9bb",x"30de",x"39f5",x"3b7d"),
(x"302f",x"3f1a",x"3710",x"a828",x"260a",x"3bfe",x"3b97",x"3b1e",x"3024",x"3f23",x"3713",x"30f4",x"19bc",x"3be7",x"3b96",x"3b25",x"3046",x"3f24",x"3711",x"2cd1",x"250b",x"3bf9",x"3b99",x"3b27"),
(x"3046",x"3f13",x"3714",x"aeb0",x"28fa",x"3bf3",x"3b9a",x"3b19",x"302b",x"3f12",x"3714",x"a949",x"1ffc",x"3bfe",x"3b97",x"3b18",x"302f",x"3f1a",x"3710",x"a828",x"260a",x"3bfe",x"3b97",x"3b1e"),
(x"3036",x"3f0b",x"3712",x"2587",x"208e",x"3bff",x"3b98",x"3b12",x"302b",x"3f12",x"3714",x"a949",x"1ffc",x"3bfe",x"3b97",x"3b18",x"3046",x"3f13",x"3714",x"aeb0",x"28fa",x"3bf3",x"3b9a",x"3b19"),
(x"3036",x"3f0b",x"3712",x"2587",x"208e",x"3bff",x"3b98",x"3b12",x"3021",x"3f0e",x"3712",x"a953",x"27ae",x"3bfd",x"3b96",x"3b14",x"302b",x"3f12",x"3714",x"a949",x"1ffc",x"3bfe",x"3b97",x"3b18"),
(x"3003",x"3f04",x"3715",x"20ea",x"2afd",x"3bfc",x"3b94",x"3b0c",x"2fe4",x"3f08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3b92",x"3b0f",x"300e",x"3f0b",x"3714",x"28bf",x"2c20",x"3bfa",x"3b95",x"3b11"),
(x"2f91",x"3f01",x"3715",x"a7e2",x"29b2",x"3bfc",x"3b8e",x"3b09",x"2f7e",x"3f06",x"3715",x"a70a",x"a779",x"3bfe",x"3b8d",x"3b0d",x"2fe4",x"3f08",x"3714",x"a31d",x"2b5f",x"3bfc",x"3b92",x"3b0f"),
(x"2f0e",x"3f04",x"3713",x"ab1d",x"aee4",x"3bf0",x"3b88",x"3b0b",x"2f19",x"3f08",x"3716",x"a4bc",x"aceb",x"3bf9",x"3b89",x"3b0e",x"2f7e",x"3f06",x"3715",x"a70a",x"a779",x"3bfe",x"3b8d",x"3b0d"),
(x"2e95",x"3f0a",x"3715",x"2266",x"9d87",x"3bff",x"3b82",x"3b10",x"2ec8",x"3f0e",x"3714",x"28e0",x"299e",x"3bfc",x"3b85",x"3b13",x"2f19",x"3f08",x"3716",x"a4bc",x"aceb",x"3bf9",x"3b89",x"3b0e"),
(x"2e5f",x"3f13",x"3715",x"2891",x"a7ce",x"3bfd",x"3b7f",x"3b17",x"2eb5",x"3f13",x"3714",x"2538",x"a9ab",x"3bfd",x"3b83",x"3b18",x"2ec8",x"3f0e",x"3714",x"28e0",x"299e",x"3bfc",x"3b85",x"3b13"),
(x"2e5f",x"3f13",x"3715",x"2891",x"a7ce",x"3bfd",x"3b7f",x"3b17",x"2e70",x"3f1b",x"3717",x"2d06",x"2793",x"3bf8",x"3b80",x"3b1e",x"2ed5",x"3f18",x"3715",x"2c67",x"28a5",x"3bf9",x"3b85",x"3b1b"),
(x"2ec0",x"3f22",x"3711",x"28d9",x"a52b",x"3bfe",x"3b83",x"3b24",x"2f14",x"3f18",x"3714",x"2a45",x"2b10",x"3bfa",x"3b88",x"3b1c",x"2ed5",x"3f18",x"3715",x"2c67",x"28a5",x"3bf9",x"3b85",x"3b1b"),
(x"2fc4",x"3f19",x"3711",x"2bef",x"a8a8",x"3bfa",x"3b90",x"3b1d",x"2f9c",x"3f16",x"3710",x"2352",x"ae7e",x"3bf5",x"3b8e",x"3b1a",x"2f4a",x"3f16",x"3711",x"2a66",x"b31a",x"3bca",x"3b8a",x"3b1a"),
(x"2f99",x"3f25",x"3713",x"341f",x"ac3c",x"3bb6",x"3b8d",x"3b26",x"2faf",x"3f23",x"3711",x"340b",x"26c2",x"3bbc",x"3b8f",x"3b25",x"2f3e",x"3f25",x"3718",x"2b65",x"b528",x"3b8f",x"3b89",x"3b27"),
(x"2f94",x"3f29",x"3714",x"2de0",x"a4c2",x"3bf6",x"3b8d",x"3b2a",x"2f55",x"3f28",x"3718",x"3420",x"1418",x"3bba",x"3b8a",x"3b29",x"2f5a",x"3f31",x"3715",x"27ae",x"a4ea",x"3bfe",x"3b8a",x"3b31"),
(x"2f94",x"3f29",x"3714",x"2de0",x"a4c2",x"3bf6",x"3b8d",x"3b2a",x"2f99",x"3f25",x"3713",x"341f",x"ac3c",x"3bb6",x"3b8d",x"3b26",x"2f55",x"3f28",x"3718",x"3420",x"1418",x"3bba",x"3b8a",x"3b29"),
(x"2fc4",x"3f19",x"3711",x"2bef",x"a8a8",x"3bfa",x"3b90",x"3b1d",x"2fd1",x"3f20",x"3710",x"2856",x"a9ab",x"3bfc",x"3b90",x"3b23",x"2fdc",x"3f1c",x"3710",x"2a8d",x"2973",x"3bfb",x"3b91",x"3b1f"),
(x"2f14",x"3f18",x"3714",x"2a45",x"2b10",x"3bfa",x"3b88",x"3b1c",x"2ec0",x"3f22",x"3711",x"28d9",x"a52b",x"3bfe",x"3b83",x"3b24",x"2fd1",x"3f20",x"3710",x"2856",x"a9ab",x"3bfc",x"3b90",x"3b23"),
(x"301e",x"3ec3",x"3718",x"224c",x"a36c",x"3bff",x"3990",x"326f",x"2fd9",x"3edf",x"3716",x"282f",x"2808",x"3bfd",x"398c",x"32b2",x"3033",x"3ee0",x"3715",x"21a1",x"23fc",x"3bff",x"3991",x"32b4"),
(x"2f9f",x"3f25",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b93",x"366c",x"2f99",x"3f25",x"3713",x"3bc2",x"33a4",x"298a",x"3b8e",x"366b",x"2f94",x"3f29",x"3714",x"3bf3",x"ae23",x"2b27",x"3b8e",x"3670"),
(x"2f94",x"3f29",x"3714",x"3bf3",x"ae23",x"2b27",x"3b8e",x"3670",x"2fb5",x"3f36",x"36eb",x"346a",x"bb91",x"316a",x"3b92",x"367e",x"2f9f",x"3f25",x"36eb",x"3bf6",x"2a70",x"2d61",x"3b93",x"366c"),
(x"3008",x"3de5",x"370e",x"2fd2",x"a717",x"3bef",x"386c",x"38b1",x"2fa8",x"3ddc",x"3712",x"342b",x"ae69",x"3bae",x"3866",x"38a6",x"2f67",x"3ddc",x"3716",x"30f9",x"28af",x"3be5",x"3862",x"38a6"),
(x"2f67",x"3ddc",x"3716",x"badd",x"b75a",x"334d",x"3b13",x"3a46",x"2f52",x"3dd9",x"36eb",x"b996",x"b95e",x"33ec",x"3b19",x"3a47",x"2eeb",x"3de9",x"36eb",x"bb99",x"b315",x"330d",x"3b18",x"3a3e"),
(x"2f72",x"3e29",x"3714",x"ac39",x"a9a5",x"3bf9",x"385b",x"38fe",x"2f3e",x"3e22",x"3713",x"ada3",x"af14",x"3beb",x"3858",x"38f5",x"2f20",x"3e21",x"3712",x"aa69",x"a87e",x"3bfc",x"3856",x"38f5"),
(x"2ef3",x"3e1f",x"3711",x"a994",x"a977",x"3bfc",x"3853",x"38f2",x"2eb1",x"3e20",x"3712",x"2a38",x"2d35",x"3bf6",x"384f",x"38f3",x"2e89",x"3e24",x"3711",x"a481",x"a546",x"3bff",x"384c",x"38f7"),
(x"2ea4",x"3e29",x"3712",x"aa73",x"aa97",x"3bfa",x"384e",x"38fd",x"2eea",x"3e2b",x"3713",x"a91b",x"ab55",x"3bfb",x"3852",x"38ff",x"2f20",x"3e21",x"3712",x"aa69",x"a87e",x"3bfc",x"3856",x"38f5"),
(x"2f2f",x"3e2e",x"3718",x"ae36",x"2160",x"3bf6",x"3857",x"3903",x"2f0a",x"3e2d",x"3716",x"af14",x"b29c",x"3bc6",x"3854",x"3902",x"2ec3",x"3e2f",x"3711",x"afec",x"2c2c",x"3beb",x"384f",x"3904"),
(x"2eec",x"3e47",x"3713",x"ae9a",x"b366",x"3bbd",x"3850",x"391f",x"2f31",x"3e42",x"370f",x"2b8a",x"b0af",x"3be6",x"3855",x"391a",x"2f2d",x"3e3f",x"370e",x"26d5",x"a5c2",x"3bfe",x"3855",x"3917"),
(x"2efb",x"3e3b",x"3713",x"a538",x"2c79",x"3bfa",x"3852",x"3912",x"2e69",x"3e40",x"370f",x"acd8",x"271d",x"3bf9",x"3848",x"3917",x"2ea1",x"3e45",x"370f",x"9df0",x"2631",x"3bff",x"384b",x"391d"),
(x"2efb",x"3e3b",x"3713",x"a538",x"2c79",x"3bfa",x"3852",x"3912",x"2efa",x"3e39",x"3713",x"a7e9",x"a849",x"3bfd",x"3852",x"390f",x"2e71",x"3e37",x"370f",x"aec5",x"9a24",x"3bf4",x"3849",x"390d"),
(x"2ec3",x"3e2f",x"3711",x"afec",x"2c2c",x"3beb",x"384f",x"3904",x"2e71",x"3e37",x"370f",x"aec5",x"9a24",x"3bf4",x"3849",x"390d",x"2efa",x"3e39",x"3713",x"a7e9",x"a849",x"3bfd",x"3852",x"390f"),
(x"2f21",x"3e36",x"3710",x"ac5b",x"30a5",x"3be5",x"3855",x"390d",x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908",x"2ec3",x"3e2f",x"3711",x"afec",x"2c2c",x"3beb",x"384f",x"3904"),
(x"2f21",x"3e36",x"3710",x"ac5b",x"30a5",x"3be5",x"3855",x"390d",x"2f61",x"3e35",x"3713",x"25b5",x"37de",x"3af6",x"385a",x"390b",x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908"),
(x"2fda",x"3e66",x"3715",x"a6c2",x"2c63",x"3bfa",x"3861",x"3943",x"2fc7",x"3e5d",x"3717",x"97c8",x"1f79",x"3c00",x"3860",x"3939",x"2fa2",x"3e5e",x"3717",x"aff2",x"2a7d",x"3bed",x"385e",x"393b"),
(x"2ecb",x"3e55",x"3716",x"acd8",x"27e2",x"3bf9",x"3850",x"3930",x"2e97",x"3e57",x"3714",x"a860",x"2f8b",x"3bf0",x"384d",x"3932",x"2e81",x"3e5b",x"3712",x"b162",x"2345",x"3be2",x"384b",x"3937"),
(x"2e99",x"3e5f",x"3714",x"1553",x"2b62",x"3bfc",x"384d",x"393c",x"2f21",x"3e62",x"3711",x"240b",x"2d5c",x"3bf8",x"3855",x"393f",x"2f0c",x"3e56",x"3716",x"2818",x"2d04",x"3bf8",x"3854",x"3931"),
(x"2f79",x"3e5c",x"3714",x"b036",x"273e",x"3bed",x"385b",x"3939",x"2f4f",x"3e59",x"3714",x"a4fd",x"2dab",x"3bf7",x"3858",x"3935",x"2f21",x"3e62",x"3711",x"240b",x"2d5c",x"3bf8",x"3855",x"393f"),
(x"2f3f",x"3e64",x"3711",x"b27d",x"975f",x"3bd5",x"3857",x"3941",x"2fa2",x"3e5e",x"3717",x"aff2",x"2a7d",x"3bed",x"385e",x"393b",x"2f79",x"3e5c",x"3714",x"b036",x"273e",x"3bed",x"385b",x"3939"),
(x"2f3f",x"3e64",x"3711",x"b27d",x"975f",x"3bd5",x"3857",x"3941",x"2f4a",x"3e66",x"3712",x"af67",x"2981",x"3bf0",x"3858",x"3943",x"2fa2",x"3e5e",x"3717",x"aff2",x"2a7d",x"3bed",x"385e",x"393b"),
(x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b",x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"2f3b",x"3e6b",x"3712",x"b146",x"ac91",x"3bde",x"3857",x"3949"),
(x"2fe4",x"3e77",x"3718",x"2138",x"2e95",x"3bf4",x"3862",x"3957",x"2fd6",x"3e7d",x"3715",x"28bf",x"2fdb",x"3bef",x"3861",x"395d",x"3017",x"3e78",x"3719",x"a90e",x"2f00",x"3bf2",x"3867",x"3958"),
(x"2fd8",x"3e76",x"3718",x"2b4f",x"a525",x"3bfc",x"3861",x"3956",x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"2f6c",x"3e7b",x"3718",x"ae3b",x"9fae",x"3bf6",x"385a",x"395b"),
(x"2fd8",x"3e76",x"3718",x"2b4f",x"a525",x"3bfc",x"3861",x"3956",x"3006",x"3e73",x"3715",x"2d65",x"2c5a",x"3bf3",x"3865",x"3952",x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d"),
(x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"3006",x"3e73",x"3715",x"2d65",x"2c5a",x"3bf3",x"3865",x"3952",x"3022",x"3e6e",x"3718",x"2cf2",x"98ea",x"3bf9",x"3868",x"394c"),
(x"3027",x"3e69",x"3712",x"359c",x"b36a",x"3b42",x"3869",x"3947",x"301e",x"3e68",x"3712",x"3542",x"b0ba",x"3b76",x"3868",x"3945",x"3002",x"3e68",x"3717",x"2d2d",x"aecd",x"3bed",x"3864",x"3946"),
(x"2faf",x"3e6e",x"3718",x"abb4",x"a8d3",x"3bfa",x"385f",x"394d",x"3002",x"3e68",x"3717",x"2d2d",x"aecd",x"3bed",x"3864",x"3946",x"2fe7",x"3e67",x"3716",x"b009",x"ada8",x"3be7",x"3862",x"3945"),
(x"2f4a",x"3e66",x"3712",x"af67",x"2981",x"3bf0",x"3858",x"3943",x"2f3b",x"3e6b",x"3712",x"b146",x"ac91",x"3bde",x"3857",x"3949",x"2fe7",x"3e67",x"3716",x"b009",x"ada8",x"3be7",x"3862",x"3945"),
(x"2fc7",x"3e5d",x"3717",x"97c8",x"1f79",x"3c00",x"3860",x"3939",x"300d",x"3e5f",x"3718",x"ac00",x"a90e",x"3bfa",x"3866",x"393c",x"3008",x"3e58",x"3715",x"a518",x"ad04",x"3bf9",x"3865",x"3934"),
(x"2fc7",x"3e5d",x"3717",x"97c8",x"1f79",x"3c00",x"3860",x"3939",x"2fe5",x"3e63",x"3714",x"a581",x"2e8a",x"3bf4",x"3862",x"3940",x"300d",x"3e5f",x"3718",x"ac00",x"a90e",x"3bfa",x"3866",x"393c"),
(x"3008",x"3e58",x"3715",x"a518",x"ad04",x"3bf9",x"3865",x"3934",x"300d",x"3e5f",x"3718",x"ac00",x"a90e",x"3bfa",x"3866",x"393c",x"3041",x"3e53",x"3714",x"175f",x"ac2c",x"3bfb",x"386d",x"392f"),
(x"302a",x"3e50",x"3714",x"2dba",x"a266",x"3bf7",x"386a",x"392b",x"3041",x"3e53",x"3714",x"175f",x"ac2c",x"3bfb",x"386d",x"392f",x"3052",x"3e47",x"3712",x"3106",x"a73e",x"3be5",x"386f",x"3920"),
(x"302f",x"3e45",x"3715",x"3468",x"a47a",x"3bb0",x"386a",x"391f",x"3052",x"3e47",x"3712",x"3106",x"a73e",x"3be5",x"386f",x"3920",x"3041",x"3e3b",x"3710",x"3550",x"ae33",x"3b81",x"386c",x"3913"),
(x"3025",x"3e3d",x"3717",x"3273",x"af43",x"3bc8",x"3868",x"3915",x"3041",x"3e3b",x"3710",x"3550",x"ae33",x"3b81",x"386c",x"3913",x"3015",x"3e33",x"3712",x"2b5f",x"a345",x"3bfc",x"3867",x"390a"),
(x"2fa3",x"3e35",x"3712",x"2dd2",x"304b",x"3be4",x"385e",x"390c",x"2f75",x"3e2e",x"3716",x"2f4d",x"2a5f",x"3bf0",x"385b",x"3903",x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908"),
(x"2fa3",x"3e35",x"3712",x"2dd2",x"304b",x"3be4",x"385e",x"390c",x"3015",x"3e33",x"3712",x"2b5f",x"a345",x"3bfc",x"3867",x"390a",x"2f75",x"3e2e",x"3716",x"2f4d",x"2a5f",x"3bf0",x"385b",x"3903"),
(x"2fa3",x"3e35",x"3712",x"2dd2",x"304b",x"3be4",x"385e",x"390c",x"2fe6",x"3e36",x"3711",x"ae24",x"aa2b",x"3bf4",x"3862",x"390d",x"3015",x"3e33",x"3712",x"2b5f",x"a345",x"3bfc",x"3867",x"390a"),
(x"2f2f",x"3e2e",x"3718",x"ae36",x"2160",x"3bf6",x"3857",x"3903",x"2f67",x"3e32",x"3718",x"ac13",x"31c5",x"3bda",x"385a",x"3908",x"2f75",x"3e2e",x"3716",x"2f4d",x"2a5f",x"3bf0",x"385b",x"3903"),
(x"2f0a",x"3e2d",x"3716",x"af14",x"b29c",x"3bc6",x"3854",x"3902",x"2f72",x"3e29",x"3714",x"ac39",x"a9a5",x"3bf9",x"385b",x"38fe",x"2eea",x"3e2b",x"3713",x"a91b",x"ab55",x"3bfb",x"3852",x"38ff"),
(x"2f0a",x"3e2d",x"3716",x"af14",x"b29c",x"3bc6",x"3854",x"3902",x"2f5c",x"3e2c",x"3716",x"a553",x"b2c7",x"3bd1",x"385a",x"3901",x"2f72",x"3e29",x"3714",x"ac39",x"a9a5",x"3bf9",x"385b",x"38fe"),
(x"2f3e",x"3e22",x"3713",x"ada3",x"af14",x"3beb",x"3858",x"38f5",x"2f72",x"3e29",x"3714",x"ac39",x"a9a5",x"3bf9",x"385b",x"38fe",x"2fe6",x"3e22",x"3717",x"b0e7",x"b057",x"3bd4",x"3863",x"38f6"),
(x"2f93",x"3e1d",x"370f",x"aedc",x"acd0",x"3bee",x"385e",x"38f0",x"2fe6",x"3e22",x"3717",x"b0e7",x"b057",x"3bd4",x"3863",x"38f6",x"301b",x"3e14",x"3713",x"a9b8",x"26e9",x"3bfd",x"3869",x"38e7"),
(x"302a",x"3df8",x"370d",x"3809",x"ae09",x"3add",x"386f",x"38c7",x"301d",x"3df6",x"3713",x"2f9f",x"3907",x"3a25",x"386d",x"38c5",x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4"),
(x"2f13",x"3dea",x"3715",x"2d56",x"a0d0",x"3bf8",x"385b",x"38b5",x"2f27",x"3df7",x"3715",x"19bc",x"26cf",x"3bff",x"385b",x"38c3",x"3013",x"3def",x"3712",x"29f0",x"ab1d",x"3bfa",x"386c",x"38bd"),
(x"2f02",x"3df7",x"36eb",x"bb89",x"3473",x"31fc",x"3b17",x"3a37",x"2f8f",x"3e09",x"36eb",x"bb4a",x"3677",x"2cfa",x"3b15",x"3a2d",x"2f97",x"3e08",x"370e",x"bb5f",x"35f1",x"2f4d",x"3b10",x"3a2e"),
(x"2ece",x"3e8d",x"36eb",x"3ba1",x"34cc",x"1f45",x"3a16",x"3a29",x"2ed8",x"3e8e",x"3713",x"3ba5",x"3497",x"ac28",x"3a11",x"3a29",x"2ec4",x"3e97",x"3710",x"3bfd",x"2997",x"a09b",x"3a11",x"3a2e"),
(x"2ec4",x"3e97",x"3710",x"3bfd",x"2997",x"a09b",x"3a11",x"3a2e",x"2ec5",x"3e9c",x"36eb",x"3bf5",x"ae59",x"2467",x"3a16",x"3a31",x"2ece",x"3e8d",x"36eb",x"3ba1",x"34cc",x"1f45",x"3a16",x"3a29"),
(x"2f6c",x"3e7b",x"36eb",x"b46a",x"3b91",x"316a",x"3a15",x"3a1e",x"2f6c",x"3e7b",x"3718",x"b9e5",x"3968",x"0000",x"3a10",x"3a1e",x"2f2f",x"3e80",x"3714",x"3b1c",x"3754",x"223f",x"3a10",x"3a22"),
(x"2f2f",x"3e80",x"3714",x"3b1c",x"3754",x"223f",x"3a10",x"3a22",x"2ece",x"3e8d",x"36eb",x"3ba1",x"34cc",x"1f45",x"3a16",x"3a29",x"2f6c",x"3e7b",x"36eb",x"b46a",x"3b91",x"316a",x"3a15",x"3a1e"),
(x"2ec5",x"3e9c",x"36eb",x"3bf5",x"ae59",x"2467",x"3a16",x"3a31",x"2eca",x"3e9e",x"3714",x"3beb",x"b08b",x"98ea",x"3a11",x"3a32",x"2edf",x"3ea3",x"3712",x"3b76",x"b5c5",x"204d",x"3a11",x"3a34"),
(x"2edf",x"3ea3",x"3712",x"3b76",x"b5c5",x"204d",x"3a11",x"3a34",x"2ee8",x"3ea4",x"36eb",x"3ab1",x"b862",x"21f0",x"3a16",x"3a35",x"2ec5",x"3e9c",x"36eb",x"3bf5",x"ae59",x"2467",x"3a16",x"3a31"),
(x"2f38",x"3ea8",x"36eb",x"37e1",x"baf5",x"269a",x"3a16",x"3a38",x"2ee8",x"3ea4",x"36eb",x"3ab1",x"b862",x"21f0",x"3a16",x"3a35",x"2f06",x"3ea6",x"3714",x"395a",x"b9f1",x"2032",x"3a11",x"3a36"),
(x"2f9e",x"3eaa",x"36eb",x"303c",x"bbeb",x"299b",x"3a16",x"3a3c",x"2f38",x"3ea8",x"36eb",x"37e1",x"baf5",x"269a",x"3a16",x"3a38",x"2f3d",x"3ea8",x"3714",x"35bf",x"bb76",x"27db",x"3a11",x"3a39"),
(x"3003",x"3ea9",x"36eb",x"b868",x"baab",x"296a",x"3a16",x"3a3f",x"2f9e",x"3eaa",x"36eb",x"303c",x"bbeb",x"299b",x"3a16",x"3a3c",x"2fa3",x"3eaa",x"3715",x"a836",x"bbfd",x"294c",x"3a11",x"3a3c"),
(x"302c",x"3ea3",x"3714",x"bb01",x"b7b5",x"2839",x"3a12",x"3a44",x"3029",x"3ea2",x"36eb",x"baf3",x"b7df",x"2b38",x"3a17",x"3a43",x"3003",x"3ea9",x"36eb",x"b868",x"baab",x"296a",x"3a16",x"3a3f"),
(x"3036",x"3e9d",x"36eb",x"bbf9",x"ad11",x"2511",x"3a17",x"3a46",x"3029",x"3ea2",x"36eb",x"baf3",x"b7df",x"2b38",x"3a17",x"3a43",x"302c",x"3ea3",x"3714",x"bb01",x"b7b5",x"2839",x"3a12",x"3a44"),
(x"3029",x"3e99",x"36eb",x"b90c",x"3a34",x"2532",x"3a17",x"3a49",x"3036",x"3e9d",x"36eb",x"bbf9",x"ad11",x"2511",x"3a17",x"3a46",x"3036",x"3e9d",x"3714",x"bbe6",x"310f",x"9bfc",x"3a12",x"3a47"),
(x"3006",x"3e98",x"3714",x"2fe2",x"3bee",x"28fd",x"3a12",x"3a4b",x"3004",x"3e98",x"36eb",x"35dd",x"3b6d",x"2be9",x"3a17",x"3a4b",x"3029",x"3e99",x"36eb",x"b90c",x"3a34",x"2532",x"3a17",x"3a49"),
(x"2fd7",x"3e9a",x"3711",x"364f",x"3b52",x"2d1b",x"3a13",x"3a4d",x"2fdd",x"3e9b",x"36eb",x"32b1",x"3bc8",x"2e54",x"3a18",x"3a4d",x"3004",x"3e98",x"36eb",x"35dd",x"3b6d",x"2be9",x"3a17",x"3a4b"),
(x"2f82",x"3e8c",x"36eb",x"bbf6",x"aa70",x"2d60",x"3a17",x"3a5a",x"2f71",x"3e8d",x"36eb",x"b9db",x"b96c",x"2c1a",x"3a17",x"3a59",x"2f73",x"3e8e",x"3711",x"ba7a",x"b8af",x"2839",x"3a12",x"3a58"),
(x"2f85",x"3e9a",x"3710",x"b416",x"3bad",x"2f8d",x"3a13",x"3a50",x"2f79",x"3e9b",x"36eb",x"b37e",x"3bba",x"2ef6",x"3a18",x"3a50",x"2fdd",x"3e9b",x"36eb",x"32b1",x"3bc8",x"2e54",x"3a18",x"3a4d"),
(x"2efa",x"3e48",x"36eb",x"35e4",x"3b4d",x"31a2",x"3b21",x"3b72",x"2f46",x"3e42",x"36eb",x"3b7d",x"3521",x"3096",x"3b1f",x"3b6f",x"2f31",x"3e42",x"370f",x"3a9c",x"3854",x"30fa",x"3b1b",x"3b71"),
(x"2f13",x"3dea",x"3715",x"bbc5",x"ab9a",x"3358",x"3b13",x"3a3f",x"2eeb",x"3de9",x"36eb",x"bb99",x"b315",x"330d",x"3b18",x"3a3e",x"2f02",x"3df7",x"36eb",x"bb89",x"3473",x"31fc",x"3b17",x"3a37"),
(x"2f51",x"3e90",x"3710",x"a856",x"29ab",x"3bfc",x"3858",x"3973",x"3030",x"3e8e",x"3711",x"a8d9",x"252b",x"3bfe",x"386a",x"3972",x"2fe3",x"3e8b",x"3718",x"ab65",x"3528",x"3b8f",x"3862",x"396d"),
(x"300a",x"3df5",x"36eb",x"3be3",x"ace8",x"30c3",x"3b11",x"3a58",x"3013",x"3def",x"3712",x"3bcf",x"3082",x"3141",x"3b0f",x"3a53",x"3006",x"3df4",x"3715",x"3bd7",x"31f9",x"2c2a",x"3b0d",x"3a55"),
(x"300a",x"3df5",x"36eb",x"3be3",x"ace8",x"30c3",x"3b11",x"3a58",x"3023",x"3def",x"36eb",x"3bdb",x"9c67",x"320a",x"3b13",x"3a55",x"3013",x"3def",x"3712",x"3bcf",x"3082",x"3141",x"3b0f",x"3a53"),
(x"3041",x"3e3b",x"3710",x"3b6a",x"b5bb",x"2efe",x"3a23",x"3a52",x"3046",x"3e3a",x"36eb",x"3b75",x"b5a2",x"2d46",x"3a27",x"3a52",x"301f",x"3e33",x"36eb",x"3958",x"b9de",x"2fe4",x"3a27",x"3a4d"),
(x"2f4e",x"3e99",x"36eb",x"baa4",x"3859",x"2fe4",x"3a18",x"3a52",x"2f79",x"3e9b",x"36eb",x"b37e",x"3bba",x"2ef6",x"3a18",x"3a50",x"2f85",x"3e9a",x"3710",x"b416",x"3bad",x"2f8d",x"3a13",x"3a50"),
(x"2fd8",x"3e89",x"36eb",x"3be6",x"b08e",x"2c41",x"3b49",x"38d4",x"2fd4",x"3e7f",x"36eb",x"3bfa",x"20b5",x"2cbc",x"3b47",x"38d2",x"2fc7",x"3e7f",x"3715",x"3bfa",x"2710",x"2c48",x"3b44",x"38d3"),
(x"2f45",x"3e94",x"3710",x"bbcc",x"3227",x"2f2e",x"3a13",x"3a54",x"2f36",x"3e94",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3a18",x"3a55",x"2f4e",x"3e99",x"36eb",x"baa4",x"3859",x"2fe4",x"3a18",x"3a52"),
(x"2f46",x"3e42",x"36eb",x"3b7d",x"3521",x"3096",x"3b1f",x"3b6f",x"2f3c",x"3e3f",x"36eb",x"3b19",x"b744",x"2cf7",x"3b1e",x"3b6d",x"2f2d",x"3e3f",x"370e",x"3b25",x"b70d",x"2d6a",x"3b1a",x"3b70"),
(x"2e90",x"3e61",x"36eb",x"b6fe",x"3b25",x"2ea4",x"3b4e",x"38fe",x"2f2b",x"3e63",x"36eb",x"b7d8",x"3af6",x"2a35",x"3b4f",x"38fc",x"2f21",x"3e62",x"3711",x"b4dc",x"3b97",x"2d61",x"3b4b",x"38fc"),
(x"2f71",x"3e8d",x"36eb",x"b9db",x"b96c",x"2c1a",x"3a17",x"3a59",x"2f41",x"3e90",x"36eb",x"bb02",x"b776",x"2fc8",x"3a17",x"3a57",x"2f51",x"3e90",x"3710",x"bb2f",x"b6d9",x"2e52",x"3a13",x"3a56"),
(x"3015",x"3e33",x"3712",x"384e",x"bab0",x"2ec8",x"3a23",x"3a4d",x"301f",x"3e33",x"36eb",x"3958",x"b9de",x"2fe4",x"3a27",x"3a4d",x"2f6d",x"3e2d",x"36eb",x"3776",x"bb0b",x"2d41",x"3a27",x"3a45"),
(x"2fc7",x"3e7f",x"3715",x"3bfa",x"2710",x"2c48",x"3b44",x"38d3",x"2fd4",x"3e7f",x"36eb",x"3bfa",x"20b5",x"2cbc",x"3b47",x"38d2",x"2fd9",x"3e7e",x"36eb",x"39df",x"3964",x"2d28",x"3b47",x"38d2"),
(x"2f2d",x"3e3f",x"370e",x"3b25",x"b70d",x"2d6a",x"3b1a",x"3b70",x"2f3c",x"3e3f",x"36eb",x"3b19",x"b744",x"2cf7",x"3b1e",x"3b6d",x"2f02",x"3e3a",x"36eb",x"3ad3",x"b822",x"2c4d",x"3b1c",x"3b6b"),
(x"2f97",x"3e08",x"370e",x"bb5f",x"35f1",x"2f4d",x"3b10",x"3a2e",x"2f8f",x"3e09",x"36eb",x"bb4a",x"3677",x"2cfa",x"3b15",x"3a2d",x"2fc6",x"3e13",x"36eb",x"bbfe",x"9ea7",x"2828",x"3b13",x"3a27"),
(x"2f6d",x"3e2d",x"36eb",x"3776",x"bb0b",x"2d41",x"3a27",x"3a45",x"2f62",x"3e2c",x"36eb",x"3b24",x"371c",x"2cde",x"3a27",x"3a45",x"2f5c",x"3e2c",x"3716",x"3bde",x"b1b5",x"2825",x"3a22",x"3a45"),
(x"2fd6",x"3e7d",x"3715",x"395d",x"39e3",x"2de3",x"3b44",x"38d3",x"2fd9",x"3e7e",x"36eb",x"39df",x"3964",x"2d28",x"3b47",x"38d2",x"3026",x"3e78",x"36eb",x"39ed",x"394b",x"2f45",x"3b46",x"38cf"),
(x"2f3c",x"3e66",x"36eb",x"bbf8",x"2379",x"2d44",x"3b4f",x"38fb",x"2f4a",x"3e66",x"3712",x"bbf7",x"a83f",x"2d8f",x"3b4b",x"38fb",x"2f3f",x"3e64",x"3711",x"bb12",x"3763",x"2ca3",x"3b4b",x"38fb"),
(x"2f3f",x"3e64",x"3711",x"bb12",x"3763",x"2ca3",x"3b4b",x"38fb",x"2f2b",x"3e63",x"36eb",x"b7d8",x"3af6",x"2a35",x"3b4f",x"38fc",x"2f3c",x"3e66",x"36eb",x"bbf8",x"2379",x"2d44",x"3b4f",x"38fb"),
(x"2efb",x"3e3b",x"3713",x"3b5b",x"b634",x"2c08",x"3b41",x"3917",x"2f02",x"3e3a",x"36eb",x"3ad3",x"b822",x"2c4d",x"3b45",x"3917",x"2f01",x"3e39",x"36eb",x"39e9",x"3955",x"2e31",x"3b45",x"3917"),
(x"2fc6",x"3e13",x"36eb",x"bbfe",x"9ea7",x"2828",x"3b13",x"3a27",x"2f8f",x"3e1d",x"36eb",x"bab4",x"b859",x"2a59",x"3b12",x"3a22",x"2f93",x"3e1d",x"370f",x"bad7",x"b821",x"29e6",x"3b0e",x"3a23"),
(x"2f62",x"3e2c",x"36eb",x"3b24",x"371c",x"2cde",x"3a27",x"3a45",x"2f83",x"3e2a",x"36eb",x"397a",x"39b6",x"3099",x"3a27",x"3a44",x"2f72",x"3e29",x"3714",x"39e8",x"3951",x"2f27",x"3a22",x"3a44"),
(x"3026",x"3e78",x"36eb",x"39ed",x"394b",x"2f45",x"3b46",x"38cf",x"3021",x"3e76",x"36eb",x"32cb",x"bbc1",x"2fc5",x"3b45",x"38cf",x"3017",x"3e77",x"3719",x"3250",x"bbca",x"2f22",x"3b42",x"38d1"),
(x"2f3c",x"3e66",x"36eb",x"bbf8",x"2379",x"2d44",x"3b4f",x"38fb",x"2f33",x"3e6a",x"36eb",x"bb57",x"b625",x"2e99",x"3b4f",x"38f9",x"2f3b",x"3e6b",x"3712",x"bb92",x"b509",x"2cb4",x"3b4c",x"38f9"),
(x"2f69",x"3e35",x"36eb",x"3046",x"3be8",x"2cb7",x"3b45",x"3914",x"2f61",x"3e35",x"3713",x"30a8",x"3be9",x"22dc",x"3b42",x"3914",x"2f21",x"3e36",x"3710",x"3833",x"3ac7",x"2d1d",x"3b42",x"3915"),
(x"2f21",x"3e36",x"3710",x"3833",x"3ac7",x"2d1d",x"3b42",x"3915",x"2f01",x"3e39",x"36eb",x"39e9",x"3955",x"2e31",x"3b45",x"3917",x"2f69",x"3e35",x"36eb",x"3046",x"3be8",x"2cb7",x"3b45",x"3914"),
(x"2f93",x"3e1d",x"370f",x"bad7",x"b821",x"29e6",x"3b0e",x"3a23",x"2f8f",x"3e1d",x"36eb",x"bab4",x"b859",x"2a59",x"3b12",x"3a22",x"2f33",x"3e21",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3b11",x"3a1e"),
(x"2f83",x"3e2a",x"36eb",x"397a",x"39b6",x"3099",x"3a27",x"3a44",x"3000",x"3e23",x"36eb",x"3aff",x"373c",x"3197",x"3a27",x"3a3e",x"2fe6",x"3e22",x"3717",x"3a77",x"3889",x"310c",x"3a22",x"3a3e"),
(x"3017",x"3e77",x"3719",x"3250",x"bbca",x"2f22",x"3b42",x"38d1",x"3021",x"3e76",x"36eb",x"32cb",x"bbc1",x"2fc5",x"3b45",x"38cf",x"2fda",x"3e76",x"36eb",x"3b01",x"b745",x"3141",x"3b44",x"38ce"),
(x"2f33",x"3e6a",x"36eb",x"bb57",x"b625",x"2e99",x"3b4f",x"38f9",x"2ea7",x"3e7d",x"36eb",x"bb99",x"b45f",x"30d6",x"3b50",x"38f4",x"2ec5",x"3e7c",x"3711",x"bb70",x"b585",x"3014",x"3b4c",x"38f4"),
(x"2fdf",x"3e37",x"36eb",x"b74a",x"3b15",x"2de4",x"3b46",x"3912",x"2fe6",x"3e36",x"3711",x"b934",x"3a0e",x"2c16",x"3b43",x"3912",x"2fa3",x"3e35",x"3712",x"b2e8",x"3bcb",x"2c10",x"3b42",x"3913"),
(x"2fa3",x"3e35",x"3712",x"b2e8",x"3bcb",x"2c10",x"3b42",x"3913",x"2f69",x"3e35",x"36eb",x"3046",x"3be8",x"2cb7",x"3b45",x"3914",x"2fdf",x"3e37",x"36eb",x"b74a",x"3b15",x"2de4",x"3b46",x"3912"),
(x"2f33",x"3e21",x"36eb",x"b73f",x"bb1a",x"2d3c",x"3b1d",x"3b96",x"2f19",x"3e20",x"36eb",x"38ae",x"ba73",x"2d49",x"3b1d",x"3b95",x"2f20",x"3e21",x"3712",x"3721",x"bb24",x"2bf2",x"3b19",x"3b92"),
(x"3000",x"3e23",x"36eb",x"3aff",x"373c",x"3197",x"3a27",x"3a3e",x"302b",x"3e14",x"36eb",x"3bbf",x"3113",x"322d",x"3a27",x"3a36",x"301b",x"3e14",x"3713",x"3bc6",x"31be",x"30de",x"3a22",x"3a37"),
(x"2ea7",x"3e7d",x"36eb",x"bb99",x"b45f",x"30d6",x"3b50",x"38f4",x"2e7f",x"3e8c",x"36eb",x"bbe6",x"ac77",x"308b",x"3b50",x"38f0",x"2e95",x"3e8c",x"3711",x"bbe4",x"ad1e",x"308c",x"3b4d",x"38f0"),
(x"2fe6",x"3e36",x"3711",x"b934",x"3a0e",x"2c16",x"3b43",x"3912",x"2fdf",x"3e37",x"36eb",x"b74a",x"3b15",x"2de4",x"3b46",x"3912",x"3021",x"3e3d",x"36eb",x"baaf",x"3860",x"2a70",x"3b47",x"3910"),
(x"2f19",x"3e20",x"36eb",x"38ae",x"ba73",x"2d49",x"3b1d",x"3b95",x"2efa",x"3e1e",x"36eb",x"2e29",x"bbe6",x"3005",x"3b1e",x"3b94",x"2ef3",x"3e1f",x"3711",x"35dd",x"bb65",x"2eae",x"3b1a",x"3b91"),
(x"301b",x"3e14",x"3713",x"3bc6",x"31be",x"30de",x"3a22",x"3a37",x"302b",x"3e14",x"36eb",x"3bbf",x"3113",x"322d",x"3a27",x"3a36",x"3025",x"3e07",x"36eb",x"3bea",x"2e09",x"2f12",x"3a26",x"3a2f"),
(x"2fda",x"3e76",x"36eb",x"3b01",x"b745",x"3141",x"3b83",x"3670",x"3006",x"3e73",x"3715",x"39d1",x"3974",x"2cc6",x"3b7e",x"366a",x"2fd8",x"3e76",x"3718",x"3af6",x"37e0",x"2460",x"3b7d",x"366f"),
(x"2fda",x"3e76",x"36eb",x"3b01",x"b745",x"3141",x"3b83",x"3670",x"3016",x"3e72",x"36eb",x"3a0e",x"3929",x"2e76",x"3b83",x"3669",x"3006",x"3e73",x"3715",x"39d1",x"3974",x"2cc6",x"3b7e",x"366a"),
(x"2e95",x"3e8c",x"3711",x"bbe4",x"ad1e",x"308c",x"3b4d",x"38f0",x"2e7f",x"3e8c",x"36eb",x"bbe6",x"ac77",x"308b",x"3b50",x"38f0",x"2e82",x"3e9d",x"36eb",x"bbe8",x"2d66",x"3010",x"3b50",x"38eb"),
(x"3025",x"3e3d",x"3717",x"bb6f",x"35e5",x"261e",x"3b43",x"390f",x"3021",x"3e3d",x"36eb",x"baaf",x"3860",x"2a70",x"3b47",x"3910",x"302e",x"3e45",x"36eb",x"bbfa",x"2c62",x"2617",x"3b48",x"390e"),
(x"2efa",x"3e1e",x"36eb",x"2e29",x"bbe6",x"3005",x"3b1e",x"3b94",x"2e9b",x"3e1f",x"36eb",x"b913",x"ba0d",x"310f",x"3b20",x"3b91",x"2eb1",x"3e20",x"3712",x"b5a6",x"bb63",x"30cc",x"3b1b",x"3b8f"),
(x"3025",x"3e07",x"36eb",x"3bea",x"2e09",x"2f12",x"3a26",x"3a2f",x"303b",x"3dfc",x"36eb",x"3be4",x"2adf",x"30ee",x"3a26",x"3a29",x"3031",x"3dfc",x"370f",x"3bdd",x"30de",x"2e6c",x"3a21",x"3a2a"),
(x"3016",x"3e72",x"36eb",x"3a0e",x"3929",x"2e76",x"3b83",x"3669",x"302e",x"3e6e",x"36eb",x"3bbf",x"3333",x"2ed0",x"3b83",x"3663",x"3022",x"3e6e",x"3718",x"3b13",x"3732",x"2fec",x"3b7d",x"3663"),
(x"2e82",x"3e9d",x"36eb",x"bbe8",x"2d66",x"3010",x"3b50",x"38eb",x"2ea5",x"3ea6",x"36eb",x"bab2",x"3834",x"30cf",x"3b50",x"38e8",x"2eb5",x"3ea5",x"3712",x"bb45",x"3640",x"30a6",x"3b4d",x"38e9"),
(x"2f51",x"3e90",x"3710",x"bb2f",x"b6d9",x"2e52",x"3a13",x"3a56",x"2f41",x"3e90",x"36eb",x"bb02",x"b776",x"2fc8",x"3a17",x"3a57",x"2f36",x"3e94",x"36eb",x"bbf4",x"1edc",x"2eb6",x"3a18",x"3a55"),
(x"302f",x"3e45",x"3715",x"bbfe",x"a412",x"2867",x"3b44",x"390d",x"302e",x"3e45",x"36eb",x"bbfa",x"2c62",x"2617",x"3b48",x"390e",x"3025",x"3e4f",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"3b49",x"390b"),
(x"2e9b",x"3e1f",x"36eb",x"b913",x"ba0d",x"310f",x"3b20",x"3b91",x"2e73",x"3e23",x"36eb",x"bbe5",x"2dbc",x"3036",x"3b20",x"3b8e",x"2e89",x"3e24",x"3711",x"bbb2",x"b32f",x"30f4",x"3b1c",x"3b8d"),
(x"303b",x"3dfc",x"36eb",x"3be4",x"2adf",x"30ee",x"3a26",x"3a29",x"3035",x"3df6",x"36eb",x"3af6",x"b714",x"32f0",x"3a25",x"3a26",x"302a",x"3df8",x"370d",x"3b0d",x"b70c",x"3169",x"3a21",x"3a28"),
(x"302e",x"3e6e",x"36eb",x"3bbf",x"3333",x"2ed0",x"3b83",x"3663",x"302b",x"3e68",x"36eb",x"3bbf",x"b371",x"2dad",x"3b83",x"365d",x"3027",x"3e69",x"3712",x"3bf0",x"ac20",x"2e95",x"3b7e",x"365f"),
(x"2ea5",x"3ea6",x"36eb",x"bab2",x"3834",x"30cf",x"3b50",x"38e8",x"2f13",x"3eae",x"36eb",x"b7cb",x"3ae6",x"3068",x"3b50",x"38e6",x"2f1a",x"3eac",x"3715",x"b93c",x"39e9",x"311d",x"3b4d",x"38e6"),
(x"302a",x"3e50",x"3714",x"bb81",x"b558",x"2da6",x"3b46",x"390a",x"3025",x"3e4f",x"36eb",x"bbcf",x"b2aa",x"2bc5",x"3b49",x"390b",x"3001",x"3e57",x"36eb",x"bac2",x"b833",x"2e85",x"3b4a",x"3909"),
(x"2e73",x"3e23",x"36eb",x"bbe5",x"2dbc",x"3036",x"3b20",x"3b8e",x"2e9a",x"3e2b",x"36eb",x"b902",x"3a23",x"306a",x"3b21",x"3b8a",x"2ea4",x"3e29",x"3712",x"bae4",x"37c3",x"30c9",x"3b1c",x"3b8a"),
(x"302a",x"3df8",x"370d",x"3b0d",x"b70c",x"3169",x"3a21",x"3a28",x"3035",x"3df6",x"36eb",x"3af6",x"b714",x"32f0",x"3a25",x"3a26",x"3020",x"3df5",x"36eb",x"3571",x"bb6d",x"30cc",x"3a25",x"3a25"),
(x"302b",x"3e68",x"36eb",x"3bbf",x"b371",x"2dad",x"3b83",x"365d",x"3025",x"3e67",x"36eb",x"2eda",x"bbea",x"2e47",x"3b83",x"365c",x"301e",x"3e68",x"3712",x"3297",x"bbcc",x"2d84",x"3b7e",x"365d"),
(x"2f13",x"3eae",x"36eb",x"b7cb",x"3ae6",x"3068",x"3b50",x"38e6",x"2f91",x"3eb0",x"36eb",x"96f6",x"3bf5",x"2e99",x"3b50",x"38e3",x"2f91",x"3eaf",x"3715",x"9ef6",x"3bee",x"302a",x"3b4c",x"38e4"),
(x"3008",x"3e58",x"3715",x"ba65",x"b8c1",x"2d9e",x"3b47",x"3908",x"3001",x"3e57",x"36eb",x"bac2",x"b833",x"2e85",x"3b4a",x"3909",x"2fc1",x"3e5c",x"36eb",x"b9cd",x"b979",x"2caa",x"3b4b",x"3907"),
(x"2e9a",x"3e2b",x"36eb",x"b902",x"3a23",x"306a",x"3b21",x"3b8a",x"2ef3",x"3e2c",x"36eb",x"b3f1",x"3bbc",x"2b5c",x"3b22",x"3b87",x"2eea",x"3e2b",x"3713",x"b607",x"3b5e",x"2e4f",x"3b1d",x"3b87"),
(x"301d",x"3df6",x"3713",x"3451",x"bbac",x"2d81",x"3a20",x"3a27",x"3020",x"3df5",x"36eb",x"3571",x"bb6d",x"30cc",x"3a25",x"3a25",x"300a",x"3df5",x"36eb",x"3be3",x"ace8",x"30c3",x"3a24",x"3a23"),
(x"301e",x"3e68",x"3712",x"3297",x"bbcc",x"2d84",x"3b7e",x"365d",x"3025",x"3e67",x"36eb",x"2eda",x"bbea",x"2e47",x"3b83",x"365c",x"2ffe",x"3e67",x"36eb",x"2c58",x"bbf7",x"2bc5",x"3b82",x"3657"),
(x"2f91",x"3eaf",x"3715",x"9ef6",x"3bee",x"302a",x"3b4c",x"38e4",x"2f91",x"3eb0",x"36eb",x"96f6",x"3bf5",x"2e99",x"3b50",x"38e3",x"3007",x"3eae",x"36eb",x"366a",x"3b44",x"2f81",x"3b4f",x"38e1"),
(x"2fc7",x"3e5d",x"3717",x"b939",x"ba0b",x"29e0",x"3b47",x"3906",x"2fc1",x"3e5c",x"36eb",x"b9cd",x"b979",x"2caa",x"3b4b",x"3907",x"2fa3",x"3e5e",x"36eb",x"35a5",x"bb74",x"2d53",x"3b4b",x"3907"),
(x"2eea",x"3e2b",x"3713",x"b607",x"3b5e",x"2e4f",x"3b1d",x"3b87",x"2ef3",x"3e2c",x"36eb",x"b3f1",x"3bbc",x"2b5c",x"3b22",x"3b87",x"2f03",x"3e2d",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3b22",x"3b87"),
(x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4",x"2f27",x"3df7",x"3715",x"19bc",x"26cf",x"3bff",x"385b",x"38c3",x"2f97",x"3e08",x"370e",x"b004",x"271d",x"3bef",x"3860",x"38d8"),
(x"3006",x"3df4",x"3715",x"a58e",x"b07a",x"3beb",x"386a",x"38c2",x"3013",x"3def",x"3712",x"29f0",x"ab1d",x"3bfa",x"386c",x"38bd",x"2f27",x"3df7",x"3715",x"19bc",x"26cf",x"3bff",x"385b",x"38c3"),
(x"2f27",x"3df7",x"3715",x"19bc",x"26cf",x"3bff",x"385b",x"38c3",x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4",x"3006",x"3df4",x"3715",x"a58e",x"b07a",x"3beb",x"386a",x"38c2"),
(x"2f97",x"3e08",x"370e",x"b004",x"271d",x"3bef",x"3860",x"38d8",x"3020",x"3e07",x"3717",x"abf6",x"a5ae",x"3bfb",x"386b",x"38d8",x"3008",x"3df6",x"3716",x"a0ea",x"2786",x"3bfe",x"386a",x"38c4"),
(x"2ffe",x"3e67",x"36eb",x"2c58",x"bbf7",x"2bc5",x"3b82",x"3657",x"2fea",x"3e66",x"36eb",x"3a75",x"b8ad",x"2ccc",x"3b82",x"3655",x"2fe7",x"3e67",x"3716",x"38f4",x"ba42",x"2c09",x"3b7d",x"3657"),
(x"300a",x"3ead",x"3713",x"382e",x"3aba",x"306c",x"3b4c",x"38e2",x"3007",x"3eae",x"36eb",x"366a",x"3b44",x"2f81",x"3b4f",x"38e1",x"3051",x"3ea8",x"36eb",x"39f2",x"3938",x"30b5",x"3b4e",x"38de"),
(x"2f4c",x"3e58",x"36eb",x"3976",x"b9cc",x"2dcc",x"3b4c",x"3905",x"2f4f",x"3e59",x"3714",x"397e",x"b9c5",x"2dbf",x"3b49",x"3904",x"2f79",x"3e5c",x"3714",x"39a7",x"b99f",x"2d1e",x"3b48",x"3905"),
(x"2f79",x"3e5c",x"3714",x"39a7",x"b99f",x"2d1e",x"3b48",x"3905",x"2fa3",x"3e5e",x"36eb",x"35a5",x"bb74",x"2d53",x"3b4b",x"3907",x"2f4c",x"3e58",x"36eb",x"3976",x"b9cc",x"2dcc",x"3b4c",x"3905"),
(x"2f03",x"3e2d",x"36eb",x"b94d",x"b9f2",x"2dc5",x"3b22",x"3b87",x"2ea2",x"3e2e",x"36eb",x"b9ec",x"b92b",x"31e4",x"3b22",x"3b83",x"2ec3",x"3e2f",x"3711",x"b8c8",x"ba4e",x"30a8",x"3b1d",x"3b84"),
(x"3046",x"3ea6",x"3715",x"3ae0",x"37cf",x"30d4",x"3b4b",x"38df",x"3051",x"3ea8",x"36eb",x"39f2",x"3938",x"30b5",x"3b4e",x"38de",x"306a",x"3e9e",x"36eb",x"3bc4",x"327a",x"3012",x"3b4d",x"38dc"),
(x"2f4c",x"3e58",x"36eb",x"3976",x"b9cc",x"2dcc",x"3b4c",x"3905",x"2f11",x"3e55",x"36eb",x"353f",x"bb87",x"2d28",x"3b4d",x"3904",x"2f0c",x"3e56",x"3716",x"37d5",x"baf0",x"2d8e",x"3b4a",x"3903"),
(x"2ea2",x"3e2e",x"36eb",x"b9ec",x"b92b",x"31e4",x"3b22",x"3b83",x"2e56",x"3e37",x"36eb",x"bbbc",x"b212",x"3175",x"3b22",x"3b7e",x"2e71",x"3e37",x"370f",x"bb4b",x"b5cc",x"3223",x"3b1e",x"3b7f"),
(x"3023",x"3def",x"36eb",x"3bdb",x"9c67",x"320a",x"3b13",x"3a55",x"3014",x"3de3",x"36eb",x"3ade",x"b7ab",x"31d3",x"3b16",x"3a50",x"3008",x"3de5",x"370e",x"3b7b",x"b4a9",x"3270",x"3b12",x"3a4e"),
(x"2fda",x"3e66",x"3715",x"3a5f",x"3873",x"3389",x"3a20",x"3a6a",x"3025",x"3e5f",x"36eb",x"3afe",x"375c",x"30f4",x"3a26",x"3a65",x"300d",x"3e5f",x"3718",x"3ac6",x"37dc",x"3286",x"3a20",x"3a66"),
(x"3061",x"3e9d",x"3715",x"3bec",x"2be2",x"2fce",x"3b4a",x"38dc",x"306a",x"3e9e",x"36eb",x"3bc4",x"327a",x"3012",x"3b4d",x"38dc",x"3065",x"3e94",x"36eb",x"3b6e",x"b575",x"309e",x"3b4c",x"38d9"),
(x"2f2f",x"3e80",x"3714",x"b05e",x"a194",x"3bec",x"3856",x"3961",x"2e95",x"3e8c",x"3711",x"acd1",x"a504",x"3bf9",x"384b",x"396e",x"2ed8",x"3e8e",x"3713",x"b0f4",x"9987",x"3be7",x"3850",x"3970"),
(x"2f2f",x"3e80",x"3714",x"b05e",x"a194",x"3bec",x"3856",x"3961",x"2ec5",x"3e7c",x"3711",x"b115",x"a7d5",x"3be4",x"384f",x"395c",x"2e95",x"3e8c",x"3711",x"acd1",x"a504",x"3bf9",x"384b",x"396e"),
(x"2f11",x"3e55",x"36eb",x"353f",x"bb87",x"2d28",x"3b4d",x"3904",x"2ec4",x"3e54",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"3b4d",x"3902",x"2ecb",x"3e55",x"3716",x"a345",x"bbf7",x"2dcc",x"3b4a",x"3901"),
(x"2e56",x"3e37",x"36eb",x"bbbc",x"b212",x"3175",x"3b22",x"3b7e",x"2e52",x"3e41",x"36eb",x"bb61",x"35a0",x"3119",x"3b22",x"3b79",x"2e69",x"3e40",x"370f",x"bbd3",x"2f46",x"3182",x"3b1d",x"3b7a"),
(x"3025",x"3e5f",x"36eb",x"3afe",x"375c",x"30f4",x"3a26",x"3a65",x"304c",x"3e53",x"36eb",x"3bba",x"3376",x"2f14",x"3a26",x"3a5f",x"3041",x"3e53",x"3714",x"3b6b",x"3587",x"3096",x"3a21",x"3a5f"),
(x"3065",x"3e94",x"36eb",x"3b6e",x"b575",x"309e",x"3b4c",x"38d9",x"303a",x"3e8d",x"36eb",x"3884",x"ba69",x"324a",x"3b4b",x"38d7",x"3030",x"3e8e",x"3711",x"38a4",x"ba69",x"309a",x"3b48",x"38d8"),
(x"2ec4",x"3e54",x"36eb",x"b3e5",x"bbb4",x"2ec2",x"3b4d",x"3902",x"2e81",x"3e56",x"36eb",x"bacb",x"b812",x"3065",x"3b4e",x"3901",x"2e97",x"3e57",x"3714",x"b976",x"b9c0",x"3023",x"3b4b",x"3901"),
(x"2e52",x"3e41",x"36eb",x"bb61",x"35a0",x"3119",x"3b22",x"3b79",x"2e9d",x"3e47",x"36eb",x"b86e",x"3a87",x"313e",x"3b21",x"3b75",x"2ea1",x"3e45",x"370f",x"b891",x"3a72",x"30f5",x"3b1d",x"3b77"),
(x"3014",x"3de3",x"36eb",x"3ade",x"b7ab",x"31d3",x"3b16",x"3a50",x"2fa3",x"3dd9",x"36eb",x"38a6",x"ba54",x"3207",x"3b18",x"3a49",x"2fa8",x"3ddc",x"3712",x"38b5",x"ba3e",x"32bd",x"3b13",x"3a49"),
(x"304c",x"3e53",x"36eb",x"3bba",x"3376",x"2f14",x"3a26",x"3a5f",x"305b",x"3e46",x"36eb",x"3bef",x"ad09",x"2e69",x"3a27",x"3a58",x"3052",x"3e47",x"3712",x"3bf0",x"2a00",x"2f46",x"3a22",x"3a58"),
(x"3030",x"3e8e",x"3711",x"38a4",x"ba69",x"309a",x"3b48",x"38d8",x"303a",x"3e8d",x"36eb",x"3884",x"ba69",x"324a",x"3b4b",x"38d7",x"2fed",x"3e8b",x"36eb",x"360d",x"bb5a",x"2ef3",x"3b49",x"38d5"),
(x"2e81",x"3e56",x"36eb",x"bacb",x"b812",x"3065",x"3b4e",x"3901",x"2e6a",x"3e5c",x"36eb",x"bbcf",x"3174",x"3043",x"3b4e",x"3900",x"2e81",x"3e5b",x"3712",x"bbe0",x"ae5e",x"30a3",x"3b4b",x"38ff"),
(x"2ea1",x"3e45",x"370f",x"b891",x"3a72",x"30f5",x"3b1d",x"3b77",x"2e9d",x"3e47",x"36eb",x"b86e",x"3a87",x"313e",x"3b21",x"3b75",x"2efa",x"3e48",x"36eb",x"35e4",x"3b4d",x"31a2",x"3b21",x"3b72"),
(x"2fa8",x"3ddc",x"3712",x"38b5",x"ba3e",x"32bd",x"3b13",x"3a49",x"2fa3",x"3dd9",x"36eb",x"38a6",x"ba54",x"3207",x"3b18",x"3a49",x"2f52",x"3dd9",x"36eb",x"b996",x"b95e",x"33ec",x"3b19",x"3a47"),
(x"305b",x"3e46",x"36eb",x"3bef",x"ad09",x"2e69",x"3a27",x"3a58",x"3046",x"3e3a",x"36eb",x"3b75",x"b5a2",x"2d46",x"3a27",x"3a52",x"3041",x"3e3b",x"3710",x"3b6a",x"b5bb",x"2efe",x"3a23",x"3a52"),
(x"2fe3",x"3e8b",x"3718",x"38ae",x"ba78",x"2b79",x"3b46",x"38d6",x"2fed",x"3e8b",x"36eb",x"360d",x"bb5a",x"2ef3",x"3b49",x"38d5",x"2fd8",x"3e89",x"36eb",x"3be6",x"b08e",x"2c41",x"3b49",x"38d4"),
(x"2e6a",x"3e5c",x"36eb",x"bbcf",x"3174",x"3043",x"3b4e",x"3900",x"2e90",x"3e61",x"36eb",x"b6fe",x"3b25",x"2ea4",x"3b4e",x"38fe",x"2e99",x"3e5f",x"3714",x"b972",x"39bb",x"30de",x"3b4b",x"38fe"),
(x"2ec4",x"3e97",x"3710",x"2828",x"a60a",x"3bfe",x"384e",x"397a",x"2ed8",x"3e8e",x"3713",x"b0f4",x"9987",x"3be7",x"3850",x"3970",x"2e95",x"3e8c",x"3711",x"acd1",x"a504",x"3bf9",x"384b",x"396e"),
(x"2e95",x"3e9d",x"3714",x"2eb0",x"a8fa",x"3bf3",x"384b",x"3981",x"2eca",x"3e9e",x"3714",x"2946",x"9ffc",x"3bfe",x"384e",x"3982",x"2ec4",x"3e97",x"3710",x"2828",x"a60a",x"3bfe",x"384e",x"397a"),
(x"2eb5",x"3ea5",x"3712",x"a587",x"a08e",x"3bff",x"384c",x"398a",x"2eca",x"3e9e",x"3714",x"2946",x"9ffc",x"3bfe",x"384e",x"3982",x"2e95",x"3e9d",x"3714",x"2eb0",x"a8fa",x"3bf3",x"384b",x"3981"),
(x"2eb5",x"3ea5",x"3712",x"a587",x"a08e",x"3bff",x"384c",x"398a",x"2edf",x"3ea3",x"3712",x"2953",x"a7ae",x"3bfd",x"384f",x"3987",x"2eca",x"3e9e",x"3714",x"2946",x"9ffc",x"3bfe",x"384e",x"3982"),
(x"2f1a",x"3eac",x"3715",x"a0ea",x"aafd",x"3bfc",x"3853",x"3993",x"2f3d",x"3ea8",x"3714",x"231d",x"ab5f",x"3bfc",x"3855",x"398e",x"2f06",x"3ea6",x"3714",x"a8bf",x"ac22",x"3bfa",x"3852",x"398b"),
(x"2f91",x"3eaf",x"3715",x"27db",x"a9b2",x"3bfc",x"385a",x"3996",x"2fa3",x"3eaa",x"3715",x"270a",x"2779",x"3bfe",x"385c",x"3991",x"2f3d",x"3ea8",x"3714",x"231d",x"ab5f",x"3bfc",x"3855",x"398e"),
(x"300a",x"3ead",x"3713",x"2b1d",x"2ee4",x"3bf0",x"3863",x"3994",x"3004",x"3ea9",x"3716",x"24bc",x"2ceb",x"3bf9",x"3862",x"3990",x"2fa3",x"3eaa",x"3715",x"270a",x"2779",x"3bfe",x"385c",x"3991"),
(x"3046",x"3ea6",x"3715",x"a266",x"1d87",x"3bff",x"386b",x"398d",x"302c",x"3ea3",x"3714",x"a8e0",x"a99e",x"3bfc",x"3868",x"3989",x"3004",x"3ea9",x"3716",x"24bc",x"2ceb",x"3bf9",x"3862",x"3990"),
(x"3061",x"3e9d",x"3715",x"a891",x"27ce",x"3bfd",x"386f",x"3983",x"3036",x"3e9d",x"3714",x"a538",x"29ab",x"3bfd",x"386a",x"3983",x"302c",x"3ea3",x"3714",x"a8e0",x"a99e",x"3bfc",x"3868",x"3989"),
(x"3061",x"3e9d",x"3715",x"a891",x"27ce",x"3bfd",x"386f",x"3983",x"3058",x"3e95",x"3717",x"ad06",x"a793",x"3bf8",x"386f",x"397a",x"3026",x"3e98",x"3715",x"ac67",x"a8a5",x"3bf9",x"3868",x"397d"),
(x"3030",x"3e8e",x"3711",x"a8d9",x"252b",x"3bfe",x"386a",x"3972",x"3006",x"3e98",x"3714",x"aa45",x"ab10",x"3bfa",x"3864",x"397c",x"3026",x"3e98",x"3715",x"ac67",x"a8a5",x"3bf9",x"3868",x"397d"),
(x"2f5e",x"3e98",x"3711",x"abef",x"28a8",x"3bfa",x"3858",x"397c",x"2f85",x"3e9a",x"3710",x"a352",x"2e80",x"3bf5",x"385b",x"397f",x"2fd7",x"3e9a",x"3711",x"aa66",x"331a",x"3bca",x"3860",x"397f"),
(x"2f89",x"3e8c",x"3713",x"b41f",x"2c3a",x"3bb6",x"385b",x"396e",x"2f73",x"3e8e",x"3711",x"b40c",x"a6c2",x"3bbc",x"385a",x"3970",x"2fe3",x"3e8b",x"3718",x"ab65",x"3528",x"3b8f",x"3862",x"396d"),
(x"2f8e",x"3e87",x"3714",x"ade0",x"24c2",x"3bf6",x"385c",x"3969",x"2fcc",x"3e88",x"3718",x"b420",x"9418",x"3bba",x"3860",x"396a",x"2fc7",x"3e7f",x"3715",x"a7ae",x"24ea",x"3bfe",x"3860",x"395f"),
(x"2f8e",x"3e87",x"3714",x"ade0",x"24c2",x"3bf6",x"385c",x"3969",x"2f89",x"3e8c",x"3713",x"b41f",x"2c3a",x"3bb6",x"385b",x"396e",x"2fcc",x"3e88",x"3718",x"b420",x"9418",x"3bba",x"3860",x"396a"),
(x"2f5e",x"3e98",x"3711",x"abef",x"28a8",x"3bfa",x"3858",x"397c",x"2f51",x"3e90",x"3710",x"a856",x"29ab",x"3bfc",x"3858",x"3973",x"2f45",x"3e94",x"3710",x"aa8d",x"a973",x"3bfb",x"3857",x"3978"),
(x"3006",x"3e98",x"3714",x"aa45",x"ab10",x"3bfa",x"3864",x"397c",x"3030",x"3e8e",x"3711",x"a8d9",x"252b",x"3bfe",x"386a",x"3972",x"2f51",x"3e90",x"3710",x"a856",x"29ab",x"3bfc",x"3858",x"3973"),
(x"2f82",x"3e8c",x"36eb",x"bbf6",x"aa70",x"2d60",x"3a17",x"3a5a",x"2f89",x"3e8c",x"3713",x"bbc2",x"b3a4",x"298a",x"3a12",x"3a59",x"2f8e",x"3e87",x"3714",x"bbf3",x"2e23",x"2b27",x"3a11",x"3a5b"),
(x"2f8e",x"3e87",x"3714",x"bbf3",x"2e23",x"2b27",x"3a11",x"3a5b",x"2f6c",x"3e7b",x"36eb",x"b46a",x"3b91",x"316a",x"3a15",x"3a63",x"2f82",x"3e8c",x"36eb",x"bbf6",x"aa70",x"2d60",x"3a17",x"3a5a"),
(x"3a25",x"4041",x"3710",x"3bd6",x"2604",x"3256",x"39c5",x"33c0",x"3a26",x"4036",x"3710",x"3bcf",x"2680",x"32dc",x"39b2",x"33ca",x"3a20",x"4036",x"3732",x"3b18",x"2439",x"3763",x"39b1",x"33aa"),
(x"3a1f",x"4041",x"3733",x"3b23",x"251e",x"3738",x"39c4",x"339f",x"3a20",x"4036",x"3732",x"3b18",x"2439",x"3763",x"39b1",x"33aa",x"3a19",x"4036",x"3749",x"3871",x"2587",x"3aa6",x"39b0",x"3392"),
(x"3a18",x"4041",x"3748",x"36c9",x"29dc",x"3b3c",x"39c4",x"3388",x"3a19",x"4036",x"3749",x"3871",x"2587",x"3aa6",x"39b0",x"3392",x"3a14",x"4036",x"374e",x"2fa2",x"2997",x"3bef",x"39b0",x"3387"),
(x"3a10",x"4041",x"3749",x"b4de",x"2b76",x"3b9b",x"39c3",x"337b",x"3a14",x"4036",x"374e",x"2fa2",x"2997",x"3bef",x"39b0",x"3387",x"3a0d",x"4036",x"374b",x"b745",x"2966",x"3b1e",x"39b0",x"337b"),
(x"3a09",x"4041",x"373b",x"b7a6",x"3a67",x"35ca",x"3b1c",x"3899",x"39fc",x"4042",x"3713",x"af5f",x"3bdb",x"30c1",x"3b21",x"38a0",x"3a03",x"4042",x"370e",x"ae5c",x"3b3a",x"36a9",x"3b1f",x"38a1"),
(x"3a09",x"4042",x"373a",x"baf6",x"2b34",x"37d2",x"3b1b",x"3899",x"3a11",x"4042",x"374a",x"b548",x"b37f",x"3b50",x"3b18",x"3896",x"3a10",x"4041",x"3749",x"b3ab",x"a4bc",x"3bc3",x"3b1a",x"3895"),
(x"39fc",x"4036",x"3710",x"ba72",x"9a8d",x"38bc",x"39b0",x"333e",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e",x"3a02",x"4036",x"3724",x"bb1f",x"1a24",x"3747",x"39b0",x"3352"),
(x"3a02",x"404d",x"3711",x"bbe1",x"a6cf",x"3179",x"3bfb",x"399f",x"3a04",x"404d",x"3727",x"bbc5",x"a901",x"3377",x"3bfb",x"39a3",x"3a03",x"4042",x"370e",x"bbc2",x"ab4f",x"338c",x"3bea",x"399f"),
(x"3a08",x"404d",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"39a7",x"3a0f",x"404d",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"39ab",x"3a11",x"4042",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"39ac"),
(x"3a0f",x"404d",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"39ab",x"3a17",x"404d",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3bfc",x"39af",x"3a19",x"4043",x"374d",x"3400",x"aa73",x"3bbc",x"3bec",x"39af"),
(x"3a1d",x"404d",x"374d",x"3802",x"a90b",x"3aea",x"3bfc",x"39b1",x"3a21",x"4043",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"39b3",x"3a19",x"4043",x"374d",x"3400",x"aa73",x"3bbc",x"3bec",x"39af"),
(x"3a24",x"404d",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"39b5",x"3a25",x"4043",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"39b6",x"3a21",x"4043",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"39b3"),
(x"3a2a",x"404d",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"39ba",x"3a2d",x"4042",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"39be",x"3a25",x"4043",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"39b6"),
(x"3a2d",x"4042",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"39be",x"3a2a",x"404d",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"39ba",x"3a2f",x"404d",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"39bf"),
(x"3a25",x"4043",x"3738",x"36f3",x"bae7",x"3422",x"3b16",x"388d",x"3a2d",x"4042",x"3710",x"3644",x"bb4c",x"2f83",x"3b19",x"3884",x"3a25",x"4041",x"3710",x"3700",x"bb23",x"2f05",x"3b1b",x"3887"),
(x"3a0d",x"4036",x"374b",x"b745",x"2966",x"3b1e",x"39b0",x"337b",x"3a07",x"4036",x"373c",x"bac4",x"2853",x"3841",x"39b0",x"336a",x"3a09",x"4041",x"373b",x"b9d7",x"2404",x"3976",x"39c3",x"3369"),
(x"3a11",x"4042",x"374a",x"b548",x"b37f",x"3b50",x"3b18",x"3896",x"3a19",x"4043",x"374d",x"3243",x"b807",x"3aba",x"3b16",x"3893",x"3a18",x"4041",x"3748",x"2918",x"b8de",x"3a57",x"3b18",x"3893"),
(x"3a18",x"4041",x"3748",x"2918",x"b8de",x"3a57",x"3b18",x"3893",x"3a19",x"4043",x"374d",x"3243",x"b807",x"3aba",x"3b16",x"3893",x"3a21",x"4043",x"3744",x"37e0",x"ba17",x"36be",x"3b16",x"388f"),
(x"3a25",x"4043",x"3738",x"36f3",x"bae7",x"3422",x"3b16",x"388d",x"3a1f",x"4041",x"3733",x"37fe",x"ba99",x"3438",x"3b19",x"388d",x"3a21",x"4043",x"3744",x"37e0",x"ba17",x"36be",x"3b16",x"388f"),
(x"3a2a",x"404d",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3821",x"3a20",x"404d",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3827",x"3a26",x"404d",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3820"),
(x"3a24",x"404d",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3826",x"3a1a",x"404d",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"382b",x"3a20",x"404d",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3827"),
(x"3a1d",x"404d",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"382a",x"3a15",x"404d",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"382d",x"3a1a",x"404d",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"382b"),
(x"3a17",x"404d",x"3751",x"2fd8",x"39a6",x"3994",x"3b24",x"382d",x"3a15",x"404d",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"382d",x"3a1d",x"404d",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"382a"),
(x"3a0f",x"404d",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3830",x"3a0f",x"404e",x"3749",x"b6e3",x"3561",x"3ab3",x"3b21",x"382f",x"3a15",x"404d",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"382d"),
(x"3a08",x"404d",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3832",x"3a09",x"404e",x"373e",x"ba28",x"9df0",x"391a",x"3b1e",x"3831",x"3a0f",x"404e",x"3749",x"b6e3",x"3561",x"3ab3",x"3b21",x"382f"),
(x"3a04",x"404d",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3835",x"3a01",x"404d",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3835",x"3a09",x"404e",x"373e",x"ba28",x"9df0",x"391a",x"3b1e",x"3831"),
(x"3a02",x"404d",x"3711",x"b40e",x"bb3a",x"3585",x"3b18",x"3838",x"3a01",x"404d",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3835",x"3a04",x"404d",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3835"),
(x"3a02",x"404d",x"3711",x"b40e",x"bb3a",x"3585",x"3b18",x"3838",x"39fb",x"404d",x"3713",x"aedc",x"bb7b",x"3565",x"3b16",x"3836",x"3a01",x"404d",x"371c",x"b97c",x"b976",x"340b",x"3b19",x"3835"),
(x"3a02",x"404d",x"3711",x"315a",x"2bae",x"3bdf",x"39d6",x"3349",x"3a03",x"4042",x"370e",x"34eb",x"a6e9",x"3b9c",x"39c4",x"334b",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e"),
(x"3a24",x"4059",x"372b",x"3b86",x"a8a8",x"3564",x"39eb",x"33b1",x"3a27",x"4059",x"3710",x"3bea",x"a4d6",x"30a2",x"39ea",x"33c9",x"3a26",x"404d",x"3710",x"3bed",x"a7ae",x"3024",x"39d7",x"33c4"),
(x"3a24",x"4059",x"372b",x"3b86",x"a8a8",x"3564",x"39eb",x"33b1",x"3a20",x"404d",x"3739",x"3abd",x"a8b5",x"384c",x"39d7",x"339e",x"3a21",x"4059",x"373a",x"3acd",x"a5ae",x"3834",x"39eb",x"33a3"),
(x"3a20",x"404d",x"3739",x"3abd",x"a8b5",x"384c",x"39d7",x"339e",x"3a1a",x"404d",x"3746",x"38a5",x"a839",x"3a81",x"39d8",x"338e",x"3a1a",x"4059",x"3749",x"38cd",x"a812",x"3a64",x"39eb",x"3391"),
(x"3a15",x"404d",x"374b",x"2e57",x"a8d3",x"3bf4",x"39d8",x"3385",x"3a14",x"4059",x"374f",x"32be",x"a89e",x"3bd0",x"39eb",x"3384",x"3a1a",x"4059",x"3749",x"38cd",x"a812",x"3a64",x"39eb",x"3391"),
(x"3a0f",x"404e",x"3749",x"b771",x"a91b",x"3b13",x"39d8",x"3379",x"3a0d",x"4059",x"374b",x"b6cb",x"a758",x"3b3d",x"39eb",x"3378",x"3a14",x"4059",x"374f",x"32be",x"a89e",x"3bd0",x"39eb",x"3384"),
(x"3a09",x"404e",x"373e",x"ba21",x"a786",x"3921",x"39d8",x"336a",x"3a07",x"4059",x"373c",x"baa0",x"a6bb",x"3879",x"39eb",x"3366",x"3a0d",x"4059",x"374b",x"b6cb",x"a758",x"3b3d",x"39eb",x"3378"),
(x"3a09",x"404e",x"373e",x"ba21",x"a786",x"3921",x"39d8",x"336a",x"3a01",x"404d",x"371c",x"b9f4",x"a495",x"3957",x"39d7",x"334a",x"3a00",x"4059",x"3722",x"ba6c",x"a860",x"38c2",x"39ea",x"334c"),
(x"3a01",x"404d",x"371c",x"b9f4",x"a495",x"3957",x"39d7",x"334a",x"39fb",x"404d",x"3713",x"a9a8",x"a460",x"3bfd",x"39d7",x"333d",x"39fc",x"4059",x"3718",x"b8fc",x"a86a",x"3a40",x"39eb",x"3340"),
(x"3475",x"404a",x"3710",x"0000",x"0000",x"3c00",x"39d1",x"2450",x"3485",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"24c1",x"3485",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"24c1"),
(x"3485",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"24c1",x"3485",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"24c1",x"349b",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"255f"),
(x"349b",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"255f",x"349b",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"255f",x"34bb",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2642"),
(x"34bb",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2642",x"34cb",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"26b3",x"34cb",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"26b3"),
(x"34cb",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"26b3",x"34cb",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"26b3",x"34e9",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"278b"),
(x"34e9",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"278b",x"3501",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"281a",x"3501",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"281a"),
(x"3501",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"281a",x"351b",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"2878",x"351b",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39be",x"2878"),
(x"351b",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"2878",x"353f",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"28fa",x"353f",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"28fa"),
(x"353f",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"28fa",x"353f",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"28fa",x"3555",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2949"),
(x"3555",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2949",x"357d",x"404b",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"29d7",x"357d",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"29d7"),
(x"357d",x"404b",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"29d7",x"3592",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"2a20",x"3592",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2a20"),
(x"36f7",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2d8d",x"363b",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2c3f",x"363b",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2c3f"),
(x"363b",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2c3f",x"363b",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2c3f",x"362c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2c23"),
(x"362c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2c23",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b"),
(x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b",x"3592",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2a20",x"3592",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"2a20"),
(x"35f5",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2b83",x"35fd",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"2ba0",x"35fd",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2ba0"),
(x"35e4",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2b47",x"35fd",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2ba0",x"35f3",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2b7d"),
(x"35d3",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"2b0a",x"35f3",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2b7d",x"35f1",x"4052",x"3710",x"0000",x"0000",x"3c00",x"39df",x"2b76"),
(x"35f5",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2b83",x"35e4",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2b47",x"35fd",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2ba0"),
(x"35e4",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2b47",x"35d3",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2b0a",x"35f3",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2b7d"),
(x"35d3",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2b0a",x"35bd",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"2ab9",x"35f1",x"403d",x"3710",x"868d",x"8cea",x"3c00",x"39bb",x"2b76"),
(x"35bd",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"2ab9",x"359e",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2a4d",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b"),
(x"35bd",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2ab9",x"35f1",x"4052",x"3710",x"0000",x"0000",x"3c00",x"39df",x"2b76",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b"),
(x"359e",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2a4d",x"358a",x"403d",x"3710",x"0000",x"0000",x"3c00",x"39bb",x"2a0d",x"3593",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2a27"),
(x"3593",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2a24",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b",x"3592",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"2a20"),
(x"36f7",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2d8d",x"36f7",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2d8d",x"3710",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2dbb"),
(x"380a",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2f8b",x"37b8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2ee7",x"37b8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ee7"),
(x"37b8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ee7",x"37b8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2ee7",x"37a8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2ec9"),
(x"37a8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2ec9",x"378c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2e97",x"378c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2e97"),
(x"378c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2e97",x"378c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2e97",x"376c",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"2e5e"),
(x"376c",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"2e5e",x"3752",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2e30",x"3752",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2e30"),
(x"36f7",x"405b",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e",x"3716",x"405a",x"3710",x"0000",x"0000",x"3c00",x"39ed",x"2dc4",x"36df",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"2d63"),
(x"3716",x"405a",x"3710",x"0000",x"0000",x"3c00",x"39ed",x"2dc4",x"372e",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2df0",x"36dc",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2d5e"),
(x"36df",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"2d63",x"3716",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ad",x"2dc4",x"36f7",x"4034",x"3710",x"0000",x"0000",x"3c00",x"39ac",x"2d8e"),
(x"36dc",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2d5e",x"372e",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2df0",x"3716",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ad",x"2dc4"),
(x"3753",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b0",x"2e32",x"3742",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2e14",x"375f",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2e47"),
(x"3742",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2e14",x"372e",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2df0",x"3754",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"2e33"),
(x"3753",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39ea",x"2e32",x"3760",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e7",x"2e49",x"375f",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e4",x"2e47"),
(x"3742",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2e14",x"375f",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e4",x"2e47",x"3754",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"2e33"),
(x"36cb",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2d3f",x"36c2",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"2d2f",x"36c4",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"2d33"),
(x"36cb",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39be",x"2d3f",x"3705",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"2da6",x"36c4",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"2d33"),
(x"3705",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"2da6",x"3713",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"2dbf",x"36dc",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2d5e"),
(x"3705",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"2da6",x"36c4",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"2d33",x"36dc",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2d5e"),
(x"3713",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2dbf",x"36dc",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2d5e",x"372e",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2df0"),
(x"372e",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2df0",x"36dc",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2d5e",x"3713",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"2dbf"),
(x"3713",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2dbf",x"3754",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"2e33",x"3752",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2e30"),
(x"3713",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"2dbf",x"3716",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2dc5",x"3752",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2e30"),
(x"3710",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2dbb",x"3710",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2dbb",x"3716",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2dc5"),
(x"3716",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2dc5",x"3752",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2e30",x"3752",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2e30"),
(x"3813",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2fac",x"3813",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2fac",x"380a",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2f8b"),
(x"382a",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2ffc",x"382a",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2ffc",x"3813",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2fac"),
(x"3885",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30a2",x"3885",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30a2",x"382a",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2ffc"),
(x"3885",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30a2",x"388c",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30ad",x"388c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30ad"),
(x"38bf",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"3109",x"38bf",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"3109",x"38d5",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"3130"),
(x"38bf",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"3109",x"38b2",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"30f1",x"38b2",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"30f1"),
(x"38b2",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"30f1",x"38b0",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"30ed",x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed"),
(x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed",x"38b0",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"30ed",x"388c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30ad"),
(x"3872",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"3080",x"3877",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3088",x"386d",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3076"),
(x"3885",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"30a2",x"3894",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ae",x"30bc",x"3877",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3088"),
(x"386d",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3076",x"3877",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3088",x"3872",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"3080"),
(x"3877",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3088",x"3894",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39ec",x"30bc",x"3885",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"30a2"),
(x"3894",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39ec",x"30bc",x"38b7",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"30f9",x"388c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"30ae"),
(x"388c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"30ae",x"38b7",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"30f9",x"3894",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ae",x"30bc"),
(x"38d8",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3135",x"38c7",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"3117",x"38d4",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"312d"),
(x"38d8",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3135",x"38d9",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e4",x"3136",x"38d4",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"312d"),
(x"38c7",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"3117",x"38d4",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"312d",x"38c9",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"311a"),
(x"38c7",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"3117",x"38b7",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"30f9",x"38c9",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"311a"),
(x"388c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"30ae",x"388c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30ad",x"38b0",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"30ed"),
(x"388c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"30ae",x"38b2",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"30f2",x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed"),
(x"38b2",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"30f2",x"38b7",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"30f9",x"388c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"30ae"),
(x"38b7",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"30f9",x"38b2",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"30f2",x"388c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"30ae"),
(x"38c9",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"311a",x"38b7",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"30f9",x"38bd",x"403d",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"3107"),
(x"38b2",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"30f2",x"38b7",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"30f9",x"38bd",x"4052",x"3710",x"0000",x"0000",x"3c00",x"39de",x"3107"),
(x"38f6",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"316b",x"38f6",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"316b",x"38d5",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"3130"),
(x"38f6",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"316b",x"3915",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"31a2",x"3915",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"31a2"),
(x"392f",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"31d0",x"392f",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"31d0",x"3915",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"31a2"),
(x"393f",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"31ed",x"393f",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"31ed",x"392f",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"31d0"),
(x"3953",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3211",x"3953",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3211",x"393f",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"31ed"),
(x"3953",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3211",x"395a",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"321d",x"395a",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"321d"),
(x"395d",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"3222",x"395d",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"3222",x"395a",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"321d"),
(x"395d",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"3222",x"3963",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"322d",x"3963",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"322d"),
(x"3972",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"3248",x"3972",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"3248",x"3963",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"322d"),
(x"3985",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3269",x"3985",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3269",x"3972",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"3248"),
(x"3985",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3269",x"3994",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3284",x"3994",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3284"),
(x"3999",x"4058",x"3710",x"935f",x"1e0a",x"3c00",x"39e9",x"328d",x"3999",x"4037",x"3710",x"975f",x"9f93",x"3c00",x"39b1",x"328d",x"3994",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3284"),
(x"3999",x"4058",x"3710",x"935f",x"1e0a",x"3c00",x"39e9",x"328d",x"39fb",x"404d",x"3713",x"a9a8",x"a460",x"3bfd",x"39d7",x"333d",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e"),
(x"39f5",x"4059",x"3710",x"b60b",x"25b5",x"3b67",x"39eb",x"3331",x"39fc",x"4059",x"3718",x"b8fc",x"a86a",x"3a40",x"39eb",x"3340",x"39fb",x"404d",x"3713",x"a9a8",x"a460",x"3bfd",x"39d7",x"333d"),
(x"3999",x"4037",x"3710",x"975f",x"9f93",x"3c00",x"39b1",x"328d",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e",x"39fc",x"4036",x"3710",x"ba72",x"9a8d",x"38bc",x"39b0",x"333e"),
(x"3a0d",x"4059",x"374b",x"a412",x"3bfd",x"295c",x"3a18",x"3ba9",x"3a07",x"4059",x"373c",x"a752",x"3bff",x"9bfc",x"3a1b",x"3ba6",x"3a1a",x"4059",x"3749",x"a2b5",x"3bfe",x"281b",x"3a18",x"3bae"),
(x"3a07",x"4059",x"373c",x"a752",x"3bff",x"9bfc",x"3a1b",x"3ba6",x"3a00",x"4059",x"3722",x"23fc",x"3bf8",x"2d58",x"3a1f",x"3ba4",x"3a21",x"4059",x"373a",x"a884",x"3bfe",x"253f",x"3a1b",x"3bb1"),
(x"3a00",x"4059",x"3722",x"23fc",x"3bf8",x"2d58",x"3a1f",x"3ba4",x"39fc",x"4059",x"3718",x"135f",x"3bfd",x"29a5",x"3a21",x"3ba2",x"3a24",x"4059",x"372b",x"a504",x"3bff",x"9a59",x"3a1e",x"3bb2"),
(x"39fc",x"4059",x"3718",x"135f",x"3bfd",x"29a5",x"3a21",x"3ba2",x"39f5",x"4059",x"3710",x"a4e3",x"3bff",x"1818",x"3a23",x"3b9f",x"3a27",x"4059",x"3710",x"a3ef",x"3bff",x"9818",x"3a23",x"3bb3"),
(x"3a19",x"4036",x"3749",x"208e",x"bc00",x"135f",x"3a12",x"3bab",x"3a07",x"4036",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a0f",x"3ba4",x"3a0d",x"4036",x"374b",x"1481",x"bbff",x"26ae",x"3a12",x"3ba6"),
(x"3a20",x"4036",x"3732",x"1f93",x"bc00",x"975f",x"3a0d",x"3bae",x"3a02",x"4036",x"3724",x"1c81",x"bbff",x"a1c9",x"3a0b",x"3ba2",x"3a07",x"4036",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a0f",x"3ba4"),
(x"3a26",x"4036",x"3710",x"1f45",x"bbff",x"a032",x"3a07",x"3bb0",x"39fc",x"4036",x"3710",x"9bc8",x"bc00",x"200b",x"3a07",x"3b9f",x"3a02",x"4036",x"3724",x"1c81",x"bbff",x"a1c9",x"3a0b",x"3ba2"),
(x"34e9",x"403f",x"36da",x"b698",x"bb49",x"8000",x"3a50",x"3b8e",x"34e9",x"403f",x"3710",x"b50d",x"bb97",x"0000",x"3a5a",x"3b8e",x"3501",x"403e",x"3710",x"2d0c",x"bbf9",x"0000",x"3a5a",x"3b93"),
(x"3872",x"403e",x"36da",x"b902",x"3a3c",x"0000",x"3a72",x"3ad4",x"3872",x"403e",x"3710",x"b9d1",x"397d",x"8000",x"3a7c",x"3ad4",x"386c",x"403c",x"3710",x"bbdd",x"31e1",x"0000",x"3a7c",x"3ad8"),
(x"3813",x"404e",x"36da",x"27fc",x"3bfe",x"0000",x"3a8b",x"3b47",x"3813",x"404e",x"3710",x"a8bf",x"3bfe",x"8000",x"3a96",x"3b47",x"380a",x"404d",x"3710",x"ae11",x"3bf6",x"0000",x"3a96",x"3b4a"),
(x"34cb",x"4041",x"36da",x"b501",x"bb99",x"0000",x"3a50",x"3b87",x"34cb",x"4041",x"3710",x"b64c",x"bb5a",x"0000",x"3a5a",x"3b87",x"34e9",x"403f",x"3710",x"b50d",x"bb97",x"0000",x"3a5a",x"3b8e"),
(x"39fc",x"4036",x"36da",x"a111",x"bc00",x"0000",x"39fd",x"3b9f",x"39fc",x"4036",x"3710",x"9bc8",x"bc00",x"200b",x"3a07",x"3b9f",x"3a26",x"4036",x"3710",x"1f45",x"bbff",x"a032",x"3a07",x"3bb0"),
(x"3885",x"4040",x"36da",x"b83d",x"3ac8",x"0000",x"3a72",x"3acc",x"3885",x"4040",x"3710",x"b7eb",x"3af3",x"0000",x"3a7c",x"3acc",x"3872",x"403e",x"3710",x"b9d1",x"397d",x"8000",x"3a7c",x"3ad4"),
(x"375f",x"4055",x"36da",x"3b14",x"b774",x"0000",x"3a8b",x"3b77",x"375f",x"4055",x"3710",x"3bc1",x"b3d8",x"0000",x"3a96",x"3b77",x"3760",x"4056",x"3710",x"3b92",x"3528",x"8000",x"3a96",x"3b79"),
(x"34bb",x"4042",x"36da",x"b13f",x"bbe4",x"0000",x"3a50",x"3b84",x"34bb",x"4042",x"3710",x"b31c",x"bbcc",x"0000",x"3a5a",x"3b84",x"34cb",x"4041",x"3710",x"b64c",x"bb5a",x"0000",x"3a5a",x"3b87"),
(x"388c",x"4041",x"36da",x"bbfd",x"29ab",x"0000",x"3a72",x"3ac9",x"388c",x"4041",x"3710",x"bb54",x"3669",x"8000",x"3a7c",x"3ac9",x"3885",x"4040",x"3710",x"b7eb",x"3af3",x"0000",x"3a7c",x"3acc"),
(x"380a",x"404d",x"36da",x"ad54",x"3bf8",x"8000",x"3a8b",x"3b4a",x"380a",x"404d",x"3710",x"ae11",x"3bf6",x"0000",x"3a96",x"3b4a",x"37b8",x"404c",x"3710",x"30d0",x"3be8",x"0000",x"3a96",x"3b5c"),
(x"349b",x"4042",x"36da",x"b4a8",x"bba7",x"8000",x"3a50",x"3b7e",x"349b",x"4042",x"3710",x"b221",x"bbda",x"0000",x"3a5a",x"3b7e",x"34bb",x"4042",x"3710",x"b31c",x"bbcc",x"0000",x"3a5a",x"3b84"),
(x"388c",x"4042",x"36da",x"b967",x"b9e6",x"0000",x"3a72",x"3ac8",x"388c",x"4042",x"3710",x"bb52",x"b671",x"0000",x"3a7c",x"3ac8",x"388c",x"4041",x"3710",x"bb54",x"3669",x"8000",x"3a7c",x"3ac9"),
(x"37b8",x"404c",x"36da",x"2df3",x"3bf7",x"0000",x"3a8b",x"3b5c",x"37b8",x"404c",x"3710",x"30d0",x"3be8",x"0000",x"3a96",x"3b5c",x"37a8",x"404c",x"3710",x"3580",x"3b83",x"0000",x"3a96",x"3b5f"),
(x"3485",x"4043",x"36da",x"b92c",x"ba1a",x"8000",x"3a50",x"3b7a",x"3485",x"4043",x"3710",x"b819",x"bade",x"0000",x"3a5a",x"3b7a",x"349b",x"4042",x"3710",x"b221",x"bbda",x"0000",x"3a5a",x"3b7e"),
(x"3885",x"4042",x"36da",x"b25f",x"bbd7",x"0000",x"3a42",x"3bad",x"3885",x"4042",x"3710",x"b304",x"bbce",x"0000",x"3a4c",x"3bad",x"388c",x"4042",x"3710",x"bb52",x"b671",x"0000",x"3a4c",x"3bb0"),
(x"37a8",x"404c",x"36da",x"33d5",x"3bc1",x"0000",x"3a8b",x"3b5f",x"37a8",x"404c",x"3710",x"3580",x"3b83",x"0000",x"3a96",x"3b5f",x"378c",x"404e",x"3710",x"3688",x"3b4d",x"8000",x"3a96",x"3b65"),
(x"3a2f",x"404d",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"3816",x"3a2f",x"404d",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"381d",x"3a26",x"404d",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3820"),
(x"3475",x"4045",x"36da",x"bbab",x"b48e",x"0000",x"3a50",x"3b75",x"3475",x"4045",x"3710",x"baeb",x"b803",x"0000",x"3a5a",x"3b75",x"3485",x"4043",x"3710",x"b819",x"bade",x"0000",x"3a5a",x"3b7a"),
(x"3753",x"4037",x"36da",x"37e4",x"baf5",x"8000",x"3a42",x"3b48",x"3753",x"4037",x"3710",x"38fe",x"ba3f",x"0000",x"3a4c",x"3b48",x"3760",x"4038",x"3710",x"3bfa",x"acac",x"868d",x"3a4c",x"3b4c"),
(x"378c",x"404e",x"36da",x"373a",x"3b23",x"0000",x"3a8b",x"3b65",x"378c",x"404e",x"3710",x"3688",x"3b4d",x"8000",x"3a96",x"3b65",x"376c",x"4050",x"3710",x"3899",x"3a8b",x"0000",x"3a96",x"3b6c"),
(x"382a",x"4042",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b89",x"382a",x"4042",x"3710",x"2f40",x"bbf2",x"0000",x"3a4c",x"3b89",x"3885",x"4042",x"3710",x"b304",x"bbce",x"0000",x"3a4c",x"3bad"),
(x"376c",x"4050",x"36da",x"3787",x"3b0e",x"0000",x"3a8b",x"3b6c",x"376c",x"4050",x"3710",x"3899",x"3a8b",x"0000",x"3a96",x"3b6c",x"3752",x"4053",x"3710",x"3bfd",x"aac2",x"0000",x"3a96",x"3b72"),
(x"3999",x"4037",x"36da",x"b32b",x"bbcb",x"0000",x"39fd",x"3b78",x"3999",x"4037",x"3710",x"b2ba",x"bbd2",x"0000",x"3a07",x"3b78",x"39fc",x"4036",x"3710",x"9bc8",x"bc00",x"200b",x"3a07",x"3b9f"),
(x"3813",x"4041",x"36da",x"a8bf",x"bbfe",x"8000",x"3a42",x"3b80",x"3813",x"4041",x"3710",x"27fc",x"bbfe",x"0000",x"3a4c",x"3b80",x"382a",x"4042",x"3710",x"2f40",x"bbf2",x"0000",x"3a4c",x"3b89"),
(x"3753",x"4058",x"36da",x"38fe",x"3a3f",x"8000",x"3a8b",x"3b7d",x"3753",x"4058",x"3710",x"37e4",x"3af5",x"8000",x"3a96",x"3b7d",x"3742",x"4059",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b80"),
(x"380a",x"4041",x"36da",x"ae12",x"bbf6",x"0000",x"3a42",x"3b7c",x"380a",x"4041",x"3710",x"ad56",x"bbf8",x"0000",x"3a4c",x"3b7c",x"3813",x"4041",x"3710",x"27fc",x"bbfe",x"0000",x"3a4c",x"3b80"),
(x"3742",x"4059",x"36da",x"342c",x"3bb9",x"8000",x"3a8b",x"3b80",x"3742",x"4059",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b80",x"372e",x"4059",x"3710",x"338a",x"3bc6",x"0000",x"3a96",x"3b84"),
(x"3760",x"4038",x"36da",x"3b92",x"b528",x"0000",x"3a42",x"3b4c",x"3760",x"4038",x"3710",x"3bfa",x"acac",x"868d",x"3a4c",x"3b4c",x"375f",x"403a",x"3710",x"3b14",x"3774",x"8000",x"3a4c",x"3b4e"),
(x"372e",x"4059",x"36da",x"2fc6",x"3bf0",x"0000",x"3a8b",x"3b84",x"372e",x"4059",x"3710",x"338a",x"3bc6",x"0000",x"3a96",x"3b84",x"3716",x"405a",x"3710",x"32c2",x"3bd1",x"8000",x"3a96",x"3b89"),
(x"37b8",x"4043",x"36da",x"30d0",x"bbe8",x"0000",x"3a42",x"3b6a",x"37b8",x"4043",x"3710",x"2df5",x"bbf7",x"0000",x"3a4c",x"3b6a",x"380a",x"4041",x"3710",x"ad56",x"bbf8",x"0000",x"3a4c",x"3b7c"),
(x"3716",x"405a",x"36da",x"34b5",x"3ba5",x"8000",x"3a8b",x"3b89",x"3716",x"405a",x"3710",x"32c2",x"3bd1",x"8000",x"3a96",x"3b89",x"36f7",x"405b",x"3710",x"b463",x"3bb1",x"8000",x"3a96",x"3b8f"),
(x"37a8",x"4043",x"36da",x"3580",x"bb83",x"0000",x"3a42",x"3b66",x"37a8",x"4043",x"3710",x"33d5",x"bbc1",x"0000",x"3a4c",x"3b66",x"37b8",x"4043",x"3710",x"2df5",x"bbf7",x"0000",x"3a4c",x"3b6a"),
(x"36f7",x"405b",x"36da",x"ae6b",x"3bf5",x"0000",x"3a8b",x"3b8f",x"36f7",x"405b",x"3710",x"b463",x"3bb1",x"8000",x"3a96",x"3b8f",x"36e3",x"405a",x"3710",x"bb17",x"3766",x"868d",x"3a96",x"3b93"),
(x"378c",x"4041",x"36da",x"3688",x"bb4d",x"8000",x"3a42",x"3b60",x"378c",x"4041",x"3710",x"373a",x"bb23",x"0000",x"3a4c",x"3b60",x"37a8",x"4043",x"3710",x"33d5",x"bbc1",x"0000",x"3a4c",x"3b66"),
(x"36e3",x"405a",x"36da",x"b9b5",x"399a",x"0000",x"3a8b",x"3b93",x"36e3",x"405a",x"3710",x"bb17",x"3766",x"868d",x"3a96",x"3b93",x"36df",x"4058",x"3710",x"bbc6",x"338f",x"8000",x"3a96",x"3b96"),
(x"376c",x"403f",x"36da",x"3899",x"ba8b",x"0000",x"3a42",x"3b59",x"376c",x"403f",x"3710",x"3787",x"bb0e",x"0000",x"3a4c",x"3b59",x"378c",x"4041",x"3710",x"373a",x"bb23",x"0000",x"3a4c",x"3b60"),
(x"36df",x"4058",x"36da",x"bbbc",x"3412",x"0000",x"3a8b",x"3b96",x"36df",x"4058",x"3710",x"bbc6",x"338f",x"8000",x"3a96",x"3b96",x"36dc",x"4056",x"3710",x"bb3a",x"36da",x"0000",x"3a96",x"3b98"),
(x"3a26",x"404d",x"36da",x"3bff",x"a4d0",x"0000",x"39d6",x"33f3",x"3a26",x"404d",x"3710",x"3bed",x"a7ae",x"3024",x"39d7",x"33c4",x"3a27",x"4059",x"3710",x"3bea",x"a4d6",x"30a2",x"39ea",x"33c9"),
(x"39f5",x"4059",x"36da",x"a49b",x"3bff",x"8000",x"3a2d",x"3b9f",x"39f5",x"4059",x"3710",x"a4e3",x"3bff",x"1818",x"3a23",x"3b9f",x"3999",x"4058",x"3710",x"b329",x"3bcb",x"8000",x"3a23",x"3b7b"),
(x"3752",x"403c",x"36da",x"3bfd",x"2ac2",x"0000",x"3a42",x"3b53",x"3752",x"403c",x"3710",x"3be0",x"b1a3",x"068d",x"3a4c",x"3b53",x"376c",x"403f",x"3710",x"3787",x"bb0e",x"0000",x"3a4c",x"3b59"),
(x"36dc",x"4056",x"36da",x"bba4",x"34ba",x"0000",x"3a8b",x"3b98",x"36dc",x"4056",x"3710",x"bb3a",x"36da",x"0000",x"3a96",x"3b98",x"36c4",x"4053",x"3710",x"bbc5",x"339b",x"068d",x"3a96",x"3b9f"),
(x"3999",x"4058",x"36da",x"b2b0",x"3bd2",x"0000",x"3a2d",x"3b7b",x"3999",x"4058",x"3710",x"b329",x"3bcb",x"8000",x"3a23",x"3b7b",x"3994",x"4058",x"3710",x"b59f",x"3b7d",x"0000",x"3a23",x"3b79"),
(x"3742",x"4036",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b44",x"3742",x"4036",x"3710",x"342c",x"bbb9",x"0000",x"3a4c",x"3b44",x"3753",x"4037",x"3710",x"38fe",x"ba3f",x"0000",x"3a4c",x"3b48"),
(x"36c4",x"4053",x"36da",x"bb61",x"362a",x"0000",x"3a8b",x"3b9f",x"36c4",x"4053",x"3710",x"bbc5",x"339b",x"068d",x"3a96",x"3b9f",x"36c2",x"4051",x"3710",x"bafe",x"b7c2",x"0000",x"3a96",x"3ba1"),
(x"3994",x"4058",x"36da",x"b458",x"3bb2",x"8000",x"3a2d",x"3b79",x"3994",x"4058",x"3710",x"b59f",x"3b7d",x"0000",x"3a23",x"3b79",x"3985",x"4055",x"3710",x"b796",x"3b0b",x"0000",x"3a23",x"3b72"),
(x"372e",x"4036",x"36da",x"338a",x"bbc6",x"0000",x"3a42",x"3b40",x"372e",x"4036",x"3710",x"2fc6",x"bbf0",x"0000",x"3a4c",x"3b40",x"3742",x"4036",x"3710",x"342c",x"bbb9",x"0000",x"3a4c",x"3b44"),
(x"36c2",x"4051",x"36da",x"bbe7",x"b0ec",x"0000",x"3a8b",x"3ba1",x"36c2",x"4051",x"3710",x"bafe",x"b7c2",x"0000",x"3a96",x"3ba1",x"36cb",x"4050",x"3710",x"b86c",x"baa9",x"0000",x"3a96",x"3ba3"),
(x"3985",x"4055",x"36da",x"b817",x"3adf",x"0000",x"3a2d",x"3b72",x"3985",x"4055",x"3710",x"b796",x"3b0b",x"0000",x"3a23",x"3b72",x"3972",x"4053",x"3710",x"b0a0",x"3bea",x"0000",x"3a23",x"3b6a"),
(x"3716",x"4035",x"36da",x"32c2",x"bbd1",x"0000",x"3a42",x"3b3b",x"3716",x"4035",x"3710",x"34b5",x"bba5",x"0000",x"3a4c",x"3b3b",x"372e",x"4036",x"3710",x"2fc6",x"bbf0",x"0000",x"3a4c",x"3b40"),
(x"36cb",x"4050",x"36da",x"b922",x"ba22",x"068d",x"3a8b",x"3ba3",x"36cb",x"4050",x"3710",x"b86c",x"baa9",x"0000",x"3a96",x"3ba3",x"3705",x"404f",x"3710",x"b675",x"bb51",x"0000",x"3a96",x"3bae"),
(x"3972",x"4053",x"36da",x"b475",x"3bae",x"0000",x"3a2d",x"3b6a",x"3972",x"4053",x"3710",x"b0a0",x"3bea",x"0000",x"3a23",x"3b6a",x"3963",x"4053",x"3710",x"36c5",x"3b3f",x"0000",x"3a23",x"3b64"),
(x"36f7",x"4034",x"36da",x"b463",x"bbb1",x"8000",x"3a42",x"3b35",x"36f7",x"4034",x"3710",x"ae6b",x"bbf5",x"0000",x"3a4c",x"3b35",x"3716",x"4035",x"3710",x"34b5",x"bba5",x"0000",x"3a4c",x"3b3b"),
(x"3705",x"404f",x"36da",x"b599",x"bb7e",x"0000",x"3a8b",x"3bae",x"3705",x"404f",x"3710",x"b675",x"bb51",x"0000",x"3a96",x"3bae",x"3713",x"404e",x"3710",x"ba37",x"b909",x"0000",x"3a96",x"3bb1"),
(x"3963",x"4053",x"36da",x"3420",x"3bba",x"0000",x"3a2d",x"3b64",x"3963",x"4053",x"3710",x"36c5",x"3b3f",x"0000",x"3a23",x"3b64",x"395d",x"4054",x"3710",x"3ac1",x"3849",x"0000",x"3a23",x"3b61"),
(x"36e3",x"4035",x"36da",x"bb17",x"b766",x"068d",x"3a42",x"3b31",x"36e3",x"4035",x"3710",x"b9b5",x"b99a",x"0000",x"3a4c",x"3b31",x"36f7",x"4034",x"3710",x"ae6b",x"bbf5",x"0000",x"3a4c",x"3b35"),
(x"3713",x"404e",x"36da",x"b972",x"b9db",x"8000",x"3a8b",x"3bb1",x"3713",x"404e",x"3710",x"ba37",x"b909",x"0000",x"3a96",x"3bb1",x"3716",x"404e",x"3710",x"bbad",x"3480",x"0000",x"3a96",x"3bb2"),
(x"395d",x"4054",x"36da",x"399d",x"39b2",x"0000",x"3a2d",x"3b61",x"395d",x"4054",x"3710",x"3ac1",x"3849",x"0000",x"3a23",x"3b61",x"395a",x"4055",x"3710",x"3af1",x"37f3",x"0000",x"3a23",x"3b5e"),
(x"36df",x"4037",x"36da",x"bbc6",x"b38f",x"8000",x"3a42",x"3b2e",x"36df",x"4037",x"3710",x"bbbc",x"b412",x"0000",x"3a4c",x"3b2e",x"36e3",x"4035",x"3710",x"b9b5",x"b99a",x"0000",x"3a4c",x"3b31"),
(x"3716",x"404e",x"36da",x"bbb8",x"b42d",x"0000",x"3b11",x"39ae",x"3716",x"404e",x"3710",x"bbad",x"3480",x"0000",x"3b1c",x"39ae",x"3710",x"404d",x"3710",x"b80d",x"3ae5",x"0000",x"3b1c",x"39af"),
(x"395a",x"4055",x"36da",x"3b46",x"36a7",x"8000",x"3a2d",x"3b5e",x"395a",x"4055",x"3710",x"3af1",x"37f3",x"0000",x"3a23",x"3b5e",x"3953",x"4058",x"3710",x"3857",x"3ab8",x"8000",x"3a23",x"3b5a"),
(x"36dc",x"4038",x"36da",x"bb3a",x"b6d9",x"0000",x"3a42",x"3b2b",x"36dc",x"4038",x"3710",x"bba4",x"b4ba",x"0000",x"3a4c",x"3b2b",x"36df",x"4037",x"3710",x"bbbc",x"b412",x"0000",x"3a4c",x"3b2e"),
(x"3710",x"404d",x"36da",x"b8f7",x"3a45",x"0000",x"3b11",x"39af",x"3710",x"404d",x"3710",x"b80d",x"3ae5",x"0000",x"3b1c",x"39af",x"36f7",x"404c",x"3710",x"b05b",x"3bec",x"8000",x"3b1c",x"39b4"),
(x"3475",x"404a",x"36da",x"baeb",x"3803",x"8000",x"3a50",x"3b6f",x"3475",x"404a",x"3710",x"bbab",x"348e",x"8000",x"3a5a",x"3b6f",x"3475",x"4045",x"3710",x"baeb",x"b803",x"0000",x"3a5a",x"3b75"),
(x"3953",x"4058",x"36da",x"39a8",x"39a7",x"868d",x"3a2d",x"3b5a",x"3953",x"4058",x"3710",x"3857",x"3ab8",x"8000",x"3a23",x"3b5a",x"393f",x"4059",x"3710",x"b2bb",x"3bd2",x"868d",x"3a23",x"3b51"),
(x"36c4",x"403c",x"36da",x"bbc5",x"b39b",x"0000",x"3a42",x"3b24",x"36c4",x"403c",x"3710",x"bb61",x"b62a",x"0000",x"3a4c",x"3b24",x"36dc",x"4038",x"3710",x"bba4",x"b4ba",x"0000",x"3a4c",x"3b2b"),
(x"363b",x"404c",x"36da",x"3439",x"3bb7",x"0000",x"3b11",x"39d8",x"363b",x"404c",x"3710",x"34bd",x"3ba4",x"0000",x"3b1c",x"39d8",x"362c",x"404d",x"3710",x"3609",x"3b68",x"8000",x"3b1c",x"39db"),
(x"3994",x"4037",x"36da",x"b59f",x"bb7d",x"0000",x"39fd",x"3b76",x"3994",x"4037",x"3710",x"b459",x"bbb2",x"068d",x"3a07",x"3b76",x"3999",x"4037",x"3710",x"b2ba",x"bbd2",x"0000",x"3a07",x"3b78"),
(x"393f",x"4059",x"36da",x"1cea",x"3c00",x"0000",x"3a2d",x"3b51",x"393f",x"4059",x"3710",x"b2bb",x"3bd2",x"868d",x"3a23",x"3b51",x"392f",x"4057",x"3710",x"b874",x"3aa4",x"0000",x"3a23",x"3b4b"),
(x"36c2",x"403d",x"36da",x"bafe",x"37c2",x"8000",x"3a42",x"3b22",x"36c2",x"403d",x"3710",x"bbe7",x"30ec",x"868d",x"3a4c",x"3b22",x"36c4",x"403c",x"3710",x"bb61",x"b62a",x"0000",x"3a4c",x"3b24"),
(x"36f7",x"404c",x"36da",x"b12d",x"3be4",x"0000",x"3b11",x"39b4",x"36f7",x"404c",x"3710",x"b05b",x"3bec",x"8000",x"3b1c",x"39b4",x"363b",x"404c",x"3710",x"34bd",x"3ba4",x"0000",x"3b1c",x"39d8"),
(x"3985",x"403a",x"36da",x"b796",x"bb0b",x"0000",x"39fd",x"3b6f",x"3985",x"403a",x"3710",x"b817",x"badf",x"0000",x"3a07",x"3b6f",x"3994",x"4037",x"3710",x"b459",x"bbb2",x"068d",x"3a07",x"3b76"),
(x"3752",x"4053",x"36da",x"3be0",x"31a3",x"8000",x"3a8b",x"3b72",x"3752",x"4053",x"3710",x"3bfd",x"aac2",x"0000",x"3a96",x"3b72",x"3754",x"4054",x"3710",x"3afe",x"b7c4",x"0000",x"3a96",x"3b74"),
(x"36cb",x"403e",x"36da",x"b86c",x"3aaa",x"0000",x"3a42",x"3b1f",x"36cb",x"403e",x"3710",x"b922",x"3a22",x"0000",x"3a4c",x"3b1f",x"36c2",x"403d",x"3710",x"bbe7",x"30ec",x"868d",x"3a4c",x"3b22"),
(x"362c",x"404d",x"36da",x"3550",x"3b8b",x"0000",x"3b11",x"39db",x"362c",x"404d",x"3710",x"3609",x"3b68",x"8000",x"3b1c",x"39db",x"35f7",x"4051",x"3710",x"3a6a",x"38c7",x"0000",x"3b1c",x"39e6"),
(x"3972",x"403c",x"36da",x"b0a0",x"bbea",x"0000",x"39fd",x"3b67",x"3972",x"403c",x"3710",x"b475",x"bbae",x"0000",x"3a07",x"3b67",x"3985",x"403a",x"3710",x"b817",x"badf",x"0000",x"3a07",x"3b6f"),
(x"392f",x"4057",x"36da",x"b73b",x"3b22",x"8000",x"3a2d",x"3b4b",x"392f",x"4057",x"3710",x"b874",x"3aa4",x"0000",x"3a23",x"3b4b",x"3915",x"4051",x"3710",x"b845",x"3ac3",x"0000",x"3a23",x"3b3c"),
(x"3705",x"4040",x"36da",x"b675",x"3b51",x"0000",x"3a42",x"3b14",x"3705",x"4040",x"3710",x"b599",x"3b7e",x"0000",x"3a4c",x"3b14",x"36cb",x"403e",x"3710",x"b922",x"3a22",x"0000",x"3a4c",x"3b1f"),
(x"35f7",x"4051",x"36da",x"3a05",x"3944",x"868d",x"3b11",x"39e6",x"35f7",x"4051",x"3710",x"3a6a",x"38c7",x"0000",x"3b1c",x"39e6",x"35f1",x"4052",x"3710",x"3bf9",x"ad20",x"0000",x"3b1c",x"39e8"),
(x"3963",x"403c",x"36da",x"36c5",x"bb3f",x"0000",x"39fd",x"3b61",x"3963",x"403c",x"3710",x"3420",x"bbba",x"0000",x"3a07",x"3b61",x"3972",x"403c",x"3710",x"b475",x"bbae",x"0000",x"3a07",x"3b67"),
(x"3754",x"4054",x"36da",x"3ba5",x"b4b5",x"0000",x"3a8b",x"3b74",x"3754",x"4054",x"3710",x"3afe",x"b7c4",x"0000",x"3a96",x"3b74",x"375f",x"4055",x"3710",x"3bc1",x"b3d8",x"0000",x"3a96",x"3b77"),
(x"3713",x"4041",x"36da",x"ba37",x"3909",x"0000",x"3a42",x"3b11",x"3713",x"4041",x"3710",x"b972",x"39db",x"0000",x"3a4c",x"3b11",x"3705",x"4040",x"3710",x"b599",x"3b7e",x"0000",x"3a4c",x"3b14"),
(x"35f1",x"4052",x"36da",x"3bcd",x"3318",x"0000",x"3b11",x"39e8",x"35f1",x"4052",x"3710",x"3bf9",x"ad20",x"0000",x"3b1c",x"39e8",x"35f3",x"4053",x"3710",x"3b36",x"b6ea",x"8000",x"3b1c",x"39e9"),
(x"395d",x"403b",x"36da",x"3ac1",x"b849",x"0000",x"39fd",x"3b5e",x"395d",x"403b",x"3710",x"399d",x"b9b2",x"0000",x"3a07",x"3b5e",x"3963",x"403c",x"3710",x"3420",x"bbba",x"0000",x"3a07",x"3b61"),
(x"3915",x"4051",x"36da",x"b90a",x"3a36",x"0000",x"3a2d",x"3b3c",x"3915",x"4051",x"3710",x"b845",x"3ac3",x"0000",x"3a23",x"3b3c",x"38f6",x"404d",x"3710",x"b324",x"3bcc",x"0000",x"3a23",x"3b2e"),
(x"3716",x"4041",x"36da",x"bbad",x"b480",x"0000",x"3a42",x"3b10",x"3716",x"4041",x"3710",x"bbb8",x"342d",x"0000",x"3a4c",x"3b10",x"3713",x"4041",x"3710",x"b972",x"39db",x"0000",x"3a4c",x"3b11"),
(x"35f3",x"4053",x"36da",x"3b84",x"b57a",x"0000",x"3b11",x"39e9",x"35f3",x"4053",x"3710",x"3b36",x"b6ea",x"8000",x"3b1c",x"39e9",x"35fd",x"4054",x"3710",x"3bf0",x"aff4",x"868d",x"3b1c",x"39ed"),
(x"395a",x"4039",x"36da",x"3af1",x"b7f3",x"0000",x"39fd",x"3b5b",x"395a",x"4039",x"3710",x"3b46",x"b6a7",x"8000",x"3a07",x"3b5b",x"395d",x"403b",x"3710",x"399d",x"b9b2",x"0000",x"3a07",x"3b5e"),
(x"38f6",x"404d",x"36da",x"b551",x"3b8b",x"0000",x"3a2d",x"3b2e",x"38f6",x"404d",x"3710",x"b324",x"3bcc",x"0000",x"3a23",x"3b2e",x"38d5",x"404c",x"3710",x"2dde",x"3bf7",x"0000",x"3a23",x"3b21"),
(x"3710",x"4042",x"36da",x"b80d",x"bae5",x"8000",x"3af0",x"3a0f",x"3710",x"4042",x"3710",x"b8f7",x"ba45",x"0000",x"3afb",x"3a0f",x"3716",x"4041",x"3710",x"bbb8",x"342d",x"0000",x"3afb",x"3a11"),
(x"35fd",x"4054",x"36da",x"3b91",x"b530",x"8000",x"3b11",x"39ed",x"35fd",x"4054",x"3710",x"3bf0",x"aff4",x"868d",x"3b1c",x"39ed",x"35fd",x"4055",x"3710",x"3a08",x"3941",x"0000",x"3b1c",x"39ee"),
(x"3953",x"4037",x"36da",x"3857",x"bab8",x"8000",x"39fd",x"3b57",x"3953",x"4037",x"3710",x"39a8",x"b9a7",x"0000",x"3a07",x"3b57",x"395a",x"4039",x"3710",x"3b46",x"b6a7",x"8000",x"3a07",x"3b5b"),
(x"38d5",x"404c",x"36da",x"1987",x"3c00",x"0000",x"3a2d",x"3b21",x"38d5",x"404c",x"3710",x"2dde",x"3bf7",x"0000",x"3a23",x"3b21",x"38bf",x"404d",x"3710",x"35f3",x"3b6c",x"0000",x"3a23",x"3b18"),
(x"36f7",x"4042",x"36da",x"b05b",x"bbec",x"8000",x"3af0",x"3a0a",x"36f7",x"4042",x"3710",x"b12d",x"bbe4",x"0000",x"3afb",x"3a0a",x"3710",x"4042",x"3710",x"b8f7",x"ba45",x"0000",x"3afb",x"3a0f"),
(x"35fd",x"4055",x"36da",x"3b87",x"3567",x"8000",x"3b11",x"39ee",x"35fd",x"4055",x"3710",x"3a08",x"3941",x"0000",x"3b1c",x"39ee",x"35f5",x"4056",x"3710",x"32d5",x"3bd0",x"0000",x"3b1c",x"39f0"),
(x"393f",x"4036",x"36da",x"b2bc",x"bbd2",x"8000",x"39fd",x"3b4e",x"393f",x"4036",x"3710",x"1cea",x"bc00",x"8000",x"3a07",x"3b4e",x"3953",x"4037",x"3710",x"39a8",x"b9a7",x"0000",x"3a07",x"3b57"),
(x"38bf",x"404d",x"36da",x"3489",x"3bac",x"0000",x"3a2d",x"3b18",x"38bf",x"404d",x"3710",x"35f3",x"3b6c",x"0000",x"3a23",x"3b18",x"38b2",x"404e",x"3710",x"3af2",x"37f0",x"0000",x"3a23",x"3b13"),
(x"362c",x"4042",x"36da",x"3609",x"bb68",x"0000",x"3af0",x"39e4",x"362c",x"4042",x"3710",x"3550",x"bb8b",x"0000",x"3afb",x"39e4",x"363b",x"4042",x"3710",x"3439",x"bbb7",x"8000",x"3afb",x"39e7"),
(x"35f5",x"4056",x"36da",x"364c",x"3b5a",x"868d",x"3b11",x"39f0",x"35f5",x"4056",x"3710",x"32d5",x"3bd0",x"0000",x"3b1c",x"39f0",x"35e4",x"4056",x"3710",x"b3c3",x"3bc2",x"0000",x"3b1c",x"39f3"),
(x"392f",x"4037",x"36da",x"b874",x"baa4",x"0000",x"39fd",x"3b48",x"392f",x"4037",x"3710",x"b73b",x"bb22",x"0000",x"3a07",x"3b48",x"393f",x"4036",x"3710",x"1cea",x"bc00",x"8000",x"3a07",x"3b4e"),
(x"38b2",x"404e",x"36da",x"3a0a",x"393e",x"8000",x"3a2d",x"3b13",x"38b2",x"404e",x"3710",x"3af2",x"37f0",x"0000",x"3a23",x"3b13",x"38b0",x"4050",x"3710",x"3ba6",x"b4ab",x"0000",x"3a23",x"3b10"),
(x"363b",x"4042",x"36da",x"34be",x"bba4",x"0000",x"3af0",x"39e7",x"363b",x"4042",x"3710",x"3439",x"bbb7",x"8000",x"3afb",x"39e7",x"36f7",x"4042",x"3710",x"b12d",x"bbe4",x"0000",x"3afb",x"3a0a"),
(x"35e4",x"4056",x"36da",x"b0fa",x"3be7",x"8000",x"3b11",x"39f3",x"35e4",x"4056",x"3710",x"b3c3",x"3bc2",x"0000",x"3b1c",x"39f3",x"35d3",x"4055",x"3710",x"1c81",x"3c00",x"0000",x"3b1c",x"39f7"),
(x"3754",x"403b",x"36da",x"3afe",x"37c4",x"0000",x"3a42",x"3b51",x"3754",x"403b",x"3710",x"3ba5",x"34b5",x"0000",x"3a4c",x"3b51",x"3752",x"403c",x"3710",x"3be0",x"b1a3",x"068d",x"3a4c",x"3b53"),
(x"38b0",x"4050",x"36da",x"3bfc",x"2b27",x"0000",x"3a2d",x"3b10",x"38b0",x"4050",x"3710",x"3ba6",x"b4ab",x"0000",x"3a23",x"3b10",x"38b2",x"4051",x"3710",x"399c",x"b9b3",x"0000",x"3a23",x"3b0f"),
(x"35f7",x"403e",x"36da",x"3a6a",x"b8c7",x"0000",x"3af0",x"39d8",x"35f7",x"403e",x"3710",x"3a05",x"b944",x"0000",x"3afb",x"39d8",x"362c",x"4042",x"3710",x"3550",x"bb8b",x"0000",x"3afb",x"39e4"),
(x"35d3",x"4055",x"36da",x"b1d2",x"3bdd",x"0000",x"3b11",x"39f7",x"35d3",x"4055",x"3710",x"1c81",x"3c00",x"0000",x"3b1c",x"39f7",x"35bd",x"4056",x"3710",x"afcb",x"3bf0",x"8000",x"3b1c",x"39fb"),
(x"3915",x"403e",x"36da",x"b845",x"bac3",x"0000",x"39fd",x"3b39",x"3915",x"403e",x"3710",x"b90a",x"ba36",x"0000",x"3a07",x"3b39",x"392f",x"4037",x"3710",x"b73b",x"bb22",x"0000",x"3a07",x"3b48"),
(x"38b2",x"4051",x"36da",x"3a58",x"b8de",x"0000",x"3a88",x"3ac5",x"38b2",x"4051",x"3710",x"399c",x"b9b3",x"0000",x"3a93",x"3ac5",x"38bd",x"4052",x"3710",x"3456",x"bbb3",x"0000",x"3a93",x"3ac9"),
(x"35f1",x"403d",x"36da",x"3bf9",x"2d20",x"0000",x"3af0",x"39d6",x"35f1",x"403d",x"3710",x"3bcd",x"b318",x"0000",x"3afb",x"39d6",x"35f7",x"403e",x"3710",x"3a05",x"b944",x"0000",x"3afb",x"39d8"),
(x"35bd",x"4056",x"36da",x"2c75",x"3bfb",x"068d",x"3b11",x"39fb",x"35bd",x"4056",x"3710",x"afcb",x"3bf0",x"8000",x"3b1c",x"39fb",x"359e",x"4054",x"3710",x"b925",x"3a1f",x"0000",x"3b1c",x"3a01"),
(x"375f",x"403a",x"36da",x"3bc1",x"33d8",x"868d",x"3a42",x"3b4e",x"375f",x"403a",x"3710",x"3b14",x"3774",x"8000",x"3a4c",x"3b4e",x"3754",x"403b",x"3710",x"3ba5",x"34b5",x"0000",x"3a4c",x"3b51"),
(x"38bd",x"4052",x"36da",x"35fc",x"bb6b",x"0000",x"3a88",x"3ac9",x"38bd",x"4052",x"3710",x"3456",x"bbb3",x"0000",x"3a93",x"3ac9",x"38c9",x"4053",x"3710",x"34cb",x"bba1",x"0000",x"3a93",x"3ace"),
(x"35f3",x"403c",x"36da",x"3b36",x"36ea",x"8000",x"3af0",x"39d5",x"35f3",x"403c",x"3710",x"3b84",x"3579",x"0000",x"3afb",x"39d5",x"35f1",x"403d",x"3710",x"3bcd",x"b318",x"0000",x"3afb",x"39d6"),
(x"359e",x"4054",x"36da",x"b80b",x"3ae7",x"8000",x"3b11",x"3a01",x"359e",x"4054",x"3710",x"b925",x"3a1f",x"0000",x"3b1c",x"3a01",x"358a",x"4051",x"3710",x"bbad",x"3481",x"0000",x"3b1c",x"3a07"),
(x"38f6",x"4042",x"36da",x"b324",x"bbcc",x"0000",x"39fd",x"3b2b",x"38f6",x"4042",x"3710",x"b551",x"bb8b",x"0000",x"3a07",x"3b2b",x"3915",x"403e",x"3710",x"b90a",x"ba36",x"0000",x"3a07",x"3b39"),
(x"38c9",x"4053",x"36da",x"3385",x"bbc6",x"0000",x"3a88",x"3ace",x"38c9",x"4053",x"3710",x"34cb",x"bba1",x"0000",x"3a93",x"3ace",x"38d4",x"4054",x"3710",x"38a8",x"ba80",x"8000",x"3a93",x"3ad2"),
(x"35fd",x"403a",x"36da",x"3bf0",x"2ff4",x"868d",x"3af0",x"39d2",x"35fd",x"403a",x"3710",x"3b91",x"3530",x"0000",x"3afb",x"39d2",x"35f3",x"403c",x"3710",x"3b84",x"3579",x"0000",x"3afb",x"39d5"),
(x"358a",x"4051",x"36da",x"bb1e",x"374c",x"8000",x"3b11",x"3a07",x"358a",x"4051",x"3710",x"bbad",x"3481",x"0000",x"3b1c",x"3a07",x"3587",x"404f",x"3710",x"bb8b",x"b553",x"868d",x"3b1c",x"3a0b"),
(x"38d5",x"4043",x"36da",x"2dde",x"bbf7",x"0000",x"39fd",x"3b1e",x"38d5",x"4043",x"3710",x"1987",x"bc00",x"0000",x"3a07",x"3b1e",x"38f6",x"4042",x"3710",x"b551",x"bb8b",x"0000",x"3a07",x"3b2b"),
(x"38d4",x"4054",x"36da",x"37f2",x"baf1",x"8000",x"3a88",x"3ad2",x"38d4",x"4054",x"3710",x"38a8",x"ba80",x"8000",x"3a93",x"3ad2",x"38d9",x"4055",x"3710",x"3bfc",x"ab03",x"8a8d",x"3a93",x"3ad5"),
(x"3a26",x"4036",x"36da",x"3bff",x"26b5",x"0000",x"39b3",x"33fa",x"3a26",x"4036",x"3710",x"3bcf",x"2680",x"32dc",x"39b2",x"33ca",x"3a25",x"4041",x"3710",x"3bd6",x"2604",x"3256",x"39c5",x"33c0"),
(x"35fd",x"4039",x"36da",x"3a08",x"b941",x"8000",x"3af0",x"39d0",x"35fd",x"4039",x"3710",x"3b87",x"b567",x"868d",x"3afb",x"39d0",x"35fd",x"403a",x"3710",x"3b91",x"3530",x"0000",x"3afb",x"39d2"),
(x"3587",x"404f",x"36da",x"bbf7",x"adba",x"8000",x"3b11",x"3a0b",x"3587",x"404f",x"3710",x"bb8b",x"b553",x"868d",x"3b1c",x"3a0b",x"3593",x"404d",x"3710",x"bc00",x"15bc",x"0000",x"3b1c",x"3a0f"),
(x"38bf",x"4042",x"36da",x"35f3",x"bb6c",x"0000",x"39fd",x"3b15",x"38bf",x"4042",x"3710",x"3489",x"bbab",x"0000",x"3a07",x"3b15",x"38d5",x"4043",x"3710",x"1987",x"bc00",x"0000",x"3a07",x"3b1e"),
(x"38d9",x"4055",x"36da",x"3b88",x"b564",x"0000",x"3a88",x"3ad5",x"38d9",x"4055",x"3710",x"3bfc",x"ab03",x"8a8d",x"3a93",x"3ad5",x"38d8",x"4055",x"3710",x"3b96",x"350f",x"0000",x"3a93",x"3ad6"),
(x"35f5",x"4039",x"36da",x"32d5",x"bbd0",x"0000",x"3af0",x"39ce",x"35f5",x"4039",x"3710",x"364b",x"bb5a",x"0000",x"3afb",x"39ce",x"35fd",x"4039",x"3710",x"3b87",x"b567",x"868d",x"3afb",x"39d0"),
(x"3593",x"404d",x"36da",x"bbda",x"b21b",x"0000",x"3b11",x"3a0f",x"3593",x"404d",x"3710",x"bc00",x"15bc",x"0000",x"3b1c",x"3a0f",x"3592",x"404c",x"3710",x"ba08",x"3941",x"0000",x"3b1c",x"3a11"),
(x"38b2",x"4040",x"36da",x"3af2",x"b7f0",x"0000",x"39fd",x"3b10",x"38b2",x"4040",x"3710",x"3a0a",x"b93e",x"0000",x"3a07",x"3b10",x"38bf",x"4042",x"3710",x"3489",x"bbab",x"0000",x"3a07",x"3b15"),
(x"38d8",x"4055",x"36da",x"3be4",x"312f",x"8000",x"3a88",x"3ad6",x"38d8",x"4055",x"3710",x"3b96",x"350f",x"0000",x"3a93",x"3ad6",x"38c7",x"4057",x"3710",x"364a",x"3b5b",x"0000",x"3a93",x"3add"),
(x"35e4",x"4039",x"36da",x"b3c3",x"bbc2",x"0000",x"3af0",x"39cb",x"35e4",x"4039",x"3710",x"b0fa",x"bbe7",x"8000",x"3afb",x"39cb",x"35f5",x"4039",x"3710",x"364b",x"bb5a",x"0000",x"3afb",x"39ce"),
(x"3592",x"404c",x"36da",x"bba4",x"34bb",x"0000",x"3a50",x"3b34",x"3592",x"404c",x"3710",x"ba08",x"3941",x"0000",x"3a5a",x"3b34",x"357d",x"404b",x"3710",x"26bb",x"3bff",x"0000",x"3a5a",x"3b38"),
(x"38b0",x"403f",x"36da",x"3ba6",x"34ac",x"0000",x"3b18",x"38a2",x"38b0",x"403f",x"3710",x"3bfc",x"ab27",x"0000",x"3b18",x"38ac",x"38b2",x"4040",x"3710",x"3a0a",x"b93e",x"0000",x"3b16",x"38ac"),
(x"38c7",x"4057",x"36da",x"3653",x"3b59",x"0000",x"3a88",x"3add",x"38c7",x"4057",x"3710",x"364a",x"3b5b",x"0000",x"3a93",x"3add",x"38b7",x"4059",x"3710",x"32f7",x"3bce",x"0000",x"3a93",x"3ae4"),
(x"35d3",x"403a",x"36da",x"1c81",x"bc00",x"0000",x"3af0",x"39c8",x"35d3",x"403a",x"3710",x"b1d2",x"bbdd",x"0000",x"3afb",x"39c8",x"35e4",x"4039",x"3710",x"b0fa",x"bbe7",x"8000",x"3afb",x"39cb"),
(x"357d",x"404b",x"36da",x"a8c9",x"3bfe",x"0000",x"3a50",x"3b38",x"357d",x"404b",x"3710",x"26bb",x"3bff",x"0000",x"3a5a",x"3b38",x"3555",x"404c",x"3710",x"35eb",x"3b6e",x"0000",x"3a5a",x"3b3f"),
(x"38b2",x"403e",x"36da",x"399c",x"39b3",x"8000",x"3b1a",x"38a2",x"38b2",x"403e",x"3710",x"3a58",x"38de",x"0000",x"3b1a",x"38ac",x"38b0",x"403f",x"3710",x"3bfc",x"ab27",x"0000",x"3b18",x"38ac"),
(x"38b7",x"4059",x"36da",x"3528",x"3b92",x"068d",x"3a88",x"3ae4",x"38b7",x"4059",x"3710",x"32f7",x"3bce",x"0000",x"3a93",x"3ae4",x"3894",x"4059",x"3710",x"b036",x"3bee",x"0000",x"3a93",x"3af1"),
(x"35bd",x"4039",x"36da",x"afcb",x"bbf0",x"0000",x"3af0",x"39c3",x"35bd",x"4039",x"3710",x"2c74",x"bbfb",x"0000",x"3afb",x"39c3",x"35d3",x"403a",x"3710",x"b1d2",x"bbdd",x"0000",x"3afb",x"39c8"),
(x"3555",x"404c",x"36da",x"345b",x"3bb2",x"0000",x"3a50",x"3b3f",x"3555",x"404c",x"3710",x"35eb",x"3b6e",x"0000",x"3a5a",x"3b3f",x"353f",x"404d",x"3710",x"379f",x"3b08",x"0000",x"3a5a",x"3b44"),
(x"38bd",x"403d",x"36da",x"3456",x"3bb3",x"0000",x"3b1e",x"38a2",x"38bd",x"403d",x"3710",x"35fc",x"3b6b",x"0000",x"3b1e",x"38ac",x"38b2",x"403e",x"3710",x"3a58",x"38de",x"0000",x"3b1a",x"38ac"),
(x"3894",x"4059",x"36da",x"aa0a",x"3bfd",x"8000",x"3a88",x"3af1",x"3894",x"4059",x"3710",x"b036",x"3bee",x"0000",x"3a93",x"3af1",x"3877",x"4058",x"3710",x"b8aa",x"3a7f",x"868d",x"3a93",x"3afc"),
(x"359e",x"403a",x"36da",x"b925",x"ba1f",x"0000",x"3af0",x"39bd",x"359e",x"403a",x"3710",x"b80b",x"bae7",x"0000",x"3afb",x"39bd",x"35bd",x"4039",x"3710",x"2c74",x"bbfb",x"0000",x"3afb",x"39c3"),
(x"353f",x"404d",x"36da",x"3746",x"3b1f",x"0000",x"3a50",x"3b44",x"353f",x"404d",x"3710",x"379f",x"3b08",x"0000",x"3a5a",x"3b44",x"351b",x"4050",x"3710",x"350e",x"3b96",x"0000",x"3a5a",x"3b4c"),
(x"38c9",x"403c",x"36da",x"34cb",x"3ba1",x"8000",x"3a72",x"3b0f",x"38c9",x"403c",x"3710",x"3385",x"3bc6",x"0000",x"3a7c",x"3b0f",x"38bd",x"403d",x"3710",x"35fc",x"3b6b",x"0000",x"3a7c",x"3b13"),
(x"3877",x"4058",x"36da",x"b74e",x"3b1d",x"0000",x"3a88",x"3afc",x"3877",x"4058",x"3710",x"b8aa",x"3a7f",x"868d",x"3a93",x"3afc",x"386d",x"4056",x"3710",x"bba8",x"34a3",x"868d",x"3a93",x"3b01"),
(x"358a",x"403d",x"36da",x"bbad",x"b481",x"068d",x"3af0",x"39b7",x"358a",x"403d",x"3710",x"bb1e",x"b74c",x"0000",x"3afb",x"39b7",x"359e",x"403a",x"3710",x"b80b",x"bae7",x"0000",x"3afb",x"39bd"),
(x"351b",x"4050",x"36da",x"3664",x"3b55",x"0000",x"3a50",x"3b4c",x"351b",x"4050",x"3710",x"350e",x"3b96",x"0000",x"3a5a",x"3b4c",x"3501",x"4051",x"3710",x"ada8",x"3bf8",x"0000",x"3a5a",x"3b51"),
(x"38d4",x"403b",x"36da",x"38a8",x"3a80",x"8000",x"3a72",x"3b0b",x"38d4",x"403b",x"3710",x"37f2",x"3af1",x"8000",x"3a7c",x"3b0b",x"38c9",x"403c",x"3710",x"3385",x"3bc6",x"0000",x"3a7c",x"3b0f"),
(x"386d",x"4056",x"36da",x"bac4",x"3844",x"068d",x"3a88",x"3b01",x"386d",x"4056",x"3710",x"bba8",x"34a3",x"868d",x"3a93",x"3b01",x"386c",x"4053",x"3710",x"bb38",x"b6e2",x"868d",x"3a93",x"3b05"),
(x"3587",x"4040",x"36da",x"bb8b",x"3553",x"0000",x"3af0",x"39b3",x"3587",x"4040",x"3710",x"bbf7",x"2dba",x"868d",x"3afb",x"39b3",x"358a",x"403d",x"3710",x"bb1e",x"b74c",x"0000",x"3afb",x"39b7"),
(x"3501",x"4051",x"36da",x"2d0c",x"3bf9",x"8000",x"3a50",x"3b51",x"3501",x"4051",x"3710",x"ada8",x"3bf8",x"0000",x"3a5a",x"3b51",x"34e9",x"4050",x"3710",x"b698",x"3b49",x"0000",x"3a5a",x"3b56"),
(x"38d9",x"403a",x"36da",x"3bfc",x"2b03",x"0a8d",x"3a72",x"3b08",x"38d9",x"403a",x"3710",x"3b87",x"3565",x"0000",x"3a7c",x"3b08",x"38d4",x"403b",x"3710",x"37f2",x"3af1",x"8000",x"3a7c",x"3b0b"),
(x"386c",x"4053",x"36da",x"bbdd",x"b1e1",x"8000",x"3a88",x"3b05",x"386c",x"4053",x"3710",x"bb38",x"b6e2",x"868d",x"3a93",x"3b05",x"3872",x"4051",x"3710",x"b902",x"ba3c",x"0000",x"3a93",x"3b08"),
(x"3593",x"4042",x"36da",x"bc00",x"95bc",x"0000",x"3af0",x"39af",x"3593",x"4042",x"3710",x"bbda",x"321b",x"8000",x"3afb",x"39af",x"3587",x"4040",x"3710",x"bbf7",x"2dba",x"868d",x"3afb",x"39b3"),
(x"34e9",x"4050",x"36da",x"b50d",x"3b97",x"8000",x"3a50",x"3b56",x"34e9",x"4050",x"3710",x"b698",x"3b49",x"0000",x"3a5a",x"3b56",x"34cb",x"404e",x"3710",x"b501",x"3b99",x"0000",x"3a5a",x"3b5d"),
(x"38d8",x"4039",x"36da",x"3b96",x"b50f",x"0000",x"3a72",x"3b07",x"38d8",x"4039",x"3710",x"3be4",x"b12f",x"868d",x"3a7c",x"3b07",x"38d9",x"403a",x"3710",x"3b87",x"3565",x"0000",x"3a7c",x"3b08"),
(x"3872",x"4051",x"36da",x"b9d1",x"b97d",x"068d",x"3a88",x"3b08",x"3872",x"4051",x"3710",x"b902",x"ba3c",x"0000",x"3a93",x"3b08",x"3885",x"404f",x"3710",x"b83d",x"bac8",x"0000",x"3a93",x"3b10"),
(x"3592",x"4043",x"36da",x"ba08",x"b941",x"8000",x"3af0",x"39ae",x"3592",x"4043",x"3710",x"bba4",x"b4bb",x"0000",x"3afb",x"39ae",x"3593",x"4042",x"3710",x"bbda",x"321b",x"8000",x"3afb",x"39af"),
(x"34cb",x"404e",x"36da",x"b64c",x"3b5a",x"0000",x"3a50",x"3b5d",x"34cb",x"404e",x"3710",x"b501",x"3b99",x"0000",x"3a5a",x"3b5d",x"34bb",x"404d",x"3710",x"b141",x"3be4",x"0000",x"3a5a",x"3b60"),
(x"38c7",x"4038",x"36da",x"364a",x"bb5b",x"8000",x"3a72",x"3b00",x"38c7",x"4038",x"3710",x"3653",x"bb59",x"0000",x"3a7c",x"3b00",x"38d8",x"4039",x"3710",x"3be4",x"b12f",x"868d",x"3a7c",x"3b07"),
(x"3885",x"404f",x"36da",x"b7ea",x"baf3",x"8000",x"3a88",x"3b10",x"3885",x"404f",x"3710",x"b83d",x"bac8",x"0000",x"3a93",x"3b10",x"388c",x"404e",x"3710",x"bbfd",x"a9ab",x"0000",x"3a93",x"3b13"),
(x"357d",x"4043",x"36da",x"26c2",x"bbff",x"0000",x"3a50",x"3bac",x"357d",x"4043",x"3710",x"a8c9",x"bbfe",x"0000",x"3a5a",x"3bac",x"3592",x"4043",x"3710",x"bba4",x"b4bb",x"0000",x"3a5a",x"3bb0"),
(x"34bb",x"404d",x"36da",x"b31c",x"3bcc",x"0000",x"3a50",x"3b60",x"34bb",x"404d",x"3710",x"b141",x"3be4",x"0000",x"3a5a",x"3b60",x"349b",x"404d",x"3710",x"b4a8",x"3ba7",x"0000",x"3a5a",x"3b66"),
(x"38b7",x"4036",x"36da",x"32f6",x"bbce",x"0000",x"3a72",x"3af9",x"38b7",x"4036",x"3710",x"3528",x"bb92",x"0000",x"3a7c",x"3af9",x"38c7",x"4038",x"3710",x"3653",x"bb59",x"0000",x"3a7c",x"3b00"),
(x"388c",x"404e",x"36da",x"bb54",x"b669",x"8000",x"3a8b",x"3b18",x"388c",x"404e",x"3710",x"bbfd",x"a9ab",x"0000",x"3a96",x"3b18",x"388c",x"404d",x"3710",x"b967",x"39e6",x"0000",x"3a96",x"3b19"),
(x"3555",x"4043",x"36da",x"35eb",x"bb6e",x"0000",x"3a50",x"3ba5",x"3555",x"4043",x"3710",x"345a",x"bbb2",x"0000",x"3a5a",x"3ba5",x"357d",x"4043",x"3710",x"a8c9",x"bbfe",x"0000",x"3a5a",x"3bac"),
(x"349b",x"404d",x"36da",x"b221",x"3bda",x"0000",x"3a50",x"3b66",x"349b",x"404d",x"3710",x"b4a8",x"3ba7",x"0000",x"3a5a",x"3b66",x"3485",x"404c",x"3710",x"b92c",x"3a1a",x"0000",x"3a5a",x"3b6a"),
(x"3894",x"4035",x"36da",x"b036",x"bbee",x"0000",x"3a72",x"3aec",x"3894",x"4035",x"3710",x"aa0a",x"bbfd",x"8000",x"3a7c",x"3aec",x"38b7",x"4036",x"3710",x"3528",x"bb92",x"0000",x"3a7c",x"3af9"),
(x"388c",x"404d",x"36da",x"bb52",x"3671",x"0000",x"3a8b",x"3b19",x"388c",x"404d",x"3710",x"b967",x"39e6",x"0000",x"3a96",x"3b19",x"3885",x"404c",x"3710",x"b25f",x"3bd7",x"8000",x"3a96",x"3b1c"),
(x"353f",x"4041",x"36da",x"379f",x"bb08",x"0000",x"3a50",x"3ba0",x"353f",x"4041",x"3710",x"3746",x"bb1f",x"0000",x"3a5a",x"3ba0",x"3555",x"4043",x"3710",x"345a",x"bbb2",x"0000",x"3a5a",x"3ba5"),
(x"3485",x"404c",x"36da",x"b819",x"3ade",x"8000",x"3a50",x"3b6a",x"3485",x"404c",x"3710",x"b92c",x"3a1a",x"0000",x"3a5a",x"3b6a",x"3475",x"404a",x"3710",x"bbab",x"348e",x"8000",x"3a5a",x"3b6f"),
(x"3877",x"4037",x"36da",x"b8aa",x"ba7f",x"868d",x"3a72",x"3ae1",x"3877",x"4037",x"3710",x"b74e",x"bb1d",x"8000",x"3a7c",x"3ae1",x"3894",x"4035",x"3710",x"aa0a",x"bbfd",x"8000",x"3a7c",x"3aec"),
(x"3760",x"4056",x"36da",x"3bfa",x"2cac",x"868d",x"3a8b",x"3b79",x"3760",x"4056",x"3710",x"3b92",x"3528",x"8000",x"3a96",x"3b79",x"3753",x"4058",x"3710",x"37e4",x"3af5",x"8000",x"3a96",x"3b7d"),
(x"3a2d",x"4042",x"36da",x"3bfe",x"a8f0",x"0000",x"3bea",x"39c8",x"3a2d",x"4042",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"39be",x"3a2f",x"404d",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"39bf"),
(x"351b",x"403f",x"36da",x"350e",x"bb96",x"0000",x"3a50",x"3b98",x"351b",x"403f",x"3710",x"3664",x"bb55",x"0000",x"3a5a",x"3b98",x"353f",x"4041",x"3710",x"3746",x"bb1f",x"0000",x"3a5a",x"3ba0"),
(x"3a27",x"4059",x"36da",x"a3ae",x"3bff",x"0000",x"3a2d",x"3bb3",x"3a27",x"4059",x"3710",x"a3ef",x"3bff",x"9818",x"3a23",x"3bb3",x"39f5",x"4059",x"3710",x"a4e3",x"3bff",x"1818",x"3a23",x"3b9f"),
(x"386d",x"4039",x"36da",x"bba8",x"b4a3",x"8000",x"3a72",x"3adc",x"386d",x"4039",x"3710",x"bac4",x"b844",x"0000",x"3a7c",x"3adc",x"3877",x"4037",x"3710",x"b74e",x"bb1d",x"8000",x"3a7c",x"3ae1"),
(x"3885",x"404c",x"36da",x"b305",x"3bce",x"0000",x"3a8b",x"3b1c",x"3885",x"404c",x"3710",x"b25f",x"3bd7",x"8000",x"3a96",x"3b1c",x"382a",x"404d",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b3e"),
(x"3501",x"403e",x"36da",x"ada8",x"bbf8",x"8000",x"3a50",x"3b93",x"3501",x"403e",x"3710",x"2d0c",x"bbf9",x"0000",x"3a5a",x"3b93",x"351b",x"403f",x"3710",x"3664",x"bb55",x"0000",x"3a5a",x"3b98"),
(x"386c",x"403c",x"36da",x"bb38",x"36e2",x"868d",x"3a72",x"3ad8",x"386c",x"403c",x"3710",x"bbdd",x"31e1",x"0000",x"3a7c",x"3ad8",x"386d",x"4039",x"3710",x"bac4",x"b844",x"0000",x"3a7c",x"3adc"),
(x"382a",x"404d",x"36da",x"2f40",x"3bf2",x"8000",x"3a8b",x"3b3e",x"382a",x"404d",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b3e",x"3813",x"404e",x"3710",x"a8bf",x"3bfe",x"8000",x"3a96",x"3b47"),
(x"3a25",x"4041",x"36da",x"367a",x"bb50",x"0000",x"3b21",x"387e",x"3a25",x"4041",x"3710",x"3700",x"bb23",x"2f05",x"3b1b",x"3887",x"3a2d",x"4042",x"3710",x"3644",x"bb4c",x"2f83",x"3b19",x"3884"),
(x"3a25",x"3d5c",x"3710",x"3bd6",x"2604",x"3256",x"3a49",x"33c0",x"3a26",x"3d45",x"3710",x"3bcf",x"2680",x"32dc",x"3a36",x"33ca",x"3a20",x"3d45",x"3732",x"3b18",x"2439",x"3763",x"3a35",x"33aa"),
(x"3a1f",x"3d5c",x"3733",x"3b23",x"251e",x"3737",x"3a49",x"339f",x"3a20",x"3d45",x"3732",x"3b18",x"2439",x"3763",x"3a35",x"33aa",x"3a19",x"3d45",x"3749",x"3871",x"2587",x"3aa6",x"3a35",x"3392"),
(x"3a18",x"3d5c",x"3748",x"36c9",x"29dc",x"3b3c",x"3a48",x"3388",x"3a19",x"3d45",x"3749",x"3871",x"2587",x"3aa6",x"3a35",x"3392",x"3a14",x"3d45",x"374e",x"2fa2",x"2997",x"3bef",x"3a34",x"3387"),
(x"3a10",x"3d5c",x"3749",x"b4de",x"2b76",x"3b9b",x"3a48",x"337b",x"3a14",x"3d45",x"374e",x"2fa2",x"2997",x"3bef",x"3a34",x"3387",x"3a0d",x"3d45",x"374b",x"b745",x"2966",x"3b1e",x"3a34",x"337b"),
(x"3a09",x"3d5c",x"373b",x"b7a6",x"3a67",x"35ca",x"3bbd",x"39cf",x"39fc",x"3d5d",x"3713",x"af5f",x"3bdb",x"30c1",x"3bc3",x"39d6",x"3a03",x"3d5d",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bc0",x"39d7"),
(x"3a09",x"3d5e",x"373a",x"baf6",x"2b34",x"37d2",x"3bbc",x"39cf",x"3a11",x"3d5e",x"374a",x"b547",x"b37e",x"3b50",x"3bb9",x"39cc",x"3a10",x"3d5c",x"3749",x"b3aa",x"a4b5",x"3bc3",x"3bbb",x"39cb"),
(x"39fc",x"3d45",x"3710",x"ba72",x"9a8d",x"38bc",x"3a34",x"333e",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e",x"3a02",x"3d45",x"3724",x"bb1f",x"1a24",x"3747",x"3a34",x"3352"),
(x"3a02",x"3d73",x"3711",x"bbe1",x"a6cf",x"3179",x"3bfb",x"396f",x"3a04",x"3d73",x"3727",x"bbc5",x"a8fd",x"3377",x"3bfb",x"3974",x"3a03",x"3d5d",x"370e",x"bbc2",x"ab4f",x"338c",x"3bea",x"3970"),
(x"3a08",x"3d73",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"3978",x"3a0f",x"3d72",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"397c",x"3a11",x"3d5e",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"397d"),
(x"3a0f",x"3d72",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"397c",x"3a17",x"3d72",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3bfb",x"397f",x"3a19",x"3d5e",x"374d",x"3400",x"aa73",x"3bbc",x"3beb",x"3980"),
(x"3a1d",x"3d72",x"374d",x"3802",x"a90b",x"3aea",x"3bfb",x"3982",x"3a21",x"3d5e",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"3984",x"3a19",x"3d5e",x"374d",x"3400",x"aa73",x"3bbc",x"3beb",x"3980"),
(x"3a24",x"3d72",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"3986",x"3a25",x"3d5e",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"3986",x"3a21",x"3d5e",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"3984"),
(x"3a2a",x"3d73",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"398b",x"3a2d",x"3d5e",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"398f",x"3a25",x"3d5e",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"3986"),
(x"3a2d",x"3d5e",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"398f",x"3a2a",x"3d73",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"398b",x"3a2f",x"3d73",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"398f"),
(x"3a25",x"3d5e",x"3738",x"36f3",x"bae7",x"3422",x"3bb7",x"39c3",x"3a2d",x"3d5e",x"3710",x"3644",x"bb4c",x"2f83",x"3bba",x"39ba",x"3a25",x"3d5c",x"3710",x"3700",x"bb23",x"2f05",x"3bbd",x"39bd"),
(x"3a0d",x"3d45",x"374b",x"b745",x"2966",x"3b1e",x"3a34",x"337b",x"3a07",x"3d45",x"373c",x"bac4",x"2853",x"3841",x"3a34",x"336a",x"3a09",x"3d5c",x"373b",x"b9d7",x"2404",x"3976",x"3a48",x"3369"),
(x"3a11",x"3d5e",x"374a",x"b547",x"b37e",x"3b50",x"3bb9",x"39cc",x"3a19",x"3d5e",x"374d",x"3243",x"b807",x"3aba",x"3bb8",x"39c9",x"3a18",x"3d5c",x"3748",x"291b",x"b8de",x"3a57",x"3bba",x"39c9"),
(x"3a18",x"3d5c",x"3748",x"291b",x"b8de",x"3a57",x"3bba",x"39c9",x"3a19",x"3d5e",x"374d",x"3243",x"b807",x"3aba",x"3bb8",x"39c9",x"3a21",x"3d5e",x"3744",x"37e0",x"ba17",x"36be",x"3bb7",x"39c5"),
(x"3a25",x"3d5e",x"3738",x"36f3",x"bae7",x"3422",x"3bb7",x"39c3",x"3a1f",x"3d5c",x"3733",x"37ff",x"ba99",x"3438",x"3bba",x"39c3",x"3a21",x"3d5e",x"3744",x"37e0",x"ba17",x"36be",x"3bb7",x"39c5"),
(x"3a2a",x"3d73",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3843",x"3a20",x"3d74",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3849",x"3a26",x"3d74",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3842"),
(x"3a24",x"3d72",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3848",x"3a1a",x"3d74",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"384d",x"3a20",x"3d74",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3849"),
(x"3a1d",x"3d72",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"384c",x"3a15",x"3d74",x"374b",x"aaa7",x"39a6",x"39a5",x"3b22",x"384f",x"3a1a",x"3d74",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"384d"),
(x"3a17",x"3d72",x"3751",x"2fda",x"39a6",x"3994",x"3b24",x"384f",x"3a15",x"3d74",x"374b",x"aaa7",x"39a6",x"39a5",x"3b22",x"384f",x"3a1d",x"3d72",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"384c"),
(x"3a0f",x"3d72",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3851",x"3a0f",x"3d74",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3851",x"3a15",x"3d74",x"374b",x"aaa7",x"39a6",x"39a5",x"3b22",x"384f"),
(x"3a08",x"3d73",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3854",x"3a09",x"3d74",x"373e",x"ba28",x"9dd6",x"391a",x"3b1e",x"3853",x"3a0f",x"3d74",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3851"),
(x"3a04",x"3d73",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3857",x"3a01",x"3d74",x"371c",x"b97b",x"b976",x"340b",x"3b19",x"3857",x"3a09",x"3d74",x"373e",x"ba28",x"9dd6",x"391a",x"3b1e",x"3853"),
(x"3a02",x"3d73",x"3711",x"b40d",x"bb3a",x"3585",x"3b18",x"385a",x"3a01",x"3d74",x"371c",x"b97b",x"b976",x"340b",x"3b19",x"3857",x"3a04",x"3d73",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3857"),
(x"3a02",x"3d73",x"3711",x"b40d",x"bb3a",x"3585",x"3b18",x"385a",x"39fb",x"3d73",x"3713",x"aeda",x"bb7b",x"3565",x"3b16",x"3858",x"3a01",x"3d74",x"371c",x"b97b",x"b976",x"340b",x"3b19",x"3857"),
(x"3a02",x"3d73",x"3711",x"315a",x"2bae",x"3bdf",x"3a5b",x"3349",x"3a03",x"3d5d",x"370e",x"34eb",x"a6e9",x"3b9c",x"3a49",x"334b",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e"),
(x"3a24",x"3d8b",x"372b",x"3b86",x"a8a8",x"3564",x"3a6f",x"33b1",x"3a27",x"3d8b",x"3710",x"3bea",x"a4d6",x"30a2",x"3a6f",x"33c9",x"3a26",x"3d74",x"3710",x"3bed",x"a7ae",x"3024",x"3a5b",x"33c4"),
(x"3a24",x"3d8b",x"372b",x"3b86",x"a8a8",x"3564",x"3a6f",x"33b1",x"3a20",x"3d74",x"3739",x"3abd",x"a8b5",x"384c",x"3a5c",x"339e",x"3a21",x"3d8b",x"373a",x"3acd",x"a5ae",x"3834",x"3a6f",x"33a3"),
(x"3a20",x"3d74",x"3739",x"3abd",x"a8b5",x"384c",x"3a5c",x"339e",x"3a1a",x"3d74",x"3746",x"38a5",x"a839",x"3a81",x"3a5c",x"338e",x"3a1a",x"3d8a",x"3749",x"38cd",x"a812",x"3a64",x"3a6f",x"3391"),
(x"3a15",x"3d74",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a5c",x"3385",x"3a14",x"3d8a",x"374f",x"32be",x"a89e",x"3bd0",x"3a6f",x"3385",x"3a1a",x"3d8a",x"3749",x"38cd",x"a812",x"3a64",x"3a6f",x"3391"),
(x"3a0f",x"3d74",x"3749",x"b771",x"a91b",x"3b13",x"3a5c",x"3379",x"3a0d",x"3d8a",x"374b",x"b6cb",x"a758",x"3b3d",x"3a6f",x"3378",x"3a14",x"3d8a",x"374f",x"32be",x"a89e",x"3bd0",x"3a6f",x"3385"),
(x"3a09",x"3d74",x"373e",x"ba21",x"a786",x"3921",x"3a5c",x"336a",x"3a07",x"3d8a",x"373c",x"baa0",x"a6bb",x"3879",x"3a6f",x"3366",x"3a0d",x"3d8a",x"374b",x"b6cb",x"a758",x"3b3d",x"3a6f",x"3378"),
(x"3a09",x"3d74",x"373e",x"ba21",x"a786",x"3921",x"3a5c",x"336a",x"3a01",x"3d74",x"371c",x"b9f4",x"a495",x"3957",x"3a5c",x"334a",x"3a00",x"3d8a",x"3722",x"ba6c",x"a860",x"38c2",x"3a6f",x"334c"),
(x"3a01",x"3d74",x"371c",x"b9f4",x"a495",x"3957",x"3a5c",x"334a",x"39fb",x"3d73",x"3713",x"a9a5",x"a460",x"3bfd",x"3a5b",x"333d",x"39fc",x"3d8a",x"3718",x"b8fc",x"a86a",x"3a40",x"3a6f",x"3340"),
(x"3475",x"3d6c",x"3710",x"0000",x"0000",x"3c00",x"3a55",x"2451",x"3485",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"24c1",x"3485",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"24c1"),
(x"3485",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"24c1",x"349b",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"255f",x"349b",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"255f"),
(x"349b",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"255f",x"349b",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"255f",x"34bb",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2643"),
(x"34bb",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2643",x"34cb",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"26b3",x"34cb",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"26b3"),
(x"34cb",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"26b3",x"34e9",x"3d79",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"278b",x"34e9",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"278b"),
(x"34e9",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"278b",x"34e9",x"3d79",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"278b",x"3501",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"281a"),
(x"3501",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"281a",x"351b",x"3d79",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2878",x"351b",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2878"),
(x"351b",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2878",x"351b",x"3d79",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2878",x"353f",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"28fb"),
(x"353f",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"28fb",x"3555",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2949",x"3555",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2949"),
(x"3555",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2949",x"357d",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a58",x"29d7",x"357d",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4b",x"29d7"),
(x"357d",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4b",x"29d7",x"357d",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a58",x"29d7",x"3592",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2a20"),
(x"363b",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2c3f",x"363b",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2c3f",x"36f7",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2d8d"),
(x"363b",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2c3f",x"362c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2c23",x"362c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2c23"),
(x"362c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2c23",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b",x"3592",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2a20"),
(x"35f5",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2b84",x"35fd",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2ba0",x"35fd",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"2ba0"),
(x"35e4",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2b48",x"35fd",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"2ba0",x"35f3",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2b7d"),
(x"35d3",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2b0a",x"35f3",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2b7d",x"35f1",x"3d7d",x"3710",x"868d",x"0cea",x"3c00",x"3a63",x"2b76"),
(x"35f5",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2b84",x"35e4",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2b48",x"35fd",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2ba0"),
(x"35e4",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2b48",x"35d3",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2b0a",x"35f3",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2b7d"),
(x"35d3",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2b0a",x"35bd",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2aba",x"35f1",x"3d53",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2b76"),
(x"35bd",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2aba",x"359e",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2a4d",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b"),
(x"35bd",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2aba",x"35f1",x"3d7d",x"3710",x"868d",x"0cea",x"3c00",x"3a63",x"2b76",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"3587",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5e",x"29f9",x"358a",x"3d7c",x"3710",x"0000",x"0000",x"3c00",x"3a63",x"2a04",x"3593",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2a22"),
(x"36f7",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2d8d",x"3710",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2dbb",x"3710",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2dbb"),
(x"380a",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2f8b",x"37b8",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2ee7",x"37b8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2ee7"),
(x"37b8",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2ee7",x"37a8",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2ec9",x"37a8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ec9"),
(x"37a8",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2ec9",x"378c",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2e97",x"378c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2e97"),
(x"378c",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2e97",x"376c",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2e5e",x"376c",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2e5e"),
(x"376c",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2e5e",x"376c",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2e5e",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"36f7",x"3d8e",x"3710",x"0000",x"0000",x"3c00",x"3a72",x"2d8e",x"3716",x"3d8d",x"3710",x"0000",x"0000",x"3c00",x"3a72",x"2dc4",x"36df",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"2d63"),
(x"3716",x"3d8d",x"3710",x"0000",x"0000",x"3c00",x"3a72",x"2dc4",x"372e",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"2df0",x"36dc",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2d5e"),
(x"36df",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"2d63",x"3716",x"3d42",x"3710",x"0000",x"0000",x"3c00",x"3a31",x"2dc4",x"36f7",x"3d41",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e"),
(x"36dc",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2d5e",x"372e",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2df0",x"3716",x"3d42",x"3710",x"0000",x"0000",x"3c00",x"3a31",x"2dc4"),
(x"3753",x"3d46",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"2e32",x"3742",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2e14",x"375f",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2e47"),
(x"3742",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2e14",x"372e",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2df0",x"3754",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"2e33"),
(x"3753",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"2e32",x"3760",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2e49",x"375f",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2e47"),
(x"3742",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"2e14",x"375f",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2e47",x"3754",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"2e33"),
(x"36cb",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2d40",x"36c2",x"3d7c",x"3710",x"0000",x"0000",x"3c00",x"3a63",x"2d2f",x"36c4",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2d33"),
(x"36cb",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2d40",x"3705",x"3d58",x"3710",x"0000",x"0000",x"3c00",x"3a44",x"2da6",x"36c4",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2d33"),
(x"3705",x"3d58",x"3710",x"0000",x"0000",x"3c00",x"3a44",x"2da6",x"3713",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2dbf",x"36dc",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2d5e"),
(x"3705",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5f",x"2da6",x"36c4",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2d33",x"36dc",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2d5e"),
(x"3713",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2dbf",x"36dc",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2d5e",x"372e",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"2df0"),
(x"372e",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2df0",x"36dc",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2d5e",x"3713",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2dbf"),
(x"3713",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2dbf",x"3754",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"2e33",x"3752",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2e30"),
(x"3713",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2dbf",x"3716",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2dc5",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"3710",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2dbb",x"3710",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2dbb",x"3716",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2dc5"),
(x"3716",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2dc5",x"3752",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2e30",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"380a",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2f8b",x"3813",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2fac",x"3813",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2fac"),
(x"382a",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ffc",x"382a",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2ffc",x"3813",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2fac"),
(x"382a",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ffc",x"3885",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"30a2",x"3885",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"30a2"),
(x"388c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"30ad",x"388c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"30ad",x"3885",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"30a2"),
(x"38d5",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"3130",x"38bf",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"3109",x"38bf",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"3109"),
(x"38bf",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"3109",x"38bf",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"3109",x"38b2",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30f1"),
(x"38b2",x"3d76",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"30f1",x"38b2",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30f1",x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed"),
(x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed",x"388c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"30ad",x"388c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"30ad"),
(x"3872",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"3080",x"3877",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"3088",x"386d",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"3076"),
(x"3885",x"3d59",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30a2",x"3894",x"3d44",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30bc",x"3877",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"3088"),
(x"386d",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"3076",x"3877",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"3088",x"3872",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"3080"),
(x"3877",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"3088",x"3894",x"3d8c",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"30bc",x"3885",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5e",x"30a2"),
(x"3894",x"3d8c",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"30bc",x"38b7",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"30f9",x"388c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"30ae"),
(x"388c",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"30ae",x"38b7",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30f9",x"3894",x"3d44",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30bc"),
(x"38d8",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"3135",x"38c7",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3117",x"38d4",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3d",x"312d"),
(x"38d8",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"3135",x"38d9",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a68",x"3136",x"38d4",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"312d"),
(x"38c7",x"3d87",x"3710",x"0000",x"0000",x"3c00",x"3a6c",x"3117",x"38d4",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"312d",x"38c9",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"311a"),
(x"38c7",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3117",x"38b7",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30f9",x"38c9",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"311a"),
(x"388c",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"30ae",x"388c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"30ad",x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed"),
(x"388c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"30ae",x"38b2",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"30f2",x"38b0",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"30ed"),
(x"38b2",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"30f2",x"38b7",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30f9",x"388c",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"30ae"),
(x"38b7",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"30f9",x"38b2",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"30f2",x"388c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"30ae"),
(x"38f6",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"316b",x"38f6",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"316b",x"38d5",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"3130"),
(x"3915",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"31a2",x"3915",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"31a2",x"38f6",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"316b"),
(x"392f",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"31d0",x"392f",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"31d0",x"3915",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"31a2"),
(x"393f",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"31ed",x"393f",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"31ed",x"392f",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"31d0"),
(x"3953",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3211",x"3953",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3211",x"393f",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"31ed"),
(x"395a",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"321d",x"395a",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"321d",x"3953",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3211"),
(x"395d",x"3d81",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"3222",x"395d",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"3222",x"395a",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"321d"),
(x"395d",x"3d81",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"3222",x"3963",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"322d",x"3963",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"322d"),
(x"3972",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"3248",x"3972",x"3d50",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"3248",x"3963",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"322d"),
(x"3985",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"3269",x"3985",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"3269",x"3972",x"3d50",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"3248"),
(x"3994",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3284",x"3994",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3284",x"3985",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"3269"),
(x"3999",x"3d89",x"3710",x"935f",x"1e0a",x"3c00",x"3a6e",x"328d",x"3999",x"3d47",x"3710",x"96f6",x"9f93",x"3c00",x"3a35",x"328d",x"3994",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3284"),
(x"3999",x"3d89",x"3710",x"935f",x"1e0a",x"3c00",x"3a6e",x"328d",x"39fb",x"3d73",x"3713",x"a9a5",x"a460",x"3bfd",x"3a5b",x"333d",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e"),
(x"39f5",x"3d8a",x"3710",x"b60a",x"25b5",x"3b67",x"3a6f",x"3331",x"39fc",x"3d8a",x"3718",x"b8fc",x"a86a",x"3a40",x"3a6f",x"3340",x"39fb",x"3d73",x"3713",x"a9a5",x"a460",x"3bfd",x"3a5b",x"333d"),
(x"3999",x"3d47",x"3710",x"96f6",x"9f93",x"3c00",x"3a35",x"328d",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e",x"39fc",x"3d45",x"3710",x"ba72",x"9a8d",x"38bc",x"3a34",x"333e"),
(x"3a0d",x"3d8a",x"374b",x"a412",x"3bfd",x"2966",x"3bc0",x"3a1e",x"3a07",x"3d8a",x"373c",x"a752",x"3bff",x"9bfc",x"3bc3",x"3a1b",x"3a1a",x"3d8a",x"3749",x"a2b5",x"3bfe",x"2818",x"3bc0",x"3a23"),
(x"3a07",x"3d8a",x"373c",x"a752",x"3bff",x"9bfc",x"3bc3",x"3a1b",x"3a00",x"3d8a",x"3722",x"23fc",x"3bf8",x"2d56",x"3bc8",x"3a19",x"3a21",x"3d8b",x"373a",x"a884",x"3bfe",x"2546",x"3bc3",x"3a25"),
(x"3a00",x"3d8a",x"3722",x"23fc",x"3bf8",x"2d56",x"3bc8",x"3a19",x"39fc",x"3d8a",x"3718",x"135f",x"3bfd",x"29a1",x"3bc9",x"3a17",x"3a24",x"3d8b",x"372b",x"a504",x"3bff",x"9a24",x"3bc6",x"3a27"),
(x"39fc",x"3d8a",x"3718",x"135f",x"3bfd",x"29a1",x"3bc9",x"3a17",x"39f5",x"3d8a",x"3710",x"a4e3",x"3bff",x"1818",x"3bcb",x"3a14",x"3a27",x"3d8b",x"3710",x"a3ef",x"3bff",x"9818",x"3bcb",x"3a28"),
(x"3a19",x"3d45",x"3749",x"209b",x"bc00",x"135f",x"3a5a",x"3a5e",x"3a07",x"3d45",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a57",x"3a57",x"3a0d",x"3d45",x"374b",x"1481",x"bbff",x"26a7",x"3a5a",x"3a5a"),
(x"3a20",x"3d45",x"3732",x"1f93",x"bc00",x"975f",x"3a55",x"3a61",x"3a02",x"3d45",x"3724",x"1c81",x"bbff",x"a1d6",x"3a53",x"3a55",x"3a07",x"3d45",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a57",x"3a57"),
(x"3a26",x"3d45",x"3710",x"1f5f",x"bbff",x"a032",x"3a4f",x"3a63",x"39fc",x"3d45",x"3710",x"9bc8",x"bc00",x"200b",x"3a4f",x"3a53",x"3a02",x"3d45",x"3724",x"1c81",x"bbff",x"a1d6",x"3a53",x"3a55"),
(x"34e9",x"3d56",x"36da",x"b698",x"bb49",x"8000",x"3a5f",x"3b8f",x"34e9",x"3d56",x"3710",x"b50d",x"bb97",x"0000",x"3a6a",x"3b8f",x"3501",x"3d55",x"3710",x"2d0c",x"bbf9",x"0000",x"3a6a",x"3b94"),
(x"3872",x"3d54",x"36da",x"b902",x"3a3c",x"0000",x"3a33",x"39d2",x"3872",x"3d54",x"3710",x"b9d1",x"397d",x"8000",x"3a3e",x"39d2",x"386c",x"3d51",x"3710",x"bbdd",x"31e1",x"0000",x"3a3e",x"39d5"),
(x"3813",x"3d74",x"36da",x"27fc",x"3bfe",x"0000",x"3a3d",x"3b80",x"3813",x"3d74",x"3710",x"a8bf",x"3bfe",x"8000",x"3a32",x"3b80",x"380a",x"3d74",x"3710",x"ae12",x"3bf6",x"0000",x"3a32",x"3b7d"),
(x"34cb",x"3d5b",x"36da",x"b501",x"bb99",x"0000",x"3a5f",x"3b88",x"34cb",x"3d5b",x"3710",x"b64c",x"bb5a",x"0000",x"3a6a",x"3b88",x"34e9",x"3d56",x"3710",x"b50d",x"bb97",x"0000",x"3a6a",x"3b8f"),
(x"39fc",x"3d45",x"36da",x"a111",x"bc00",x"0000",x"3a44",x"3a53",x"39fc",x"3d45",x"3710",x"9bc8",x"bc00",x"200b",x"3a4f",x"3a53",x"3a26",x"3d45",x"3710",x"1f5f",x"bbff",x"a032",x"3a4f",x"3a63"),
(x"3885",x"3d59",x"36da",x"b83d",x"3ac8",x"0000",x"3a33",x"39ca",x"3885",x"3d59",x"3710",x"b7eb",x"3af3",x"0000",x"3a3e",x"39ca",x"3872",x"3d54",x"3710",x"b9d1",x"397d",x"8000",x"3a3e",x"39d2"),
(x"375f",x"3d83",x"36da",x"3b14",x"b774",x"068d",x"3a3d",x"3b4e",x"375f",x"3d83",x"3710",x"3bc1",x"b3d7",x"868d",x"3a32",x"3b4e",x"3760",x"3d86",x"3710",x"3b92",x"3528",x"8000",x"3a32",x"3b4c"),
(x"34bb",x"3d5c",x"36da",x"b141",x"bbe4",x"0000",x"3a5f",x"3b85",x"34bb",x"3d5c",x"3710",x"b31c",x"bbcc",x"0000",x"3a6a",x"3b85",x"34cb",x"3d5b",x"3710",x"b64c",x"bb5a",x"0000",x"3a6a",x"3b88"),
(x"388c",x"3d5b",x"36da",x"bbfd",x"29ab",x"0000",x"3a33",x"39c7",x"388c",x"3d5b",x"3710",x"bb54",x"3669",x"8000",x"3a3e",x"39c7",x"3885",x"3d59",x"3710",x"b7eb",x"3af3",x"0000",x"3a3e",x"39ca"),
(x"380a",x"3d74",x"36da",x"ad56",x"3bf8",x"8000",x"3a3d",x"3b7d",x"380a",x"3d74",x"3710",x"ae12",x"3bf6",x"0000",x"3a32",x"3b7d",x"37b8",x"3d71",x"3710",x"30d0",x"3be8",x"0000",x"3a32",x"3b6a"),
(x"349b",x"3d5d",x"36da",x"b4a8",x"bba7",x"8000",x"3a5f",x"3b7f",x"349b",x"3d5d",x"3710",x"b221",x"bbda",x"0000",x"3a6a",x"3b7f",x"34bb",x"3d5c",x"3710",x"b31c",x"bbcc",x"0000",x"3a6a",x"3b85"),
(x"388c",x"3d5d",x"36da",x"b967",x"b9e6",x"0000",x"3a33",x"39c5",x"388c",x"3d5d",x"3710",x"bb52",x"b671",x"0000",x"3a3e",x"39c5",x"388c",x"3d5b",x"3710",x"bb54",x"3669",x"8000",x"3a3e",x"39c7"),
(x"37b8",x"3d71",x"36da",x"2df5",x"3bf7",x"8000",x"3a3d",x"3b6a",x"37b8",x"3d71",x"3710",x"30d0",x"3be8",x"0000",x"3a32",x"3b6a",x"37a8",x"3d71",x"3710",x"3580",x"3b83",x"0000",x"3a32",x"3b67"),
(x"3485",x"3d5f",x"36da",x"b92c",x"ba1a",x"8000",x"3a5f",x"3b7b",x"3485",x"3d5f",x"3710",x"b819",x"bade",x"868d",x"3a6a",x"3b7b",x"349b",x"3d5d",x"3710",x"b221",x"bbda",x"0000",x"3a6a",x"3b7f"),
(x"3885",x"3d5e",x"36da",x"b25f",x"bbd7",x"0000",x"3a0c",x"3b9a",x"3885",x"3d5e",x"3710",x"b305",x"bbce",x"0000",x"3a17",x"3b9a",x"388c",x"3d5d",x"3710",x"bb52",x"b671",x"0000",x"3a17",x"3b9c"),
(x"37a8",x"3d71",x"36da",x"33d5",x"3bc1",x"0000",x"3a3d",x"3b67",x"37a8",x"3d71",x"3710",x"3580",x"3b83",x"0000",x"3a32",x"3b67",x"378c",x"3d75",x"3710",x"3688",x"3b4d",x"8000",x"3a32",x"3b60"),
(x"3a2f",x"3d73",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"3838",x"3a2f",x"3d73",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"383f",x"3a26",x"3d74",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3842"),
(x"3475",x"3d64",x"36da",x"bbab",x"b48e",x"0000",x"3a5f",x"3b76",x"3475",x"3d64",x"3710",x"baeb",x"b803",x"068d",x"3a6a",x"3b76",x"3485",x"3d5f",x"3710",x"b819",x"bade",x"868d",x"3a6a",x"3b7b"),
(x"3753",x"3d46",x"36da",x"37e4",x"baf5",x"8000",x"3a0c",x"3b39",x"3753",x"3d46",x"3710",x"38fe",x"ba3f",x"0000",x"3a17",x"3b39",x"3760",x"3d4a",x"3710",x"3bfa",x"acac",x"8000",x"3a17",x"3b3c"),
(x"378c",x"3d75",x"36da",x"373a",x"3b23",x"0000",x"3a3d",x"3b60",x"378c",x"3d75",x"3710",x"3688",x"3b4d",x"8000",x"3a32",x"3b60",x"376c",x"3d78",x"3710",x"3899",x"3a8b",x"0000",x"3a32",x"3b5a"),
(x"382a",x"3d5d",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b77",x"382a",x"3d5d",x"3710",x"2f41",x"bbf2",x"0000",x"3a17",x"3b77",x"3885",x"3d5e",x"3710",x"b305",x"bbce",x"0000",x"3a17",x"3b9a"),
(x"376c",x"3d78",x"36da",x"3787",x"3b0e",x"0000",x"3a3d",x"3b5a",x"376c",x"3d78",x"3710",x"3899",x"3a8b",x"0000",x"3a32",x"3b5a",x"3752",x"3d7e",x"3710",x"3bfd",x"aabe",x"0000",x"3a32",x"3b53"),
(x"3999",x"3d47",x"36da",x"b32b",x"bbcb",x"0000",x"3a44",x"3a2e",x"3999",x"3d47",x"3710",x"b2ba",x"bbd2",x"0000",x"3a4f",x"3a2e",x"39fc",x"3d45",x"3710",x"9bc8",x"bc00",x"200b",x"3a4f",x"3a53"),
(x"3813",x"3d5c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a0c",x"3b6e",x"3813",x"3d5c",x"3710",x"27fc",x"bbfe",x"0000",x"3a17",x"3b6e",x"382a",x"3d5d",x"3710",x"2f41",x"bbf2",x"0000",x"3a17",x"3b77"),
(x"3753",x"3d89",x"36da",x"38fe",x"3a3f",x"8000",x"3a3d",x"3b48",x"3753",x"3d89",x"3710",x"37e4",x"3af5",x"8000",x"3a32",x"3b48",x"3742",x"3d8b",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b44"),
(x"380a",x"3d5c",x"36da",x"ae12",x"bbf6",x"0000",x"3a0c",x"3b6b",x"380a",x"3d5c",x"3710",x"ad54",x"bbf8",x"0000",x"3a17",x"3b6b",x"3813",x"3d5c",x"3710",x"27fc",x"bbfe",x"0000",x"3a17",x"3b6e"),
(x"3742",x"3d8b",x"36da",x"342c",x"3bb9",x"8000",x"3a3d",x"3b44",x"3742",x"3d8b",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b44",x"372e",x"3d8b",x"3710",x"338a",x"3bc6",x"0000",x"3a32",x"3b40"),
(x"3760",x"3d4a",x"36da",x"3b92",x"b528",x"0000",x"3a0c",x"3b3c",x"3760",x"3d4a",x"3710",x"3bfa",x"acac",x"8000",x"3a17",x"3b3c",x"375f",x"3d4c",x"3710",x"3b14",x"3774",x"8000",x"3a17",x"3b3e"),
(x"372e",x"3d8b",x"36da",x"2fc6",x"3bf0",x"0000",x"3a3d",x"3b40",x"372e",x"3d8b",x"3710",x"338a",x"3bc6",x"0000",x"3a32",x"3b40",x"3716",x"3d8d",x"3710",x"32c2",x"3bd1",x"8000",x"3a32",x"3b3b"),
(x"37b8",x"3d5f",x"36da",x"30d0",x"bbe8",x"0000",x"3a0c",x"3b59",x"37b8",x"3d5f",x"3710",x"2df5",x"bbf7",x"0000",x"3a17",x"3b59",x"380a",x"3d5c",x"3710",x"ad54",x"bbf8",x"0000",x"3a17",x"3b6b"),
(x"3716",x"3d8d",x"36da",x"34b5",x"3ba5",x"8000",x"3a3d",x"3b3b",x"3716",x"3d8d",x"3710",x"32c2",x"3bd1",x"8000",x"3a32",x"3b3b",x"36f7",x"3d8e",x"3710",x"b463",x"3bb1",x"8000",x"3a32",x"3b35"),
(x"37a8",x"3d5e",x"36da",x"3580",x"bb83",x"0000",x"3a0c",x"3b56",x"37a8",x"3d5e",x"3710",x"33d5",x"bbc1",x"0000",x"3a17",x"3b56",x"37b8",x"3d5f",x"3710",x"2df5",x"bbf7",x"0000",x"3a17",x"3b59"),
(x"36f7",x"3d8e",x"36da",x"ae6b",x"3bf5",x"0000",x"3a3d",x"3b35",x"36f7",x"3d8e",x"3710",x"b463",x"3bb1",x"8000",x"3a32",x"3b35",x"36e3",x"3d8c",x"3710",x"bb17",x"3766",x"0000",x"3a32",x"3b31"),
(x"378c",x"3d5a",x"36da",x"3688",x"bb4d",x"8000",x"3a0c",x"3b50",x"378c",x"3d5a",x"3710",x"373a",x"bb23",x"0000",x"3a17",x"3b50",x"37a8",x"3d5e",x"3710",x"33d5",x"bbc1",x"0000",x"3a17",x"3b56"),
(x"36e3",x"3d8c",x"36da",x"b9b5",x"399a",x"0000",x"3a3d",x"3b31",x"36e3",x"3d8c",x"3710",x"bb17",x"3766",x"0000",x"3a32",x"3b31",x"36df",x"3d89",x"3710",x"bbc6",x"338f",x"8000",x"3a32",x"3b2e"),
(x"376c",x"3d57",x"36da",x"3899",x"ba8b",x"0000",x"3a0c",x"3b4a",x"376c",x"3d57",x"3710",x"3787",x"bb0e",x"0000",x"3a17",x"3b4a",x"378c",x"3d5a",x"3710",x"373a",x"bb23",x"0000",x"3a17",x"3b50"),
(x"36df",x"3d89",x"36da",x"bbbc",x"3412",x"0000",x"3a3d",x"3b2e",x"36df",x"3d89",x"3710",x"bbc6",x"338f",x"8000",x"3a32",x"3b2e",x"36dc",x"3d86",x"3710",x"bb3a",x"36d9",x"0000",x"3a32",x"3b2c"),
(x"3a26",x"3d74",x"36da",x"3bff",x"a4d0",x"0000",x"3a5a",x"33f3",x"3a26",x"3d74",x"3710",x"3bed",x"a7ae",x"3024",x"3a5b",x"33c4",x"3a27",x"3d8b",x"3710",x"3bea",x"a4d6",x"30a2",x"3a6f",x"33c9"),
(x"39f5",x"3d8a",x"36da",x"a49b",x"3bff",x"8000",x"3bd5",x"3a14",x"39f5",x"3d8a",x"3710",x"a4e3",x"3bff",x"1818",x"3bcb",x"3a14",x"3999",x"3d89",x"3710",x"b329",x"3bcb",x"8000",x"3bcb",x"39f0"),
(x"3752",x"3d51",x"36da",x"3bfd",x"2ac2",x"0000",x"3a0c",x"3b43",x"3752",x"3d51",x"3710",x"3be0",x"b1a3",x"868d",x"3a17",x"3b43",x"376c",x"3d57",x"3710",x"3787",x"bb0e",x"0000",x"3a17",x"3b4a"),
(x"36dc",x"3d86",x"36da",x"bba4",x"34ba",x"0000",x"3a3d",x"3b2c",x"36dc",x"3d86",x"3710",x"bb3a",x"36d9",x"0000",x"3a32",x"3b2c",x"36c4",x"3d7f",x"3710",x"bbc5",x"339b",x"0000",x"3a32",x"3b25"),
(x"3999",x"3d89",x"36da",x"b2b0",x"3bd2",x"0000",x"3bd5",x"39f0",x"3999",x"3d89",x"3710",x"b329",x"3bcb",x"8000",x"3bcb",x"39f0",x"3994",x"3d88",x"3710",x"b59f",x"3b7d",x"0000",x"3bcb",x"39ee"),
(x"3742",x"3d45",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b35",x"3742",x"3d45",x"3710",x"342c",x"bbb9",x"0000",x"3a17",x"3b35",x"3753",x"3d46",x"3710",x"38fe",x"ba3f",x"0000",x"3a17",x"3b39"),
(x"36c4",x"3d7f",x"36da",x"bb61",x"362a",x"0000",x"3a3d",x"3b25",x"36c4",x"3d7f",x"3710",x"bbc5",x"339b",x"0000",x"3a32",x"3b25",x"36c2",x"3d7c",x"3710",x"bafe",x"b7c2",x"868d",x"3a32",x"3b22"),
(x"3994",x"3d88",x"36da",x"b458",x"3bb2",x"8000",x"3bd5",x"39ee",x"3994",x"3d88",x"3710",x"b59f",x"3b7d",x"0000",x"3bcb",x"39ee",x"3985",x"3d84",x"3710",x"b796",x"3b0b",x"0000",x"3bcb",x"39e7"),
(x"372e",x"3d45",x"36da",x"338a",x"bbc6",x"0000",x"3a0c",x"3b31",x"372e",x"3d45",x"3710",x"2fc6",x"bbf0",x"0000",x"3a17",x"3b31",x"3742",x"3d45",x"3710",x"342c",x"bbb9",x"0000",x"3a17",x"3b35"),
(x"36c2",x"3d7c",x"36da",x"bbe7",x"b0ec",x"0000",x"3a3d",x"3b22",x"36c2",x"3d7c",x"3710",x"bafe",x"b7c2",x"868d",x"3a32",x"3b22",x"36cb",x"3d7a",x"3710",x"b86c",x"baaa",x"0000",x"3a32",x"3b20"),
(x"3985",x"3d84",x"36da",x"b817",x"3adf",x"0000",x"3bd5",x"39e7",x"3985",x"3d84",x"3710",x"b796",x"3b0b",x"0000",x"3bcb",x"39e7",x"3972",x"3d7f",x"3710",x"b0a0",x"3bea",x"0000",x"3bcb",x"39df"),
(x"3716",x"3d42",x"36da",x"32c2",x"bbd1",x"0000",x"3a0c",x"3b2c",x"3716",x"3d42",x"3710",x"34b5",x"bba5",x"0000",x"3a17",x"3b2c",x"372e",x"3d45",x"3710",x"2fc6",x"bbf0",x"0000",x"3a17",x"3b31"),
(x"36cb",x"3d7a",x"36da",x"b922",x"ba22",x"868d",x"3a3d",x"3b20",x"36cb",x"3d7a",x"3710",x"b86c",x"baaa",x"0000",x"3a32",x"3b20",x"3705",x"3d77",x"3710",x"b675",x"bb51",x"0000",x"3a32",x"3b14"),
(x"3972",x"3d7f",x"36da",x"b475",x"3bae",x"0000",x"3bd5",x"39df",x"3972",x"3d7f",x"3710",x"b0a0",x"3bea",x"0000",x"3bcb",x"39df",x"3963",x"3d7f",x"3710",x"36c5",x"3b3f",x"0000",x"3bcb",x"39d8"),
(x"36f7",x"3d41",x"36da",x"b463",x"bbb1",x"8000",x"3a0c",x"3b27",x"36f7",x"3d41",x"3710",x"ae6b",x"bbf5",x"0000",x"3a17",x"3b27",x"3716",x"3d42",x"3710",x"34b5",x"bba5",x"0000",x"3a17",x"3b2c"),
(x"3705",x"3d77",x"36da",x"b59a",x"bb7e",x"0000",x"3a3d",x"3b14",x"3705",x"3d77",x"3710",x"b675",x"bb51",x"0000",x"3a32",x"3b14",x"3713",x"3d75",x"3710",x"ba37",x"b909",x"0000",x"3a32",x"3b11"),
(x"3963",x"3d7f",x"36da",x"3420",x"3bba",x"0000",x"3bd5",x"39d8",x"3963",x"3d7f",x"3710",x"36c5",x"3b3f",x"0000",x"3bcb",x"39d8",x"395d",x"3d81",x"3710",x"3ac1",x"3849",x"0000",x"3bcb",x"39d5"),
(x"36e3",x"3d43",x"36da",x"bb17",x"b766",x"8000",x"3a0c",x"3b22",x"36e3",x"3d43",x"3710",x"b9b5",x"b99a",x"868d",x"3a17",x"3b22",x"36f7",x"3d41",x"3710",x"ae6b",x"bbf5",x"0000",x"3a17",x"3b27"),
(x"3713",x"3d75",x"36da",x"b972",x"b9db",x"8000",x"3a3d",x"3b11",x"3713",x"3d75",x"3710",x"ba37",x"b909",x"0000",x"3a32",x"3b11",x"3716",x"3d74",x"3710",x"bbad",x"3480",x"0000",x"3a32",x"3b10"),
(x"395d",x"3d81",x"36da",x"399d",x"39b2",x"0000",x"3bd5",x"39d5",x"395d",x"3d81",x"3710",x"3ac1",x"3849",x"0000",x"3bcb",x"39d5",x"395a",x"3d84",x"3710",x"3af1",x"37f3",x"0000",x"3bcb",x"39d3"),
(x"36df",x"3d47",x"36da",x"bbc6",x"b38f",x"8000",x"3a0c",x"3b20",x"36df",x"3d47",x"3710",x"bbbc",x"b412",x"0000",x"3a17",x"3b20",x"36e3",x"3d43",x"3710",x"b9b5",x"b99a",x"868d",x"3a17",x"3b22"),
(x"3716",x"3d74",x"36da",x"bbb8",x"b42d",x"0000",x"3b06",x"39ae",x"3716",x"3d74",x"3710",x"bbad",x"3480",x"0000",x"3b11",x"39ae",x"3710",x"3d73",x"3710",x"b80d",x"3ae5",x"0000",x"3b11",x"39af"),
(x"395a",x"3d84",x"36da",x"3b46",x"36a7",x"8000",x"3bd5",x"39d3",x"395a",x"3d84",x"3710",x"3af1",x"37f3",x"0000",x"3bcb",x"39d3",x"3953",x"3d88",x"3710",x"3857",x"3ab8",x"8000",x"3bcb",x"39ce"),
(x"36dc",x"3d4a",x"36da",x"bb3a",x"b6d9",x"0000",x"3a0c",x"3b1d",x"36dc",x"3d4a",x"3710",x"bba4",x"b4ba",x"0000",x"3a17",x"3b1d",x"36df",x"3d47",x"3710",x"bbbc",x"b412",x"0000",x"3a17",x"3b20"),
(x"3710",x"3d73",x"36da",x"b8f7",x"3a45",x"0000",x"3b06",x"39af",x"3710",x"3d73",x"3710",x"b80d",x"3ae5",x"0000",x"3b11",x"39af",x"36f7",x"3d72",x"3710",x"b05b",x"3bec",x"8000",x"3b11",x"39b4"),
(x"3475",x"3d6c",x"36da",x"baeb",x"3803",x"868d",x"3a5f",x"3b70",x"3475",x"3d6c",x"3710",x"bbab",x"348e",x"8000",x"3a6a",x"3b70",x"3475",x"3d64",x"3710",x"baeb",x"b803",x"068d",x"3a6a",x"3b76"),
(x"3953",x"3d88",x"36da",x"39a8",x"39a7",x"868d",x"3bd5",x"39ce",x"3953",x"3d88",x"3710",x"3857",x"3ab8",x"8000",x"3bcb",x"39ce",x"393f",x"3d8b",x"3710",x"b2bb",x"3bd2",x"868d",x"3bcb",x"39c6"),
(x"36c4",x"3d51",x"36da",x"bbc5",x"b39b",x"0000",x"3a0c",x"3b17",x"36c4",x"3d51",x"3710",x"bb61",x"b62a",x"0000",x"3a17",x"3b17",x"36dc",x"3d4a",x"3710",x"bba4",x"b4ba",x"0000",x"3a17",x"3b1d"),
(x"363b",x"3d72",x"36da",x"3439",x"3bb7",x"0000",x"3b06",x"39d8",x"363b",x"3d72",x"3710",x"34bd",x"3ba4",x"0000",x"3b11",x"39d8",x"362c",x"3d73",x"3710",x"3609",x"3b68",x"8000",x"3b11",x"39db"),
(x"3994",x"3d47",x"36da",x"b59f",x"bb7d",x"0000",x"3a44",x"3a2c",x"3994",x"3d47",x"3710",x"b458",x"bbb2",x"8000",x"3a4f",x"3a2c",x"3999",x"3d47",x"3710",x"b2ba",x"bbd2",x"0000",x"3a4f",x"3a2e"),
(x"393f",x"3d8b",x"36da",x"1cea",x"3c00",x"0000",x"3bd5",x"39c6",x"393f",x"3d8b",x"3710",x"b2bb",x"3bd2",x"868d",x"3bcb",x"39c6",x"392f",x"3d88",x"3710",x"b874",x"3aa4",x"0000",x"3bcb",x"39bf"),
(x"36c2",x"3d54",x"36da",x"baff",x"37c2",x"068d",x"3a0c",x"3b14",x"36c2",x"3d54",x"3710",x"bbe7",x"30ec",x"868d",x"3a17",x"3b14",x"36c4",x"3d51",x"3710",x"bb61",x"b62a",x"0000",x"3a17",x"3b17"),
(x"36f7",x"3d72",x"36da",x"b12d",x"3be4",x"0000",x"3b06",x"39b4",x"36f7",x"3d72",x"3710",x"b05b",x"3bec",x"8000",x"3b11",x"39b4",x"363b",x"3d72",x"3710",x"34bd",x"3ba4",x"0000",x"3b11",x"39d8"),
(x"3985",x"3d4c",x"36da",x"b796",x"bb0b",x"0000",x"3a44",x"3a25",x"3985",x"3d4c",x"3710",x"b817",x"badf",x"0000",x"3a4f",x"3a25",x"3994",x"3d47",x"3710",x"b458",x"bbb2",x"8000",x"3a4f",x"3a2c"),
(x"3752",x"3d7e",x"36da",x"3be0",x"31a3",x"8000",x"3a3d",x"3b53",x"3752",x"3d7e",x"3710",x"3bfd",x"aabe",x"0000",x"3a32",x"3b53",x"3754",x"3d80",x"3710",x"3afe",x"b7c4",x"0000",x"3a32",x"3b51"),
(x"36cb",x"3d56",x"36da",x"b86c",x"3aa9",x"0000",x"3a0c",x"3b12",x"36cb",x"3d56",x"3710",x"b922",x"3a22",x"0000",x"3a17",x"3b12",x"36c2",x"3d54",x"3710",x"bbe7",x"30ec",x"868d",x"3a17",x"3b14"),
(x"362c",x"3d73",x"36da",x"3550",x"3b8b",x"0000",x"3b06",x"39db",x"362c",x"3d73",x"3710",x"3609",x"3b68",x"8000",x"3b11",x"39db",x"35f7",x"3d7a",x"3710",x"3a6a",x"38c7",x"0000",x"3b11",x"39e6"),
(x"3972",x"3d50",x"36da",x"b0a0",x"bbea",x"0000",x"3a44",x"3a1d",x"3972",x"3d50",x"3710",x"b475",x"bbae",x"0000",x"3a4f",x"3a1d",x"3985",x"3d4c",x"3710",x"b817",x"badf",x"0000",x"3a4f",x"3a25"),
(x"392f",x"3d88",x"36da",x"b73b",x"3b22",x"8000",x"3bd5",x"39bf",x"392f",x"3d88",x"3710",x"b874",x"3aa4",x"0000",x"3bcb",x"39bf",x"3915",x"3d7a",x"3710",x"b845",x"3ac3",x"0000",x"3bcb",x"39b0"),
(x"3705",x"3d58",x"36da",x"b675",x"3b51",x"0000",x"3a0c",x"3b07",x"3705",x"3d58",x"3710",x"b599",x"3b7e",x"0000",x"3a17",x"3b07",x"36cb",x"3d56",x"3710",x"b922",x"3a22",x"0000",x"3a17",x"3b12"),
(x"35f7",x"3d7a",x"36da",x"3a05",x"3944",x"868d",x"3b06",x"39e6",x"35f7",x"3d7a",x"3710",x"3a6a",x"38c7",x"0000",x"3b11",x"39e6",x"35f1",x"3d7d",x"3710",x"3bf9",x"ad20",x"0000",x"3b11",x"39e8"),
(x"3963",x"3d51",x"36da",x"36c5",x"bb3f",x"0000",x"3a44",x"3a17",x"3963",x"3d51",x"3710",x"3420",x"bbba",x"0000",x"3a4f",x"3a17",x"3972",x"3d50",x"3710",x"b475",x"bbae",x"0000",x"3a4f",x"3a1d"),
(x"3754",x"3d80",x"36da",x"3ba5",x"b4b4",x"0000",x"3a3d",x"3b51",x"3754",x"3d80",x"3710",x"3afe",x"b7c4",x"0000",x"3a32",x"3b51",x"375f",x"3d83",x"3710",x"3bc1",x"b3d7",x"868d",x"3a32",x"3b4e"),
(x"3713",x"3d5a",x"36da",x"ba37",x"3909",x"0000",x"3a0c",x"3b04",x"3713",x"3d5a",x"3710",x"b972",x"39db",x"0000",x"3a17",x"3b04",x"3705",x"3d58",x"3710",x"b599",x"3b7e",x"0000",x"3a17",x"3b07"),
(x"35f1",x"3d7d",x"36da",x"3bcd",x"3318",x"0000",x"3b06",x"39e8",x"35f1",x"3d7d",x"3710",x"3bf9",x"ad20",x"0000",x"3b11",x"39e8",x"35f3",x"3d7e",x"3710",x"3b36",x"b6ea",x"8000",x"3b11",x"39e9"),
(x"395d",x"3d4f",x"36da",x"3ac1",x"b849",x"0000",x"3a44",x"3a15",x"395d",x"3d4f",x"3710",x"399d",x"b9b2",x"0000",x"3a4f",x"3a15",x"3963",x"3d51",x"3710",x"3420",x"bbba",x"0000",x"3a4f",x"3a17"),
(x"3915",x"3d7a",x"36da",x"b90a",x"3a36",x"0000",x"3bd5",x"39b0",x"3915",x"3d7a",x"3710",x"b845",x"3ac3",x"0000",x"3bcb",x"39b0",x"38f6",x"3d73",x"3710",x"b324",x"3bcc",x"0000",x"3bcb",x"39a3"),
(x"3716",x"3d5b",x"36da",x"bbad",x"b480",x"0000",x"3a0c",x"3b03",x"3716",x"3d5b",x"3710",x"bbb8",x"342d",x"0000",x"3a17",x"3b03",x"3713",x"3d5a",x"3710",x"b972",x"39db",x"0000",x"3a17",x"3b04"),
(x"35f3",x"3d7e",x"36da",x"3b84",x"b57a",x"0000",x"3b06",x"39e9",x"35f3",x"3d7e",x"3710",x"3b36",x"b6ea",x"8000",x"3b11",x"39e9",x"35fd",x"3d82",x"3710",x"3bf0",x"aff6",x"868d",x"3b11",x"39ed"),
(x"395a",x"3d4c",x"36da",x"3af1",x"b7f2",x"8000",x"3a44",x"3a12",x"395a",x"3d4c",x"3710",x"3b46",x"b6a7",x"8000",x"3a4f",x"3a12",x"395d",x"3d4f",x"3710",x"399d",x"b9b2",x"0000",x"3a4f",x"3a15"),
(x"38f6",x"3d73",x"36da",x"b551",x"3b8b",x"0000",x"3bd5",x"39a3",x"38f6",x"3d73",x"3710",x"b324",x"3bcc",x"0000",x"3bcb",x"39a3",x"38d5",x"3d71",x"3710",x"2dde",x"3bf7",x"0000",x"3bcb",x"3996"),
(x"3710",x"3d5d",x"36da",x"b80d",x"bae5",x"8000",x"3a18",x"3a1a",x"3710",x"3d5d",x"3710",x"b8f7",x"ba45",x"0000",x"3a23",x"3a1a",x"3716",x"3d5b",x"3710",x"bbb8",x"342d",x"0000",x"3a23",x"3a1b"),
(x"35fd",x"3d82",x"36da",x"3b91",x"b530",x"0000",x"3b06",x"39ed",x"35fd",x"3d82",x"3710",x"3bf0",x"aff6",x"868d",x"3b11",x"39ed",x"35fd",x"3d84",x"3710",x"3a08",x"3941",x"068d",x"3b11",x"39ee"),
(x"3953",x"3d47",x"36da",x"3857",x"bab8",x"8000",x"3a44",x"3a0e",x"3953",x"3d47",x"3710",x"39a8",x"b9a7",x"068d",x"3a4f",x"3a0e",x"395a",x"3d4c",x"3710",x"3b46",x"b6a7",x"8000",x"3a4f",x"3a12"),
(x"38d5",x"3d71",x"36da",x"1953",x"3c00",x"0000",x"3bd5",x"3996",x"38d5",x"3d71",x"3710",x"2dde",x"3bf7",x"0000",x"3bcb",x"3996",x"38bf",x"3d73",x"3710",x"35f3",x"3b6c",x"0000",x"3bcb",x"398d"),
(x"36f7",x"3d5e",x"36da",x"b05b",x"bbec",x"8000",x"3a18",x"3a15",x"36f7",x"3d5e",x"3710",x"b12d",x"bbe4",x"0000",x"3a23",x"3a15",x"3710",x"3d5d",x"3710",x"b8f7",x"ba45",x"0000",x"3a23",x"3a1a"),
(x"35fd",x"3d84",x"36da",x"3b87",x"3567",x"868d",x"3b06",x"39ee",x"35fd",x"3d84",x"3710",x"3a08",x"3941",x"068d",x"3b11",x"39ee",x"35f5",x"3d85",x"3710",x"32d5",x"3bd0",x"0000",x"3b11",x"39f0"),
(x"393f",x"3d45",x"36da",x"b2bb",x"bbd2",x"8000",x"3a44",x"3a06",x"393f",x"3d45",x"3710",x"1cea",x"bc00",x"8000",x"3a4f",x"3a06",x"3953",x"3d47",x"3710",x"39a8",x"b9a7",x"068d",x"3a4f",x"3a0e"),
(x"38bf",x"3d73",x"36da",x"3489",x"3bab",x"0000",x"3bd5",x"398d",x"38bf",x"3d73",x"3710",x"35f3",x"3b6c",x"0000",x"3bcb",x"398d",x"38b2",x"3d76",x"3710",x"3af2",x"37f0",x"0000",x"3bcb",x"3987"),
(x"362c",x"3d5d",x"36da",x"3609",x"bb68",x"0000",x"3a18",x"39ee",x"362c",x"3d5d",x"3710",x"3550",x"bb8b",x"0000",x"3a23",x"39ee",x"363b",x"3d5e",x"3710",x"3439",x"bbb7",x"868d",x"3a23",x"39f1"),
(x"35f5",x"3d85",x"36da",x"364b",x"3b5a",x"068d",x"3b06",x"39f0",x"35f5",x"3d85",x"3710",x"32d5",x"3bd0",x"0000",x"3b11",x"39f0",x"35e4",x"3d85",x"3710",x"b3c3",x"3bc2",x"0000",x"3b11",x"39f3"),
(x"392f",x"3d48",x"36da",x"b874",x"baa4",x"0000",x"3a44",x"39ff",x"392f",x"3d48",x"3710",x"b73b",x"bb22",x"0000",x"3a4f",x"39ff",x"393f",x"3d45",x"3710",x"1cea",x"bc00",x"8000",x"3a4f",x"3a06"),
(x"38b2",x"3d76",x"36da",x"3a0a",x"393e",x"8000",x"3bd5",x"3987",x"38b2",x"3d76",x"3710",x"3af2",x"37f0",x"0000",x"3bcb",x"3987",x"38b0",x"3d78",x"3710",x"3ba6",x"b4ac",x"0000",x"3bcb",x"3985"),
(x"363b",x"3d5e",x"36da",x"34bd",x"bba4",x"0000",x"3a18",x"39f1",x"363b",x"3d5e",x"3710",x"3439",x"bbb7",x"868d",x"3a23",x"39f1",x"36f7",x"3d5e",x"3710",x"b12d",x"bbe4",x"0000",x"3a23",x"3a15"),
(x"35e4",x"3d85",x"36da",x"b0fa",x"3be7",x"8000",x"3b06",x"39f3",x"35e4",x"3d85",x"3710",x"b3c3",x"3bc2",x"0000",x"3b11",x"39f3",x"35d3",x"3d83",x"3710",x"1c81",x"3c00",x"0000",x"3b11",x"39f7"),
(x"3754",x"3d4f",x"36da",x"3afe",x"37c4",x"0000",x"3a0c",x"3b41",x"3754",x"3d4f",x"3710",x"3ba5",x"34b5",x"0000",x"3a17",x"3b41",x"3752",x"3d51",x"3710",x"3be0",x"b1a3",x"868d",x"3a17",x"3b43"),
(x"38b0",x"3d78",x"36da",x"3bfc",x"2b27",x"0000",x"3bd5",x"3985",x"38b0",x"3d78",x"3710",x"3ba6",x"b4ac",x"0000",x"3bcb",x"3985",x"38b2",x"3d7a",x"3710",x"399c",x"b9b3",x"0000",x"3bcb",x"3983"),
(x"35f7",x"3d55",x"36da",x"3a6a",x"b8c7",x"0000",x"3a18",x"39e3",x"35f7",x"3d55",x"3710",x"3a05",x"b944",x"0000",x"3a23",x"39e3",x"362c",x"3d5d",x"3710",x"3550",x"bb8b",x"0000",x"3a23",x"39ee"),
(x"35d3",x"3d83",x"36da",x"b1d2",x"3bdd",x"0000",x"3b06",x"39f7",x"35d3",x"3d83",x"3710",x"1c81",x"3c00",x"0000",x"3b11",x"39f7",x"35bd",x"3d85",x"3710",x"afcb",x"3bf0",x"8000",x"3b11",x"39fb"),
(x"3915",x"3d55",x"36da",x"b845",x"bac3",x"0000",x"3a44",x"39f1",x"3915",x"3d55",x"3710",x"b90a",x"ba36",x"0000",x"3a4f",x"39f1",x"392f",x"3d48",x"3710",x"b73b",x"bb22",x"0000",x"3a4f",x"39ff"),
(x"38b2",x"3d7a",x"36da",x"3a58",x"b8de",x"0000",x"3a93",x"3ac5",x"38b2",x"3d7a",x"3710",x"399c",x"b9b3",x"0000",x"3a9e",x"3ac5",x"38bd",x"3d7d",x"3710",x"3456",x"bbb3",x"0000",x"3a9e",x"3ac9"),
(x"35f1",x"3d53",x"36da",x"3bf9",x"2d21",x"0000",x"3a18",x"39e1",x"35f1",x"3d53",x"3710",x"3bcd",x"b318",x"0000",x"3a23",x"39e1",x"35f7",x"3d55",x"3710",x"3a05",x"b944",x"0000",x"3a23",x"39e3"),
(x"35bd",x"3d85",x"36da",x"2c75",x"3bfb",x"868d",x"3b06",x"39fb",x"35bd",x"3d85",x"3710",x"afcb",x"3bf0",x"8000",x"3b11",x"39fb",x"359e",x"3d82",x"3710",x"b925",x"3a1f",x"0000",x"3b11",x"3a01"),
(x"375f",x"3d4c",x"36da",x"3bc1",x"33d7",x"068d",x"3a0c",x"3b3e",x"375f",x"3d4c",x"3710",x"3b14",x"3774",x"8000",x"3a17",x"3b3e",x"3754",x"3d4f",x"3710",x"3ba5",x"34b5",x"0000",x"3a17",x"3b41"),
(x"38bd",x"3d7d",x"36da",x"35fc",x"bb6b",x"0000",x"3a93",x"3ac9",x"38bd",x"3d7d",x"3710",x"3456",x"bbb3",x"0000",x"3a9e",x"3ac9",x"38c9",x"3d7e",x"3710",x"34cb",x"bba1",x"0000",x"3a9e",x"3ace"),
(x"35f3",x"3d51",x"36da",x"3b36",x"36ea",x"8000",x"3a18",x"39e0",x"35f3",x"3d51",x"3710",x"3b84",x"357a",x"0000",x"3a23",x"39e0",x"35f1",x"3d53",x"3710",x"3bcd",x"b318",x"0000",x"3a23",x"39e1"),
(x"359e",x"3d82",x"36da",x"b80b",x"3ae7",x"8000",x"3b06",x"3a01",x"359e",x"3d82",x"3710",x"b925",x"3a1f",x"0000",x"3b11",x"3a01",x"358a",x"3d7c",x"3710",x"bbad",x"3481",x"068d",x"3b11",x"3a07"),
(x"38f6",x"3d5d",x"36da",x"b324",x"bbcc",x"0000",x"3a44",x"39e4",x"38f6",x"3d5d",x"3710",x"b551",x"bb8b",x"0000",x"3a4f",x"39e4",x"3915",x"3d55",x"3710",x"b90a",x"ba36",x"0000",x"3a4f",x"39f1"),
(x"38c9",x"3d7e",x"36da",x"3385",x"bbc6",x"0000",x"3a93",x"3ace",x"38c9",x"3d7e",x"3710",x"34cb",x"bba1",x"0000",x"3a9e",x"3ace",x"38d4",x"3d80",x"3710",x"38a8",x"ba80",x"8000",x"3a9e",x"3ad2"),
(x"35fd",x"3d4e",x"36da",x"3bf0",x"2ff4",x"8000",x"3a18",x"39dc",x"35fd",x"3d4e",x"3710",x"3b91",x"3530",x"8000",x"3a23",x"39dc",x"35f3",x"3d51",x"3710",x"3b84",x"357a",x"0000",x"3a23",x"39e0"),
(x"358a",x"3d7c",x"36da",x"bb1e",x"374c",x"8000",x"3b06",x"3a07",x"358a",x"3d7c",x"3710",x"bbad",x"3481",x"068d",x"3b11",x"3a07",x"3587",x"3d77",x"3710",x"bb8b",x"b553",x"0000",x"3b11",x"3a0b"),
(x"38d5",x"3d5f",x"36da",x"2dde",x"bbf7",x"0000",x"3a44",x"39d8",x"38d5",x"3d5f",x"3710",x"1987",x"bc00",x"0000",x"3a4f",x"39d8",x"38f6",x"3d5d",x"3710",x"b551",x"bb8b",x"0000",x"3a4f",x"39e4"),
(x"38d4",x"3d80",x"36da",x"37f2",x"baf1",x"8000",x"3a93",x"3ad2",x"38d4",x"3d80",x"3710",x"38a8",x"ba80",x"8000",x"3a9e",x"3ad2",x"38d9",x"3d82",x"3710",x"3bfc",x"ab00",x"0000",x"3a9e",x"3ad5"),
(x"3a26",x"3d45",x"36da",x"3bff",x"26b5",x"0000",x"3a38",x"33fa",x"3a26",x"3d45",x"3710",x"3bcf",x"2680",x"32dc",x"3a36",x"33ca",x"3a25",x"3d5c",x"3710",x"3bd6",x"2604",x"3256",x"3a49",x"33c0"),
(x"35fd",x"3d4c",x"36da",x"3a08",x"b941",x"8000",x"3a18",x"39db",x"35fd",x"3d4c",x"3710",x"3b87",x"b567",x"868d",x"3a23",x"39db",x"35fd",x"3d4e",x"3710",x"3b91",x"3530",x"8000",x"3a23",x"39dc"),
(x"3587",x"3d77",x"36da",x"bbf7",x"adba",x"8000",x"3b06",x"3a0b",x"3587",x"3d77",x"3710",x"bb8b",x"b553",x"0000",x"3b11",x"3a0b",x"3593",x"3d72",x"3710",x"bc00",x"15bc",x"0000",x"3b11",x"3a0f"),
(x"38bf",x"3d5d",x"36da",x"35f3",x"bb6c",x"0000",x"3a44",x"39cf",x"38bf",x"3d5d",x"3710",x"3489",x"bbab",x"0000",x"3a4f",x"39cf",x"38d5",x"3d5f",x"3710",x"1987",x"bc00",x"0000",x"3a4f",x"39d8"),
(x"38d9",x"3d82",x"36da",x"3b88",x"b564",x"0000",x"3a93",x"3ad5",x"38d9",x"3d82",x"3710",x"3bfc",x"ab00",x"0000",x"3a9e",x"3ad5",x"38d8",x"3d84",x"3710",x"3b96",x"350f",x"0000",x"3a9e",x"3ad6"),
(x"35f5",x"3d4b",x"36da",x"32d5",x"bbd0",x"0000",x"3a18",x"39d9",x"35f5",x"3d4b",x"3710",x"364b",x"bb5a",x"0000",x"3a23",x"39d9",x"35fd",x"3d4c",x"3710",x"3b87",x"b567",x"868d",x"3a23",x"39db"),
(x"3593",x"3d72",x"36da",x"bbda",x"b21b",x"0000",x"3b06",x"3a0f",x"3593",x"3d72",x"3710",x"bc00",x"15bc",x"0000",x"3b11",x"3a0f",x"3592",x"3d70",x"3710",x"ba08",x"3941",x"0000",x"3b11",x"3a11"),
(x"38b2",x"3d5a",x"36da",x"3af2",x"b7f0",x"0000",x"3a44",x"39ca",x"38b2",x"3d5a",x"3710",x"3a0a",x"b93f",x"0000",x"3a4f",x"39ca",x"38bf",x"3d5d",x"3710",x"3489",x"bbab",x"0000",x"3a4f",x"39cf"),
(x"38d8",x"3d84",x"36da",x"3be4",x"312f",x"8000",x"3a93",x"3ad6",x"38d8",x"3d84",x"3710",x"3b96",x"350f",x"0000",x"3a9e",x"3ad6",x"38c7",x"3d87",x"3710",x"364a",x"3b5a",x"0000",x"3a9e",x"3add"),
(x"35e4",x"3d4b",x"36da",x"b3c3",x"bbc2",x"0000",x"3a18",x"39d6",x"35e4",x"3d4b",x"3710",x"b0fa",x"bbe7",x"8000",x"3a23",x"39d6",x"35f5",x"3d4b",x"3710",x"364b",x"bb5a",x"0000",x"3a23",x"39d9"),
(x"3592",x"3d70",x"36da",x"bba4",x"34bb",x"0000",x"3a5f",x"3b35",x"3592",x"3d70",x"3710",x"ba08",x"3941",x"0000",x"3a6a",x"3b35",x"357d",x"3d70",x"3710",x"26bb",x"3bff",x"0000",x"3a6a",x"3b39"),
(x"38b0",x"3d57",x"36da",x"3ba6",x"34ab",x"0000",x"3a33",x"3a17",x"38b0",x"3d57",x"3710",x"3bfc",x"ab2b",x"0000",x"3a3e",x"3a17",x"38b2",x"3d5a",x"3710",x"3a0a",x"b93f",x"0000",x"3a3e",x"3a19"),
(x"38c7",x"3d87",x"36da",x"3654",x"3b58",x"8000",x"3a93",x"3add",x"38c7",x"3d87",x"3710",x"364a",x"3b5a",x"0000",x"3a9e",x"3add",x"38b7",x"3d8b",x"3710",x"32f6",x"3bce",x"0000",x"3a9e",x"3ae4"),
(x"35d3",x"3d4c",x"36da",x"1c81",x"bc00",x"0000",x"3a18",x"39d2",x"35d3",x"3d4c",x"3710",x"b1d2",x"bbdd",x"0000",x"3a23",x"39d2",x"35e4",x"3d4b",x"3710",x"b0fa",x"bbe7",x"8000",x"3a23",x"39d6"),
(x"357d",x"3d70",x"36da",x"a8c9",x"3bfe",x"0000",x"3a5f",x"3b39",x"357d",x"3d70",x"3710",x"26bb",x"3bff",x"0000",x"3a6a",x"3b39",x"3555",x"3d71",x"3710",x"35eb",x"3b6e",x"0000",x"3a6a",x"3b40"),
(x"38b2",x"3d55",x"36da",x"399c",x"39b3",x"8000",x"3a33",x"3a15",x"38b2",x"3d55",x"3710",x"3a58",x"38de",x"0000",x"3a3e",x"3a15",x"38b0",x"3d57",x"3710",x"3bfc",x"ab2b",x"0000",x"3a3e",x"3a17"),
(x"38b7",x"3d8b",x"36da",x"3528",x"3b92",x"8000",x"3a93",x"3ae4",x"38b7",x"3d8b",x"3710",x"32f6",x"3bce",x"0000",x"3a9e",x"3ae4",x"3894",x"3d8c",x"3710",x"b036",x"3bee",x"0000",x"3a9e",x"3af1"),
(x"35bd",x"3d4b",x"36da",x"afc9",x"bbf0",x"8000",x"3a18",x"39ce",x"35bd",x"3d4b",x"3710",x"2c74",x"bbfb",x"068d",x"3a23",x"39ce",x"35d3",x"3d4c",x"3710",x"b1d2",x"bbdd",x"0000",x"3a23",x"39d2"),
(x"3555",x"3d71",x"36da",x"345a",x"3bb2",x"0000",x"3a5f",x"3b40",x"3555",x"3d71",x"3710",x"35eb",x"3b6e",x"0000",x"3a6a",x"3b40",x"353f",x"3d74",x"3710",x"379f",x"3b08",x"0000",x"3a6a",x"3b45"),
(x"38bd",x"3d52",x"36da",x"3456",x"3bb3",x"0000",x"3a33",x"3a11",x"38bd",x"3d52",x"3710",x"35fc",x"3b6b",x"0000",x"3a3e",x"3a11",x"38b2",x"3d55",x"3710",x"3a58",x"38de",x"0000",x"3a3e",x"3a15"),
(x"3894",x"3d8c",x"36da",x"aa0a",x"3bfd",x"8000",x"3a93",x"3af1",x"3894",x"3d8c",x"3710",x"b036",x"3bee",x"0000",x"3a9e",x"3af1",x"3877",x"3d89",x"3710",x"b8aa",x"3a7f",x"8000",x"3a9e",x"3afc"),
(x"359e",x"3d4e",x"36da",x"b925",x"ba1f",x"8000",x"3a18",x"39c8",x"359e",x"3d4e",x"3710",x"b80b",x"bae7",x"0000",x"3a23",x"39c8",x"35bd",x"3d4b",x"3710",x"2c74",x"bbfb",x"068d",x"3a23",x"39ce"),
(x"353f",x"3d74",x"36da",x"3746",x"3b1f",x"0000",x"3a5f",x"3b45",x"353f",x"3d74",x"3710",x"379f",x"3b08",x"0000",x"3a6a",x"3b45",x"351b",x"3d79",x"3710",x"350e",x"3b96",x"0000",x"3a6a",x"3b4d"),
(x"38c9",x"3d51",x"36da",x"34cb",x"3ba1",x"8000",x"3a33",x"3a0c",x"38c9",x"3d51",x"3710",x"3385",x"3bc6",x"0000",x"3a3e",x"3a0c",x"38bd",x"3d52",x"3710",x"35fc",x"3b6b",x"0000",x"3a3e",x"3a11"),
(x"3877",x"3d89",x"36da",x"b74e",x"3b1d",x"0000",x"3a93",x"3afc",x"3877",x"3d89",x"3710",x"b8aa",x"3a7f",x"8000",x"3a9e",x"3afc",x"386d",x"3d84",x"3710",x"bba8",x"34a3",x"0000",x"3a9e",x"3b01"),
(x"358a",x"3d54",x"36da",x"bbad",x"b481",x"8000",x"3a18",x"39c2",x"358a",x"3d54",x"3710",x"bb1e",x"b74c",x"0000",x"3a23",x"39c2",x"359e",x"3d4e",x"3710",x"b80b",x"bae7",x"0000",x"3a23",x"39c8"),
(x"351b",x"3d79",x"36da",x"3664",x"3b55",x"0000",x"3a5f",x"3b4d",x"351b",x"3d79",x"3710",x"350e",x"3b96",x"0000",x"3a6a",x"3b4d",x"3501",x"3d7b",x"3710",x"ada6",x"3bf8",x"0000",x"3a6a",x"3b52"),
(x"38d4",x"3d4f",x"36da",x"38a8",x"3a80",x"8000",x"3a33",x"3a08",x"38d4",x"3d4f",x"3710",x"37f2",x"3af1",x"8000",x"3a3e",x"3a08",x"38c9",x"3d51",x"3710",x"3385",x"3bc6",x"0000",x"3a3e",x"3a0c"),
(x"386d",x"3d84",x"36da",x"bac4",x"3844",x"8000",x"3a93",x"3b01",x"386d",x"3d84",x"3710",x"bba8",x"34a3",x"0000",x"3a9e",x"3b01",x"386c",x"3d7f",x"3710",x"bb38",x"b6e2",x"868d",x"3a9e",x"3b05"),
(x"3587",x"3d59",x"36da",x"bb8b",x"3553",x"0000",x"3a18",x"39be",x"3587",x"3d59",x"3710",x"bbf7",x"2dba",x"0000",x"3a23",x"39be",x"358a",x"3d54",x"3710",x"bb1e",x"b74c",x"0000",x"3a23",x"39c2"),
(x"3501",x"3d7b",x"36da",x"2d0c",x"3bf9",x"8000",x"3a5f",x"3b52",x"3501",x"3d7b",x"3710",x"ada6",x"3bf8",x"0000",x"3a6a",x"3b52",x"34e9",x"3d79",x"3710",x"b698",x"3b49",x"0000",x"3a6a",x"3b57"),
(x"38d9",x"3d4d",x"36da",x"3bfc",x"2b00",x"8000",x"3a33",x"3a06",x"38d9",x"3d4d",x"3710",x"3b88",x"3564",x"0000",x"3a3e",x"3a06",x"38d4",x"3d4f",x"3710",x"37f2",x"3af1",x"8000",x"3a3e",x"3a08"),
(x"386c",x"3d7f",x"36da",x"bbdd",x"b1e1",x"8000",x"3a93",x"3b05",x"386c",x"3d7f",x"3710",x"bb38",x"b6e2",x"868d",x"3a9e",x"3b05",x"3872",x"3d7b",x"3710",x"b902",x"ba3c",x"0000",x"3a9e",x"3b08"),
(x"3593",x"3d5d",x"36da",x"bc00",x"95bc",x"0000",x"3a18",x"39ba",x"3593",x"3d5d",x"3710",x"bbda",x"321b",x"8000",x"3a23",x"39ba",x"3587",x"3d59",x"3710",x"bbf7",x"2dba",x"0000",x"3a23",x"39be"),
(x"34e9",x"3d79",x"36da",x"b50d",x"3b97",x"8000",x"3a5f",x"3b57",x"34e9",x"3d79",x"3710",x"b698",x"3b49",x"0000",x"3a6a",x"3b57",x"34cb",x"3d75",x"3710",x"b501",x"3b99",x"0000",x"3a6a",x"3b5d"),
(x"38d8",x"3d4c",x"36da",x"3b96",x"b50f",x"0000",x"3a33",x"3a05",x"38d8",x"3d4c",x"3710",x"3be4",x"b12f",x"8a8d",x"3a3e",x"3a05",x"38d9",x"3d4d",x"3710",x"3b88",x"3564",x"0000",x"3a3e",x"3a06"),
(x"3872",x"3d7b",x"36da",x"b9d1",x"b97d",x"8000",x"3a93",x"3b08",x"3872",x"3d7b",x"3710",x"b902",x"ba3c",x"0000",x"3a9e",x"3b08",x"3885",x"3d77",x"3710",x"b83d",x"bac8",x"0000",x"3a9e",x"3b10"),
(x"3592",x"3d60",x"36da",x"ba08",x"b941",x"8000",x"3a18",x"39b8",x"3592",x"3d60",x"3710",x"bba4",x"b4bb",x"0000",x"3a23",x"39b8",x"3593",x"3d5d",x"3710",x"bbda",x"321b",x"8000",x"3a23",x"39ba"),
(x"34cb",x"3d75",x"36da",x"b64c",x"3b5a",x"0000",x"3a5f",x"3b5d",x"34cb",x"3d75",x"3710",x"b501",x"3b99",x"0000",x"3a6a",x"3b5d",x"34bb",x"3d73",x"3710",x"b13f",x"3be4",x"0000",x"3a6a",x"3b60"),
(x"38c7",x"3d48",x"36da",x"364a",x"bb5b",x"8000",x"3a33",x"39fd",x"38c7",x"3d48",x"3710",x"3653",x"bb59",x"0000",x"3a3e",x"39fd",x"38d8",x"3d4c",x"3710",x"3be4",x"b12f",x"8a8d",x"3a3e",x"3a05"),
(x"3885",x"3d77",x"36da",x"b7eb",x"baf3",x"0000",x"3a93",x"3b10",x"3885",x"3d77",x"3710",x"b83d",x"bac8",x"0000",x"3a9e",x"3b10",x"388c",x"3d75",x"3710",x"bbfd",x"a9ab",x"0000",x"3a9e",x"3b13"),
(x"357d",x"3d60",x"36da",x"26c8",x"bbff",x"0000",x"3a5f",x"3bad",x"357d",x"3d60",x"3710",x"a8c9",x"bbfe",x"0000",x"3a6a",x"3bad",x"3592",x"3d60",x"3710",x"bba4",x"b4bb",x"0000",x"3a6a",x"3bb1"),
(x"34bb",x"3d73",x"36da",x"b31c",x"3bcc",x"0000",x"3a5f",x"3b60",x"34bb",x"3d73",x"3710",x"b13f",x"3be4",x"0000",x"3a6a",x"3b60",x"349b",x"3d73",x"3710",x"b4a8",x"3ba7",x"0000",x"3a6a",x"3b66"),
(x"38b7",x"3d45",x"36da",x"32f6",x"bbce",x"0000",x"3a33",x"39f7",x"38b7",x"3d45",x"3710",x"3528",x"bb92",x"0000",x"3a3e",x"39f7",x"38c7",x"3d48",x"3710",x"3653",x"bb59",x"0000",x"3a3e",x"39fd"),
(x"388c",x"3d75",x"36da",x"bb54",x"b669",x"8000",x"3a3d",x"3bb1",x"388c",x"3d75",x"3710",x"bbfd",x"a9ab",x"0000",x"3a32",x"3bb1",x"388c",x"3d73",x"3710",x"b967",x"39e6",x"0000",x"3a32",x"3bb0"),
(x"3555",x"3d5f",x"36da",x"35eb",x"bb6e",x"0000",x"3a5f",x"3ba5",x"3555",x"3d5f",x"3710",x"345a",x"bbb2",x"0000",x"3a6a",x"3ba5",x"357d",x"3d60",x"3710",x"a8c9",x"bbfe",x"0000",x"3a6a",x"3bad"),
(x"349b",x"3d73",x"36da",x"b221",x"3bda",x"0000",x"3a5f",x"3b66",x"349b",x"3d73",x"3710",x"b4a8",x"3ba7",x"0000",x"3a6a",x"3b66",x"3485",x"3d71",x"3710",x"b92c",x"3a1a",x"0000",x"3a6a",x"3b6b"),
(x"3894",x"3d44",x"36da",x"b036",x"bbee",x"0000",x"3a33",x"39ea",x"3894",x"3d44",x"3710",x"aa0a",x"bbfd",x"8000",x"3a3e",x"39ea",x"38b7",x"3d45",x"3710",x"3528",x"bb92",x"0000",x"3a3e",x"39f7"),
(x"388c",x"3d73",x"36da",x"bb52",x"3671",x"0000",x"3a3d",x"3bb0",x"388c",x"3d73",x"3710",x"b967",x"39e6",x"0000",x"3a32",x"3bb0",x"3885",x"3d72",x"3710",x"b25f",x"3bd7",x"8000",x"3a32",x"3bad"),
(x"353f",x"3d5c",x"36da",x"379f",x"bb08",x"0000",x"3a5f",x"3ba1",x"353f",x"3d5c",x"3710",x"3746",x"bb1f",x"0000",x"3a6a",x"3ba1",x"3555",x"3d5f",x"3710",x"345a",x"bbb2",x"0000",x"3a6a",x"3ba5"),
(x"3485",x"3d71",x"36da",x"b819",x"3ade",x"8000",x"3a5f",x"3b6b",x"3485",x"3d71",x"3710",x"b92c",x"3a1a",x"0000",x"3a6a",x"3b6b",x"3475",x"3d6c",x"3710",x"bbab",x"348e",x"8000",x"3a6a",x"3b70"),
(x"3877",x"3d47",x"36da",x"b8aa",x"ba7f",x"8000",x"3a33",x"39de",x"3877",x"3d47",x"3710",x"b74e",x"bb1d",x"8000",x"3a3e",x"39de",x"3894",x"3d44",x"3710",x"aa0a",x"bbfd",x"8000",x"3a3e",x"39ea"),
(x"3760",x"3d86",x"36da",x"3bfa",x"2cac",x"8000",x"3a3d",x"3b4c",x"3760",x"3d86",x"3710",x"3b92",x"3528",x"8000",x"3a32",x"3b4c",x"3753",x"3d89",x"3710",x"37e4",x"3af5",x"8000",x"3a32",x"3b48"),
(x"3a2d",x"3d5e",x"36da",x"3bfe",x"a8f0",x"0000",x"3bea",x"3999",x"3a2d",x"3d5e",x"3710",x"3bde",x"a849",x"31a9",x"3beb",x"398f",x"3a2f",x"3d73",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"398f"),
(x"351b",x"3d57",x"36da",x"350e",x"bb96",x"0000",x"3a5f",x"3b99",x"351b",x"3d57",x"3710",x"3664",x"bb55",x"0000",x"3a6a",x"3b99",x"353f",x"3d5c",x"3710",x"3746",x"bb1f",x"0000",x"3a6a",x"3ba1"),
(x"3a27",x"3d8b",x"36da",x"a3ae",x"3bff",x"0000",x"3bd5",x"3a28",x"3a27",x"3d8b",x"3710",x"a3ef",x"3bff",x"9818",x"3bcb",x"3a28",x"39f5",x"3d8a",x"3710",x"a4e3",x"3bff",x"1818",x"3bcb",x"3a14"),
(x"386d",x"3d4b",x"36da",x"bba8",x"b4a3",x"868d",x"3a33",x"39d9",x"386d",x"3d4b",x"3710",x"bac4",x"b844",x"0000",x"3a3e",x"39d9",x"3877",x"3d47",x"3710",x"b74e",x"bb1d",x"8000",x"3a3e",x"39de"),
(x"3885",x"3d72",x"36da",x"b304",x"3bce",x"0000",x"3a3d",x"3bad",x"3885",x"3d72",x"3710",x"b25f",x"3bd7",x"8000",x"3a32",x"3bad",x"382a",x"3d72",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b89"),
(x"3501",x"3d55",x"36da",x"ada8",x"bbf8",x"8000",x"3a5f",x"3b94",x"3501",x"3d55",x"3710",x"2d0c",x"bbf9",x"0000",x"3a6a",x"3b94",x"351b",x"3d57",x"3710",x"3664",x"bb55",x"0000",x"3a6a",x"3b99"),
(x"386c",x"3d51",x"36da",x"bb38",x"36e2",x"068d",x"3a33",x"39d5",x"386c",x"3d51",x"3710",x"bbdd",x"31e1",x"0000",x"3a3e",x"39d5",x"386d",x"3d4b",x"3710",x"bac4",x"b844",x"0000",x"3a3e",x"39d9"),
(x"382a",x"3d72",x"36da",x"2f40",x"3bf2",x"8000",x"3a3d",x"3b89",x"382a",x"3d72",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b89",x"3813",x"3d74",x"3710",x"a8bf",x"3bfe",x"8000",x"3a32",x"3b80"),
(x"3a25",x"3d5c",x"36da",x"367a",x"bb50",x"0000",x"3bc3",x"39b4",x"3a25",x"3d5c",x"3710",x"3700",x"bb23",x"2f05",x"3bbd",x"39bd",x"3a2d",x"3d5e",x"3710",x"3644",x"bb4c",x"2f83",x"3bba",x"39ba"),
(x"3a1f",x"4041",x"3733",x"3b23",x"251e",x"3738",x"39c4",x"339f",x"3a25",x"4041",x"3710",x"3bd6",x"2604",x"3256",x"39c5",x"33c0",x"3a20",x"4036",x"3732",x"3b18",x"2439",x"3763",x"39b1",x"33aa"),
(x"3a18",x"4041",x"3748",x"36c9",x"29dc",x"3b3c",x"39c4",x"3388",x"3a1f",x"4041",x"3733",x"3b23",x"251e",x"3738",x"39c4",x"339f",x"3a19",x"4036",x"3749",x"3871",x"2587",x"3aa6",x"39b0",x"3392"),
(x"3a10",x"4041",x"3749",x"b4de",x"2b76",x"3b9b",x"39c3",x"337b",x"3a18",x"4041",x"3748",x"36c9",x"29dc",x"3b3c",x"39c4",x"3388",x"3a14",x"4036",x"374e",x"2fa2",x"2997",x"3bef",x"39b0",x"3387"),
(x"3a09",x"4041",x"373b",x"b9d7",x"2404",x"3976",x"39c3",x"3369",x"3a10",x"4041",x"3749",x"b4de",x"2b76",x"3b9b",x"39c3",x"337b",x"3a0d",x"4036",x"374b",x"b745",x"2966",x"3b1e",x"39b0",x"337b"),
(x"3a09",x"4042",x"373a",x"baf6",x"2b34",x"37d2",x"3b1b",x"3899",x"3a09",x"4041",x"373b",x"b7a6",x"3a67",x"35ca",x"3b1c",x"3899",x"3a03",x"4042",x"370e",x"ae5c",x"3b3a",x"36a9",x"3b1f",x"38a1"),
(x"3a09",x"4041",x"373b",x"b7a6",x"3a67",x"35ca",x"3b1c",x"3899",x"3a09",x"4042",x"373a",x"baf6",x"2b34",x"37d2",x"3b1b",x"3899",x"3a10",x"4041",x"3749",x"b3ab",x"a4bc",x"3bc3",x"3b1a",x"3895"),
(x"3a08",x"404d",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"39a7",x"3a09",x"4042",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"39a8",x"3a04",x"404d",x"3727",x"bbc5",x"a901",x"3377",x"3bfb",x"39a3"),
(x"3a03",x"4042",x"370e",x"bbc2",x"ab4f",x"338c",x"3bea",x"399f",x"3a04",x"404d",x"3727",x"bbc5",x"a901",x"3377",x"3bfb",x"39a3",x"3a09",x"4042",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"39a8"),
(x"3a09",x"4042",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"39a8",x"3a08",x"404d",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"39a7",x"3a11",x"4042",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"39ac"),
(x"3a11",x"4042",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"39ac",x"3a0f",x"404d",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"39ab",x"3a19",x"4043",x"374d",x"3400",x"aa73",x"3bbc",x"3bec",x"39af"),
(x"3a17",x"404d",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3bfc",x"39af",x"3a1d",x"404d",x"374d",x"3802",x"a90b",x"3aea",x"3bfc",x"39b1",x"3a19",x"4043",x"374d",x"3400",x"aa73",x"3bbc",x"3bec",x"39af"),
(x"3a1d",x"404d",x"374d",x"3802",x"a90b",x"3aea",x"3bfc",x"39b1",x"3a24",x"404d",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"39b5",x"3a21",x"4043",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"39b3"),
(x"3a24",x"404d",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"39b5",x"3a2a",x"404d",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"39ba",x"3a25",x"4043",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"39b6"),
(x"3a1f",x"4041",x"3733",x"37fe",x"ba99",x"3438",x"3b19",x"388d",x"3a25",x"4043",x"3738",x"36f3",x"bae7",x"3422",x"3b16",x"388d",x"3a25",x"4041",x"3710",x"3700",x"bb23",x"2f05",x"3b1b",x"3887"),
(x"3a02",x"4036",x"3724",x"bb1f",x"1a24",x"3747",x"39b0",x"3352",x"3a09",x"4041",x"373b",x"b9d7",x"2404",x"3976",x"39c3",x"3369",x"3a07",x"4036",x"373c",x"bac4",x"2853",x"3841",x"39b0",x"336a"),
(x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e",x"3a09",x"4041",x"373b",x"b9d7",x"2404",x"3976",x"39c3",x"3369",x"3a02",x"4036",x"3724",x"bb1f",x"1a24",x"3747",x"39b0",x"3352"),
(x"3a10",x"4041",x"3749",x"b3ab",x"a4bc",x"3bc3",x"3b1a",x"3895",x"3a11",x"4042",x"374a",x"b548",x"b37f",x"3b50",x"3b18",x"3896",x"3a18",x"4041",x"3748",x"2918",x"b8de",x"3a57",x"3b18",x"3893"),
(x"3a1f",x"4041",x"3733",x"37fe",x"ba99",x"3438",x"3b19",x"388d",x"3a18",x"4041",x"3748",x"2918",x"b8de",x"3a57",x"3b18",x"3893",x"3a21",x"4043",x"3744",x"37e0",x"ba17",x"36be",x"3b16",x"388f"),
(x"3a2f",x"404d",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"381d",x"3a2a",x"404d",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3821",x"3a26",x"404d",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3820"),
(x"3a2a",x"404d",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3821",x"3a24",x"404d",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3826",x"3a20",x"404d",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3827"),
(x"3a24",x"404d",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3826",x"3a1d",x"404d",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"382a",x"3a1a",x"404d",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"382b"),
(x"3a17",x"404d",x"3751",x"2fd8",x"39a6",x"3994",x"3b24",x"382d",x"3a0f",x"404d",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3830",x"3a15",x"404d",x"374b",x"aaab",x"39a6",x"39a5",x"3b22",x"382d"),
(x"3a0f",x"404d",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3830",x"3a08",x"404d",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3832",x"3a0f",x"404e",x"3749",x"b6e3",x"3561",x"3ab3",x"3b21",x"382f"),
(x"3a08",x"404d",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3832",x"3a04",x"404d",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3835",x"3a09",x"404e",x"373e",x"ba28",x"9df0",x"391a",x"3b1e",x"3831"),
(x"39fb",x"404d",x"3713",x"a9a8",x"a460",x"3bfd",x"39d7",x"333d",x"3a02",x"404d",x"3711",x"315a",x"2bae",x"3bdf",x"39d6",x"3349",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e"),
(x"3a20",x"404d",x"3739",x"3abd",x"a8b5",x"384c",x"39d7",x"339e",x"3a24",x"4059",x"372b",x"3b86",x"a8a8",x"3564",x"39eb",x"33b1",x"3a26",x"404d",x"3710",x"3bed",x"a7ae",x"3024",x"39d7",x"33c4"),
(x"3a21",x"4059",x"373a",x"3acd",x"a5ae",x"3834",x"39eb",x"33a3",x"3a20",x"404d",x"3739",x"3abd",x"a8b5",x"384c",x"39d7",x"339e",x"3a1a",x"4059",x"3749",x"38cd",x"a812",x"3a64",x"39eb",x"3391"),
(x"3a1a",x"404d",x"3746",x"38a5",x"a839",x"3a81",x"39d8",x"338e",x"3a15",x"404d",x"374b",x"2e57",x"a8d3",x"3bf4",x"39d8",x"3385",x"3a1a",x"4059",x"3749",x"38cd",x"a812",x"3a64",x"39eb",x"3391"),
(x"3a15",x"404d",x"374b",x"2e57",x"a8d3",x"3bf4",x"39d8",x"3385",x"3a0f",x"404e",x"3749",x"b771",x"a91b",x"3b13",x"39d8",x"3379",x"3a14",x"4059",x"374f",x"32be",x"a89e",x"3bd0",x"39eb",x"3384"),
(x"3a0f",x"404e",x"3749",x"b771",x"a91b",x"3b13",x"39d8",x"3379",x"3a09",x"404e",x"373e",x"ba21",x"a786",x"3921",x"39d8",x"336a",x"3a0d",x"4059",x"374b",x"b6cb",x"a758",x"3b3d",x"39eb",x"3378"),
(x"3a07",x"4059",x"373c",x"baa0",x"a6bb",x"3879",x"39eb",x"3366",x"3a09",x"404e",x"373e",x"ba21",x"a786",x"3921",x"39d8",x"336a",x"3a00",x"4059",x"3722",x"ba6c",x"a860",x"38c2",x"39ea",x"334c"),
(x"3a00",x"4059",x"3722",x"ba6c",x"a860",x"38c2",x"39ea",x"334c",x"3a01",x"404d",x"371c",x"b9f4",x"a495",x"3957",x"39d7",x"334a",x"39fc",x"4059",x"3718",x"b8fc",x"a86a",x"3a40",x"39eb",x"3340"),
(x"3475",x"4045",x"3710",x"0000",x"0000",x"3c00",x"39c9",x"2450",x"3475",x"404a",x"3710",x"0000",x"0000",x"3c00",x"39d1",x"2450",x"3485",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"24c1"),
(x"349b",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"255f",x"3485",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"24c1",x"349b",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"255f"),
(x"34bb",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2642",x"349b",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"255f",x"34bb",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2642"),
(x"34bb",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2642",x"34bb",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2642",x"34cb",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"26b3"),
(x"34e9",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39be",x"278b",x"34cb",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"26b3",x"34e9",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"278b"),
(x"34e9",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39be",x"278b",x"34e9",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"278b",x"3501",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"281a"),
(x"3501",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"281a",x"3501",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"281a",x"351b",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39be",x"2878"),
(x"351b",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39be",x"2878",x"351b",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dc",x"2878",x"353f",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"28fa"),
(x"3555",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2949",x"353f",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"28fa",x"3555",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2949"),
(x"3555",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2949",x"3555",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2949",x"357d",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"29d7"),
(x"357d",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"29d7",x"357d",x"404b",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"29d7",x"3592",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2a20"),
(x"36f7",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2d8d",x"36f7",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2d8d",x"363b",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2c3f"),
(x"362c",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2c23",x"363b",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2c3f",x"362c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2c23"),
(x"362c",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2c23",x"362c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2c23",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b"),
(x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b",x"3592",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d4",x"2a20"),
(x"35e4",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2b47",x"35f5",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2b83",x"35fd",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2ba0"),
(x"35d3",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"2b0a",x"35e4",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2b47",x"35f3",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2b7d"),
(x"35bd",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2ab9",x"35d3",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"2b0a",x"35f1",x"4052",x"3710",x"0000",x"0000",x"3c00",x"39df",x"2b76"),
(x"35fd",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"2ba0",x"35f5",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2b83",x"35fd",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2ba0"),
(x"35fd",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2ba0",x"35e4",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2b47",x"35f3",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2b7d"),
(x"35f3",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2b7d",x"35d3",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2b0a",x"35f1",x"403d",x"3710",x"868d",x"8cea",x"3c00",x"39bb",x"2b76"),
(x"35f1",x"403d",x"3710",x"868d",x"8cea",x"3c00",x"39bb",x"2b76",x"35bd",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"2ab9",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b"),
(x"359e",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2a4d",x"35bd",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2ab9",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b"),
(x"3587",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"29fa",x"358a",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"2a05",x"3593",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2a24"),
(x"3710",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2dbb",x"36f7",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2d8d",x"3710",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2dbb"),
(x"380a",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2f8b",x"380a",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2f8b",x"37b8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ee7"),
(x"37a8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ec9",x"37b8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ee7",x"37a8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2ec9"),
(x"37a8",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"2ec9",x"37a8",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"2ec9",x"378c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2e97"),
(x"376c",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"2e5e",x"378c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2e97",x"376c",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"2e5e"),
(x"376c",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"2e5e",x"376c",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"2e5e",x"3752",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2e30"),
(x"36e3",x"405a",x"3710",x"0000",x"0000",x"3c00",x"39ec",x"2d6a",x"36f7",x"405b",x"3710",x"0000",x"0000",x"3c00",x"39ee",x"2d8e",x"36df",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"2d63"),
(x"36df",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"2d63",x"3716",x"405a",x"3710",x"0000",x"0000",x"3c00",x"39ed",x"2dc4",x"36dc",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2d5e"),
(x"36e3",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ae",x"2d6a",x"36df",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"2d63",x"36f7",x"4034",x"3710",x"0000",x"0000",x"3c00",x"39ac",x"2d8e"),
(x"36df",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"2d63",x"36dc",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2d5e",x"3716",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ad",x"2dc4"),
(x"3760",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2e49",x"3753",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b0",x"2e32",x"375f",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2e47"),
(x"375f",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"2e47",x"3742",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2e14",x"3754",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"2e33"),
(x"3742",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2e14",x"3753",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39ea",x"2e32",x"375f",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e4",x"2e47"),
(x"372e",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2df0",x"3742",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2e14",x"3754",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"2e33"),
(x"3705",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"2da6",x"36cb",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2d3f",x"36c4",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"2d33"),
(x"36c2",x"403d",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"2d2f",x"36cb",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39be",x"2d3f",x"36c4",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"2d33"),
(x"36c4",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"2d33",x"3705",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"2da6",x"36dc",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b4",x"2d5e"),
(x"3713",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2dbf",x"3705",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"2da6",x"36dc",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e6",x"2d5e"),
(x"3754",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"2e33",x"3713",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2dbf",x"372e",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"2df0"),
(x"3754",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"2e33",x"372e",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"2df0",x"3713",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"2dbf"),
(x"3716",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2dc5",x"3713",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"2dbf",x"3752",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"2e30"),
(x"3754",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"2e33",x"3713",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"2dbf",x"3752",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2e30"),
(x"3716",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2dc5",x"3710",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2dbb",x"3716",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2dc5"),
(x"3716",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2dc5",x"3716",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2dc5",x"3752",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"2e30"),
(x"380a",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d7",x"2f8b",x"3813",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2fac",x"380a",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2f8b"),
(x"3813",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"2fac",x"382a",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2ffc",x"3813",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c3",x"2fac"),
(x"382a",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2ffc",x"3885",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30a2",x"382a",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"2ffc"),
(x"3885",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30a2",x"3885",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30a2",x"388c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30ad"),
(x"38d5",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"3130",x"38bf",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"3109",x"38d5",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"3130"),
(x"38bf",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"3109",x"38bf",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"3109",x"38b2",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"30f1"),
(x"38b2",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d9",x"30f1",x"38b2",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c1",x"30f1",x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed"),
(x"388c",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30ad",x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed",x"388c",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"30ad"),
(x"386c",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"3075",x"3872",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"3080",x"386d",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3076"),
(x"3872",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"3080",x"3885",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"30a2",x"3877",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3088"),
(x"386c",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"3075",x"386d",x"4056",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3076",x"3872",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"3080"),
(x"3872",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"3080",x"3877",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3088",x"3885",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"30a2"),
(x"3885",x"404f",x"3710",x"0000",x"0000",x"3c00",x"39da",x"30a2",x"3894",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39ec",x"30bc",x"388c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"30ae"),
(x"3885",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39c0",x"30a2",x"388c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"30ae",x"3894",x"4035",x"3710",x"0000",x"0000",x"3c00",x"39ae",x"30bc"),
(x"38d9",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b6",x"3136",x"38d8",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3135",x"38d4",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"312d"),
(x"38c7",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"3117",x"38d8",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3135",x"38d4",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"312d"),
(x"38b7",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"30f9",x"38c7",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"3117",x"38c9",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"311a"),
(x"38d4",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"312d",x"38c7",x"4038",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"3117",x"38c9",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39ba",x"311a"),
(x"38b2",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"30f2",x"388c",x"4041",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"30ae",x"38b0",x"403f",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"30ed"),
(x"388c",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"30ad",x"388c",x"404e",x"3710",x"0000",x"0000",x"3c00",x"39d8",x"30ae",x"38b0",x"4050",x"3710",x"0000",x"0000",x"3c00",x"39db",x"30ed"),
(x"38d5",x"404c",x"3710",x"0000",x"0000",x"3c00",x"39d5",x"3130",x"38f6",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"316b",x"38d5",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c5",x"3130"),
(x"38f6",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c4",x"316b",x"38f6",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"316b",x"3915",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"31a2"),
(x"3915",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"31a2",x"392f",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"31d0",x"3915",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"31a2"),
(x"392f",x"4057",x"3710",x"0000",x"0000",x"3c00",x"39e8",x"31d0",x"393f",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"31ed",x"392f",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b2",x"31d0"),
(x"393f",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"31ed",x"3953",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3211",x"393f",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"31ed"),
(x"3953",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3211",x"3953",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3211",x"395a",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"321d"),
(x"395a",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"321d",x"395d",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"3222",x"395a",x"4039",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"321d"),
(x"395d",x"403b",x"3710",x"0000",x"0000",x"3c00",x"39b8",x"3222",x"395d",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e2",x"3222",x"3963",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"322d"),
(x"3963",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"322d",x"3972",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"3248",x"3963",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"322d"),
(x"3972",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e1",x"3248",x"3985",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3269",x"3972",x"403c",x"3710",x"0000",x"0000",x"3c00",x"39b9",x"3248"),
(x"3985",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b5",x"3269",x"3985",x"4055",x"3710",x"0000",x"0000",x"3c00",x"39e5",x"3269",x"3994",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3284"),
(x"3994",x"4058",x"3710",x"0000",x"0000",x"3c00",x"39e9",x"3284",x"3999",x"4058",x"3710",x"935f",x"1e0a",x"3c00",x"39e9",x"328d",x"3994",x"4037",x"3710",x"0000",x"0000",x"3c00",x"39b1",x"3284"),
(x"3999",x"4037",x"3710",x"975f",x"9f93",x"3c00",x"39b1",x"328d",x"3999",x"4058",x"3710",x"935f",x"1e0a",x"3c00",x"39e9",x"328d",x"39fc",x"4042",x"3713",x"ac0e",x"a310",x"3bfb",x"39c4",x"333e"),
(x"3999",x"4058",x"3710",x"935f",x"1e0a",x"3c00",x"39e9",x"328d",x"39f5",x"4059",x"3710",x"b60b",x"25b5",x"3b67",x"39eb",x"3331",x"39fb",x"404d",x"3713",x"a9a8",x"a460",x"3bfd",x"39d7",x"333d"),
(x"3a14",x"4059",x"374f",x"a8f0",x"3bfa",x"ac25",x"3a17",x"3bac",x"3a0d",x"4059",x"374b",x"a412",x"3bfd",x"295c",x"3a18",x"3ba9",x"3a1a",x"4059",x"3749",x"a2b5",x"3bfe",x"281b",x"3a18",x"3bae"),
(x"3a1a",x"4059",x"3749",x"a2b5",x"3bfe",x"281b",x"3a18",x"3bae",x"3a07",x"4059",x"373c",x"a752",x"3bff",x"9bfc",x"3a1b",x"3ba6",x"3a21",x"4059",x"373a",x"a884",x"3bfe",x"253f",x"3a1b",x"3bb1"),
(x"3a21",x"4059",x"373a",x"a884",x"3bfe",x"253f",x"3a1b",x"3bb1",x"3a00",x"4059",x"3722",x"23fc",x"3bf8",x"2d58",x"3a1f",x"3ba4",x"3a24",x"4059",x"372b",x"a504",x"3bff",x"9a59",x"3a1e",x"3bb2"),
(x"3a24",x"4059",x"372b",x"a504",x"3bff",x"9a59",x"3a1e",x"3bb2",x"39fc",x"4059",x"3718",x"135f",x"3bfd",x"29a5",x"3a21",x"3ba2",x"3a27",x"4059",x"3710",x"a3ef",x"3bff",x"9818",x"3a23",x"3bb3"),
(x"3a14",x"4036",x"374e",x"a81b",x"bbe6",x"b0f3",x"3a13",x"3ba9",x"3a19",x"4036",x"3749",x"208e",x"bc00",x"135f",x"3a12",x"3bab",x"3a0d",x"4036",x"374b",x"1481",x"bbff",x"26ae",x"3a12",x"3ba6"),
(x"3a19",x"4036",x"3749",x"208e",x"bc00",x"135f",x"3a12",x"3bab",x"3a20",x"4036",x"3732",x"1f93",x"bc00",x"975f",x"3a0d",x"3bae",x"3a07",x"4036",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a0f",x"3ba4"),
(x"3a20",x"4036",x"3732",x"1f93",x"bc00",x"975f",x"3a0d",x"3bae",x"3a26",x"4036",x"3710",x"1f45",x"bbff",x"a032",x"3a07",x"3bb0",x"3a02",x"4036",x"3724",x"1c81",x"bbff",x"a1c9",x"3a0b",x"3ba2"),
(x"3501",x"403e",x"36da",x"ada8",x"bbf8",x"8000",x"3a50",x"3b93",x"34e9",x"403f",x"36da",x"b698",x"bb49",x"8000",x"3a50",x"3b8e",x"3501",x"403e",x"3710",x"2d0c",x"bbf9",x"0000",x"3a5a",x"3b93"),
(x"386c",x"403c",x"36da",x"bb38",x"36e2",x"868d",x"3a72",x"3ad8",x"3872",x"403e",x"36da",x"b902",x"3a3c",x"0000",x"3a72",x"3ad4",x"386c",x"403c",x"3710",x"bbdd",x"31e1",x"0000",x"3a7c",x"3ad8"),
(x"380a",x"404d",x"36da",x"ad54",x"3bf8",x"8000",x"3a8b",x"3b4a",x"3813",x"404e",x"36da",x"27fc",x"3bfe",x"0000",x"3a8b",x"3b47",x"380a",x"404d",x"3710",x"ae11",x"3bf6",x"0000",x"3a96",x"3b4a"),
(x"34e9",x"403f",x"36da",x"b698",x"bb49",x"8000",x"3a50",x"3b8e",x"34cb",x"4041",x"36da",x"b501",x"bb99",x"0000",x"3a50",x"3b87",x"34e9",x"403f",x"3710",x"b50d",x"bb97",x"0000",x"3a5a",x"3b8e"),
(x"3a26",x"4036",x"36da",x"1e3f",x"bc00",x"0000",x"39fd",x"3bb0",x"39fc",x"4036",x"36da",x"a111",x"bc00",x"0000",x"39fd",x"3b9f",x"3a26",x"4036",x"3710",x"1f45",x"bbff",x"a032",x"3a07",x"3bb0"),
(x"3872",x"403e",x"36da",x"b902",x"3a3c",x"0000",x"3a72",x"3ad4",x"3885",x"4040",x"36da",x"b83d",x"3ac8",x"0000",x"3a72",x"3acc",x"3872",x"403e",x"3710",x"b9d1",x"397d",x"8000",x"3a7c",x"3ad4"),
(x"3760",x"4056",x"36da",x"3bfa",x"2cac",x"868d",x"3a8b",x"3b79",x"375f",x"4055",x"36da",x"3b14",x"b774",x"0000",x"3a8b",x"3b77",x"3760",x"4056",x"3710",x"3b92",x"3528",x"8000",x"3a96",x"3b79"),
(x"34cb",x"4041",x"36da",x"b501",x"bb99",x"0000",x"3a50",x"3b87",x"34bb",x"4042",x"36da",x"b13f",x"bbe4",x"0000",x"3a50",x"3b84",x"34cb",x"4041",x"3710",x"b64c",x"bb5a",x"0000",x"3a5a",x"3b87"),
(x"3885",x"4040",x"36da",x"b83d",x"3ac8",x"0000",x"3a72",x"3acc",x"388c",x"4041",x"36da",x"bbfd",x"29ab",x"0000",x"3a72",x"3ac9",x"3885",x"4040",x"3710",x"b7eb",x"3af3",x"0000",x"3a7c",x"3acc"),
(x"37b8",x"404c",x"36da",x"2df3",x"3bf7",x"0000",x"3a8b",x"3b5c",x"380a",x"404d",x"36da",x"ad54",x"3bf8",x"8000",x"3a8b",x"3b4a",x"37b8",x"404c",x"3710",x"30d0",x"3be8",x"0000",x"3a96",x"3b5c"),
(x"34bb",x"4042",x"36da",x"b13f",x"bbe4",x"0000",x"3a50",x"3b84",x"349b",x"4042",x"36da",x"b4a8",x"bba7",x"8000",x"3a50",x"3b7e",x"34bb",x"4042",x"3710",x"b31c",x"bbcc",x"0000",x"3a5a",x"3b84"),
(x"388c",x"4041",x"36da",x"bbfd",x"29ab",x"0000",x"3a72",x"3ac9",x"388c",x"4042",x"36da",x"b967",x"b9e6",x"0000",x"3a72",x"3ac8",x"388c",x"4041",x"3710",x"bb54",x"3669",x"8000",x"3a7c",x"3ac9"),
(x"37a8",x"404c",x"36da",x"33d5",x"3bc1",x"0000",x"3a8b",x"3b5f",x"37b8",x"404c",x"36da",x"2df3",x"3bf7",x"0000",x"3a8b",x"3b5c",x"37a8",x"404c",x"3710",x"3580",x"3b83",x"0000",x"3a96",x"3b5f"),
(x"349b",x"4042",x"36da",x"b4a8",x"bba7",x"8000",x"3a50",x"3b7e",x"3485",x"4043",x"36da",x"b92c",x"ba1a",x"8000",x"3a50",x"3b7a",x"349b",x"4042",x"3710",x"b221",x"bbda",x"0000",x"3a5a",x"3b7e"),
(x"388c",x"4042",x"36da",x"b967",x"b9e6",x"0000",x"3a42",x"3bb0",x"3885",x"4042",x"36da",x"b25f",x"bbd7",x"0000",x"3a42",x"3bad",x"388c",x"4042",x"3710",x"bb52",x"b671",x"0000",x"3a4c",x"3bb0"),
(x"378c",x"404e",x"36da",x"373a",x"3b23",x"0000",x"3a8b",x"3b65",x"37a8",x"404c",x"36da",x"33d5",x"3bc1",x"0000",x"3a8b",x"3b5f",x"378c",x"404e",x"3710",x"3688",x"3b4d",x"8000",x"3a96",x"3b65"),
(x"3a26",x"404d",x"36da",x"3310",x"3bcd",x"0000",x"3b16",x"3819",x"3a2f",x"404d",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"3816",x"3a26",x"404d",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3820"),
(x"3485",x"4043",x"36da",x"b92c",x"ba1a",x"8000",x"3a50",x"3b7a",x"3475",x"4045",x"36da",x"bbab",x"b48e",x"0000",x"3a50",x"3b75",x"3485",x"4043",x"3710",x"b819",x"bade",x"0000",x"3a5a",x"3b7a"),
(x"3760",x"4038",x"36da",x"3b92",x"b528",x"0000",x"3a42",x"3b4c",x"3753",x"4037",x"36da",x"37e4",x"baf5",x"8000",x"3a42",x"3b48",x"3760",x"4038",x"3710",x"3bfa",x"acac",x"868d",x"3a4c",x"3b4c"),
(x"376c",x"4050",x"36da",x"3787",x"3b0e",x"0000",x"3a8b",x"3b6c",x"378c",x"404e",x"36da",x"373a",x"3b23",x"0000",x"3a8b",x"3b65",x"376c",x"4050",x"3710",x"3899",x"3a8b",x"0000",x"3a96",x"3b6c"),
(x"3885",x"4042",x"36da",x"b25f",x"bbd7",x"0000",x"3a42",x"3bad",x"382a",x"4042",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b89",x"3885",x"4042",x"3710",x"b304",x"bbce",x"0000",x"3a4c",x"3bad"),
(x"3752",x"4053",x"36da",x"3be0",x"31a3",x"8000",x"3a8b",x"3b72",x"376c",x"4050",x"36da",x"3787",x"3b0e",x"0000",x"3a8b",x"3b6c",x"3752",x"4053",x"3710",x"3bfd",x"aac2",x"0000",x"3a96",x"3b72"),
(x"39fc",x"4036",x"36da",x"a111",x"bc00",x"0000",x"39fd",x"3b9f",x"3999",x"4037",x"36da",x"b32b",x"bbcb",x"0000",x"39fd",x"3b78",x"39fc",x"4036",x"3710",x"9bc8",x"bc00",x"200b",x"3a07",x"3b9f"),
(x"382a",x"4042",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b89",x"3813",x"4041",x"36da",x"a8bf",x"bbfe",x"8000",x"3a42",x"3b80",x"382a",x"4042",x"3710",x"2f40",x"bbf2",x"0000",x"3a4c",x"3b89"),
(x"3742",x"4059",x"36da",x"342c",x"3bb9",x"8000",x"3a8b",x"3b80",x"3753",x"4058",x"36da",x"38fe",x"3a3f",x"8000",x"3a8b",x"3b7d",x"3742",x"4059",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b80"),
(x"3813",x"4041",x"36da",x"a8bf",x"bbfe",x"8000",x"3a42",x"3b80",x"380a",x"4041",x"36da",x"ae12",x"bbf6",x"0000",x"3a42",x"3b7c",x"3813",x"4041",x"3710",x"27fc",x"bbfe",x"0000",x"3a4c",x"3b80"),
(x"372e",x"4059",x"36da",x"2fc6",x"3bf0",x"0000",x"3a8b",x"3b84",x"3742",x"4059",x"36da",x"342c",x"3bb9",x"8000",x"3a8b",x"3b80",x"372e",x"4059",x"3710",x"338a",x"3bc6",x"0000",x"3a96",x"3b84"),
(x"375f",x"403a",x"36da",x"3bc1",x"33d8",x"868d",x"3a42",x"3b4e",x"3760",x"4038",x"36da",x"3b92",x"b528",x"0000",x"3a42",x"3b4c",x"375f",x"403a",x"3710",x"3b14",x"3774",x"8000",x"3a4c",x"3b4e"),
(x"3716",x"405a",x"36da",x"34b5",x"3ba5",x"8000",x"3a8b",x"3b89",x"372e",x"4059",x"36da",x"2fc6",x"3bf0",x"0000",x"3a8b",x"3b84",x"3716",x"405a",x"3710",x"32c2",x"3bd1",x"8000",x"3a96",x"3b89"),
(x"380a",x"4041",x"36da",x"ae12",x"bbf6",x"0000",x"3a42",x"3b7c",x"37b8",x"4043",x"36da",x"30d0",x"bbe8",x"0000",x"3a42",x"3b6a",x"380a",x"4041",x"3710",x"ad56",x"bbf8",x"0000",x"3a4c",x"3b7c"),
(x"36f7",x"405b",x"36da",x"ae6b",x"3bf5",x"0000",x"3a8b",x"3b8f",x"3716",x"405a",x"36da",x"34b5",x"3ba5",x"8000",x"3a8b",x"3b89",x"36f7",x"405b",x"3710",x"b463",x"3bb1",x"8000",x"3a96",x"3b8f"),
(x"37b8",x"4043",x"36da",x"30d0",x"bbe8",x"0000",x"3a42",x"3b6a",x"37a8",x"4043",x"36da",x"3580",x"bb83",x"0000",x"3a42",x"3b66",x"37b8",x"4043",x"3710",x"2df5",x"bbf7",x"0000",x"3a4c",x"3b6a"),
(x"36e3",x"405a",x"36da",x"b9b5",x"399a",x"0000",x"3a8b",x"3b93",x"36f7",x"405b",x"36da",x"ae6b",x"3bf5",x"0000",x"3a8b",x"3b8f",x"36e3",x"405a",x"3710",x"bb17",x"3766",x"868d",x"3a96",x"3b93"),
(x"37a8",x"4043",x"36da",x"3580",x"bb83",x"0000",x"3a42",x"3b66",x"378c",x"4041",x"36da",x"3688",x"bb4d",x"8000",x"3a42",x"3b60",x"37a8",x"4043",x"3710",x"33d5",x"bbc1",x"0000",x"3a4c",x"3b66"),
(x"36df",x"4058",x"36da",x"bbbc",x"3412",x"0000",x"3a8b",x"3b96",x"36e3",x"405a",x"36da",x"b9b5",x"399a",x"0000",x"3a8b",x"3b93",x"36df",x"4058",x"3710",x"bbc6",x"338f",x"8000",x"3a96",x"3b96"),
(x"378c",x"4041",x"36da",x"3688",x"bb4d",x"8000",x"3a42",x"3b60",x"376c",x"403f",x"36da",x"3899",x"ba8b",x"0000",x"3a42",x"3b59",x"378c",x"4041",x"3710",x"373a",x"bb23",x"0000",x"3a4c",x"3b60"),
(x"36dc",x"4056",x"36da",x"bba4",x"34ba",x"0000",x"3a8b",x"3b98",x"36df",x"4058",x"36da",x"bbbc",x"3412",x"0000",x"3a8b",x"3b96",x"36dc",x"4056",x"3710",x"bb3a",x"36da",x"0000",x"3a96",x"3b98"),
(x"3a27",x"4059",x"36da",x"3bff",x"a4d0",x"0000",x"39e9",x"33f9",x"3a26",x"404d",x"36da",x"3bff",x"a4d0",x"0000",x"39d6",x"33f3",x"3a27",x"4059",x"3710",x"3bea",x"a4d6",x"30a2",x"39ea",x"33c9"),
(x"3999",x"4058",x"36da",x"b2b0",x"3bd2",x"0000",x"3a2d",x"3b7b",x"39f5",x"4059",x"36da",x"a49b",x"3bff",x"8000",x"3a2d",x"3b9f",x"3999",x"4058",x"3710",x"b329",x"3bcb",x"8000",x"3a23",x"3b7b"),
(x"376c",x"403f",x"36da",x"3899",x"ba8b",x"0000",x"3a42",x"3b59",x"3752",x"403c",x"36da",x"3bfd",x"2ac2",x"0000",x"3a42",x"3b53",x"376c",x"403f",x"3710",x"3787",x"bb0e",x"0000",x"3a4c",x"3b59"),
(x"36c4",x"4053",x"36da",x"bb61",x"362a",x"0000",x"3a8b",x"3b9f",x"36dc",x"4056",x"36da",x"bba4",x"34ba",x"0000",x"3a8b",x"3b98",x"36c4",x"4053",x"3710",x"bbc5",x"339b",x"068d",x"3a96",x"3b9f"),
(x"3994",x"4058",x"36da",x"b458",x"3bb2",x"8000",x"3a2d",x"3b79",x"3999",x"4058",x"36da",x"b2b0",x"3bd2",x"0000",x"3a2d",x"3b7b",x"3994",x"4058",x"3710",x"b59f",x"3b7d",x"0000",x"3a23",x"3b79"),
(x"3753",x"4037",x"36da",x"37e4",x"baf5",x"8000",x"3a42",x"3b48",x"3742",x"4036",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b44",x"3753",x"4037",x"3710",x"38fe",x"ba3f",x"0000",x"3a4c",x"3b48"),
(x"36c2",x"4051",x"36da",x"bbe7",x"b0ec",x"0000",x"3a8b",x"3ba1",x"36c4",x"4053",x"36da",x"bb61",x"362a",x"0000",x"3a8b",x"3b9f",x"36c2",x"4051",x"3710",x"bafe",x"b7c2",x"0000",x"3a96",x"3ba1"),
(x"3985",x"4055",x"36da",x"b817",x"3adf",x"0000",x"3a2d",x"3b72",x"3994",x"4058",x"36da",x"b458",x"3bb2",x"8000",x"3a2d",x"3b79",x"3985",x"4055",x"3710",x"b796",x"3b0b",x"0000",x"3a23",x"3b72"),
(x"3742",x"4036",x"36da",x"30bd",x"bbe9",x"0000",x"3a42",x"3b44",x"372e",x"4036",x"36da",x"338a",x"bbc6",x"0000",x"3a42",x"3b40",x"3742",x"4036",x"3710",x"342c",x"bbb9",x"0000",x"3a4c",x"3b44"),
(x"36cb",x"4050",x"36da",x"b922",x"ba22",x"068d",x"3a8b",x"3ba3",x"36c2",x"4051",x"36da",x"bbe7",x"b0ec",x"0000",x"3a8b",x"3ba1",x"36cb",x"4050",x"3710",x"b86c",x"baa9",x"0000",x"3a96",x"3ba3"),
(x"3972",x"4053",x"36da",x"b475",x"3bae",x"0000",x"3a2d",x"3b6a",x"3985",x"4055",x"36da",x"b817",x"3adf",x"0000",x"3a2d",x"3b72",x"3972",x"4053",x"3710",x"b0a0",x"3bea",x"0000",x"3a23",x"3b6a"),
(x"372e",x"4036",x"36da",x"338a",x"bbc6",x"0000",x"3a42",x"3b40",x"3716",x"4035",x"36da",x"32c2",x"bbd1",x"0000",x"3a42",x"3b3b",x"372e",x"4036",x"3710",x"2fc6",x"bbf0",x"0000",x"3a4c",x"3b40"),
(x"3705",x"404f",x"36da",x"b599",x"bb7e",x"0000",x"3a8b",x"3bae",x"36cb",x"4050",x"36da",x"b922",x"ba22",x"068d",x"3a8b",x"3ba3",x"3705",x"404f",x"3710",x"b675",x"bb51",x"0000",x"3a96",x"3bae"),
(x"3963",x"4053",x"36da",x"3420",x"3bba",x"0000",x"3a2d",x"3b64",x"3972",x"4053",x"36da",x"b475",x"3bae",x"0000",x"3a2d",x"3b6a",x"3963",x"4053",x"3710",x"36c5",x"3b3f",x"0000",x"3a23",x"3b64"),
(x"3716",x"4035",x"36da",x"32c2",x"bbd1",x"0000",x"3a42",x"3b3b",x"36f7",x"4034",x"36da",x"b463",x"bbb1",x"8000",x"3a42",x"3b35",x"3716",x"4035",x"3710",x"34b5",x"bba5",x"0000",x"3a4c",x"3b3b"),
(x"3713",x"404e",x"36da",x"b972",x"b9db",x"8000",x"3a8b",x"3bb1",x"3705",x"404f",x"36da",x"b599",x"bb7e",x"0000",x"3a8b",x"3bae",x"3713",x"404e",x"3710",x"ba37",x"b909",x"0000",x"3a96",x"3bb1"),
(x"395d",x"4054",x"36da",x"399d",x"39b2",x"0000",x"3a2d",x"3b61",x"3963",x"4053",x"36da",x"3420",x"3bba",x"0000",x"3a2d",x"3b64",x"395d",x"4054",x"3710",x"3ac1",x"3849",x"0000",x"3a23",x"3b61"),
(x"36f7",x"4034",x"36da",x"b463",x"bbb1",x"8000",x"3a42",x"3b35",x"36e3",x"4035",x"36da",x"bb17",x"b766",x"068d",x"3a42",x"3b31",x"36f7",x"4034",x"3710",x"ae6b",x"bbf5",x"0000",x"3a4c",x"3b35"),
(x"3716",x"404e",x"36da",x"bbb8",x"b42d",x"0000",x"3a8b",x"3bb2",x"3713",x"404e",x"36da",x"b972",x"b9db",x"8000",x"3a8b",x"3bb1",x"3716",x"404e",x"3710",x"bbad",x"3480",x"0000",x"3a96",x"3bb2"),
(x"395a",x"4055",x"36da",x"3b46",x"36a7",x"8000",x"3a2d",x"3b5e",x"395d",x"4054",x"36da",x"399d",x"39b2",x"0000",x"3a2d",x"3b61",x"395a",x"4055",x"3710",x"3af1",x"37f3",x"0000",x"3a23",x"3b5e"),
(x"36e3",x"4035",x"36da",x"bb17",x"b766",x"068d",x"3a42",x"3b31",x"36df",x"4037",x"36da",x"bbc6",x"b38f",x"8000",x"3a42",x"3b2e",x"36e3",x"4035",x"3710",x"b9b5",x"b99a",x"0000",x"3a4c",x"3b31"),
(x"3710",x"404d",x"36da",x"b8f7",x"3a45",x"0000",x"3b11",x"39af",x"3716",x"404e",x"36da",x"bbb8",x"b42d",x"0000",x"3b11",x"39ae",x"3710",x"404d",x"3710",x"b80d",x"3ae5",x"0000",x"3b1c",x"39af"),
(x"3953",x"4058",x"36da",x"39a8",x"39a7",x"868d",x"3a2d",x"3b5a",x"395a",x"4055",x"36da",x"3b46",x"36a7",x"8000",x"3a2d",x"3b5e",x"3953",x"4058",x"3710",x"3857",x"3ab8",x"8000",x"3a23",x"3b5a"),
(x"36df",x"4037",x"36da",x"bbc6",x"b38f",x"8000",x"3a42",x"3b2e",x"36dc",x"4038",x"36da",x"bb3a",x"b6d9",x"0000",x"3a42",x"3b2b",x"36df",x"4037",x"3710",x"bbbc",x"b412",x"0000",x"3a4c",x"3b2e"),
(x"36f7",x"404c",x"36da",x"b12d",x"3be4",x"0000",x"3b11",x"39b4",x"3710",x"404d",x"36da",x"b8f7",x"3a45",x"0000",x"3b11",x"39af",x"36f7",x"404c",x"3710",x"b05b",x"3bec",x"8000",x"3b1c",x"39b4"),
(x"3475",x"4045",x"36da",x"bbab",x"b48e",x"0000",x"3a50",x"3b75",x"3475",x"404a",x"36da",x"baeb",x"3803",x"8000",x"3a50",x"3b6f",x"3475",x"4045",x"3710",x"baeb",x"b803",x"0000",x"3a5a",x"3b75"),
(x"393f",x"4059",x"36da",x"1cea",x"3c00",x"0000",x"3a2d",x"3b51",x"3953",x"4058",x"36da",x"39a8",x"39a7",x"868d",x"3a2d",x"3b5a",x"393f",x"4059",x"3710",x"b2bb",x"3bd2",x"868d",x"3a23",x"3b51"),
(x"36dc",x"4038",x"36da",x"bb3a",x"b6d9",x"0000",x"3a42",x"3b2b",x"36c4",x"403c",x"36da",x"bbc5",x"b39b",x"0000",x"3a42",x"3b24",x"36dc",x"4038",x"3710",x"bba4",x"b4ba",x"0000",x"3a4c",x"3b2b"),
(x"362c",x"404d",x"36da",x"3550",x"3b8b",x"0000",x"3b11",x"39db",x"363b",x"404c",x"36da",x"3439",x"3bb7",x"0000",x"3b11",x"39d8",x"362c",x"404d",x"3710",x"3609",x"3b68",x"8000",x"3b1c",x"39db"),
(x"3999",x"4037",x"36da",x"b32b",x"bbcb",x"0000",x"39fd",x"3b78",x"3994",x"4037",x"36da",x"b59f",x"bb7d",x"0000",x"39fd",x"3b76",x"3999",x"4037",x"3710",x"b2ba",x"bbd2",x"0000",x"3a07",x"3b78"),
(x"392f",x"4057",x"36da",x"b73b",x"3b22",x"8000",x"3a2d",x"3b4b",x"393f",x"4059",x"36da",x"1cea",x"3c00",x"0000",x"3a2d",x"3b51",x"392f",x"4057",x"3710",x"b874",x"3aa4",x"0000",x"3a23",x"3b4b"),
(x"36c4",x"403c",x"36da",x"bbc5",x"b39b",x"0000",x"3a42",x"3b24",x"36c2",x"403d",x"36da",x"bafe",x"37c2",x"8000",x"3a42",x"3b22",x"36c4",x"403c",x"3710",x"bb61",x"b62a",x"0000",x"3a4c",x"3b24"),
(x"363b",x"404c",x"36da",x"3439",x"3bb7",x"0000",x"3b11",x"39d8",x"36f7",x"404c",x"36da",x"b12d",x"3be4",x"0000",x"3b11",x"39b4",x"363b",x"404c",x"3710",x"34bd",x"3ba4",x"0000",x"3b1c",x"39d8"),
(x"3994",x"4037",x"36da",x"b59f",x"bb7d",x"0000",x"39fd",x"3b76",x"3985",x"403a",x"36da",x"b796",x"bb0b",x"0000",x"39fd",x"3b6f",x"3994",x"4037",x"3710",x"b459",x"bbb2",x"068d",x"3a07",x"3b76"),
(x"3754",x"4054",x"36da",x"3ba5",x"b4b5",x"0000",x"3a8b",x"3b74",x"3752",x"4053",x"36da",x"3be0",x"31a3",x"8000",x"3a8b",x"3b72",x"3754",x"4054",x"3710",x"3afe",x"b7c4",x"0000",x"3a96",x"3b74"),
(x"36c2",x"403d",x"36da",x"bafe",x"37c2",x"8000",x"3a42",x"3b22",x"36cb",x"403e",x"36da",x"b86c",x"3aaa",x"0000",x"3a42",x"3b1f",x"36c2",x"403d",x"3710",x"bbe7",x"30ec",x"868d",x"3a4c",x"3b22"),
(x"35f7",x"4051",x"36da",x"3a05",x"3944",x"868d",x"3b11",x"39e6",x"362c",x"404d",x"36da",x"3550",x"3b8b",x"0000",x"3b11",x"39db",x"35f7",x"4051",x"3710",x"3a6a",x"38c7",x"0000",x"3b1c",x"39e6"),
(x"3985",x"403a",x"36da",x"b796",x"bb0b",x"0000",x"39fd",x"3b6f",x"3972",x"403c",x"36da",x"b0a0",x"bbea",x"0000",x"39fd",x"3b67",x"3985",x"403a",x"3710",x"b817",x"badf",x"0000",x"3a07",x"3b6f"),
(x"3915",x"4051",x"36da",x"b90a",x"3a36",x"0000",x"3a2d",x"3b3c",x"392f",x"4057",x"36da",x"b73b",x"3b22",x"8000",x"3a2d",x"3b4b",x"3915",x"4051",x"3710",x"b845",x"3ac3",x"0000",x"3a23",x"3b3c"),
(x"36cb",x"403e",x"36da",x"b86c",x"3aaa",x"0000",x"3a42",x"3b1f",x"3705",x"4040",x"36da",x"b675",x"3b51",x"0000",x"3a42",x"3b14",x"36cb",x"403e",x"3710",x"b922",x"3a22",x"0000",x"3a4c",x"3b1f"),
(x"35f1",x"4052",x"36da",x"3bcd",x"3318",x"0000",x"3b11",x"39e8",x"35f7",x"4051",x"36da",x"3a05",x"3944",x"868d",x"3b11",x"39e6",x"35f1",x"4052",x"3710",x"3bf9",x"ad20",x"0000",x"3b1c",x"39e8"),
(x"3972",x"403c",x"36da",x"b0a0",x"bbea",x"0000",x"39fd",x"3b67",x"3963",x"403c",x"36da",x"36c5",x"bb3f",x"0000",x"39fd",x"3b61",x"3972",x"403c",x"3710",x"b475",x"bbae",x"0000",x"3a07",x"3b67"),
(x"375f",x"4055",x"36da",x"3b14",x"b774",x"0000",x"3a8b",x"3b77",x"3754",x"4054",x"36da",x"3ba5",x"b4b5",x"0000",x"3a8b",x"3b74",x"375f",x"4055",x"3710",x"3bc1",x"b3d8",x"0000",x"3a96",x"3b77"),
(x"3705",x"4040",x"36da",x"b675",x"3b51",x"0000",x"3a42",x"3b14",x"3713",x"4041",x"36da",x"ba37",x"3909",x"0000",x"3a42",x"3b11",x"3705",x"4040",x"3710",x"b599",x"3b7e",x"0000",x"3a4c",x"3b14"),
(x"35f3",x"4053",x"36da",x"3b84",x"b57a",x"0000",x"3b11",x"39e9",x"35f1",x"4052",x"36da",x"3bcd",x"3318",x"0000",x"3b11",x"39e8",x"35f3",x"4053",x"3710",x"3b36",x"b6ea",x"8000",x"3b1c",x"39e9"),
(x"3963",x"403c",x"36da",x"36c5",x"bb3f",x"0000",x"39fd",x"3b61",x"395d",x"403b",x"36da",x"3ac1",x"b849",x"0000",x"39fd",x"3b5e",x"3963",x"403c",x"3710",x"3420",x"bbba",x"0000",x"3a07",x"3b61"),
(x"38f6",x"404d",x"36da",x"b551",x"3b8b",x"0000",x"3a2d",x"3b2e",x"3915",x"4051",x"36da",x"b90a",x"3a36",x"0000",x"3a2d",x"3b3c",x"38f6",x"404d",x"3710",x"b324",x"3bcc",x"0000",x"3a23",x"3b2e"),
(x"3713",x"4041",x"36da",x"ba37",x"3909",x"0000",x"3a42",x"3b11",x"3716",x"4041",x"36da",x"bbad",x"b480",x"0000",x"3a42",x"3b10",x"3713",x"4041",x"3710",x"b972",x"39db",x"0000",x"3a4c",x"3b11"),
(x"35fd",x"4054",x"36da",x"3b91",x"b530",x"8000",x"3b11",x"39ed",x"35f3",x"4053",x"36da",x"3b84",x"b57a",x"0000",x"3b11",x"39e9",x"35fd",x"4054",x"3710",x"3bf0",x"aff4",x"868d",x"3b1c",x"39ed"),
(x"395d",x"403b",x"36da",x"3ac1",x"b849",x"0000",x"39fd",x"3b5e",x"395a",x"4039",x"36da",x"3af1",x"b7f3",x"0000",x"39fd",x"3b5b",x"395d",x"403b",x"3710",x"399d",x"b9b2",x"0000",x"3a07",x"3b5e"),
(x"38d5",x"404c",x"36da",x"1987",x"3c00",x"0000",x"3a2d",x"3b21",x"38f6",x"404d",x"36da",x"b551",x"3b8b",x"0000",x"3a2d",x"3b2e",x"38d5",x"404c",x"3710",x"2dde",x"3bf7",x"0000",x"3a23",x"3b21"),
(x"3716",x"4041",x"36da",x"bbad",x"b480",x"0000",x"3af0",x"3a11",x"3710",x"4042",x"36da",x"b80d",x"bae5",x"8000",x"3af0",x"3a0f",x"3716",x"4041",x"3710",x"bbb8",x"342d",x"0000",x"3afb",x"3a11"),
(x"35fd",x"4055",x"36da",x"3b87",x"3567",x"8000",x"3b11",x"39ee",x"35fd",x"4054",x"36da",x"3b91",x"b530",x"8000",x"3b11",x"39ed",x"35fd",x"4055",x"3710",x"3a08",x"3941",x"0000",x"3b1c",x"39ee"),
(x"395a",x"4039",x"36da",x"3af1",x"b7f3",x"0000",x"39fd",x"3b5b",x"3953",x"4037",x"36da",x"3857",x"bab8",x"8000",x"39fd",x"3b57",x"395a",x"4039",x"3710",x"3b46",x"b6a7",x"8000",x"3a07",x"3b5b"),
(x"38bf",x"404d",x"36da",x"3489",x"3bac",x"0000",x"3a2d",x"3b18",x"38d5",x"404c",x"36da",x"1987",x"3c00",x"0000",x"3a2d",x"3b21",x"38bf",x"404d",x"3710",x"35f3",x"3b6c",x"0000",x"3a23",x"3b18"),
(x"3710",x"4042",x"36da",x"b80d",x"bae5",x"8000",x"3af0",x"3a0f",x"36f7",x"4042",x"36da",x"b05b",x"bbec",x"8000",x"3af0",x"3a0a",x"3710",x"4042",x"3710",x"b8f7",x"ba45",x"0000",x"3afb",x"3a0f"),
(x"35f5",x"4056",x"36da",x"364c",x"3b5a",x"868d",x"3b11",x"39f0",x"35fd",x"4055",x"36da",x"3b87",x"3567",x"8000",x"3b11",x"39ee",x"35f5",x"4056",x"3710",x"32d5",x"3bd0",x"0000",x"3b1c",x"39f0"),
(x"3953",x"4037",x"36da",x"3857",x"bab8",x"8000",x"39fd",x"3b57",x"393f",x"4036",x"36da",x"b2bc",x"bbd2",x"8000",x"39fd",x"3b4e",x"3953",x"4037",x"3710",x"39a8",x"b9a7",x"0000",x"3a07",x"3b57"),
(x"38b2",x"404e",x"36da",x"3a0a",x"393e",x"8000",x"3a2d",x"3b13",x"38bf",x"404d",x"36da",x"3489",x"3bac",x"0000",x"3a2d",x"3b18",x"38b2",x"404e",x"3710",x"3af2",x"37f0",x"0000",x"3a23",x"3b13"),
(x"363b",x"4042",x"36da",x"34be",x"bba4",x"0000",x"3af0",x"39e7",x"362c",x"4042",x"36da",x"3609",x"bb68",x"0000",x"3af0",x"39e4",x"363b",x"4042",x"3710",x"3439",x"bbb7",x"8000",x"3afb",x"39e7"),
(x"35e4",x"4056",x"36da",x"b0fa",x"3be7",x"8000",x"3b11",x"39f3",x"35f5",x"4056",x"36da",x"364c",x"3b5a",x"868d",x"3b11",x"39f0",x"35e4",x"4056",x"3710",x"b3c3",x"3bc2",x"0000",x"3b1c",x"39f3"),
(x"393f",x"4036",x"36da",x"b2bc",x"bbd2",x"8000",x"39fd",x"3b4e",x"392f",x"4037",x"36da",x"b874",x"baa4",x"0000",x"39fd",x"3b48",x"393f",x"4036",x"3710",x"1cea",x"bc00",x"8000",x"3a07",x"3b4e"),
(x"38b0",x"4050",x"36da",x"3bfc",x"2b27",x"0000",x"3a2d",x"3b10",x"38b2",x"404e",x"36da",x"3a0a",x"393e",x"8000",x"3a2d",x"3b13",x"38b0",x"4050",x"3710",x"3ba6",x"b4ab",x"0000",x"3a23",x"3b10"),
(x"36f7",x"4042",x"36da",x"b05b",x"bbec",x"8000",x"3af0",x"3a0a",x"363b",x"4042",x"36da",x"34be",x"bba4",x"0000",x"3af0",x"39e7",x"36f7",x"4042",x"3710",x"b12d",x"bbe4",x"0000",x"3afb",x"3a0a"),
(x"35d3",x"4055",x"36da",x"b1d2",x"3bdd",x"0000",x"3b11",x"39f7",x"35e4",x"4056",x"36da",x"b0fa",x"3be7",x"8000",x"3b11",x"39f3",x"35d3",x"4055",x"3710",x"1c81",x"3c00",x"0000",x"3b1c",x"39f7"),
(x"3752",x"403c",x"36da",x"3bfd",x"2ac2",x"0000",x"3a42",x"3b53",x"3754",x"403b",x"36da",x"3afe",x"37c4",x"0000",x"3a42",x"3b51",x"3752",x"403c",x"3710",x"3be0",x"b1a3",x"068d",x"3a4c",x"3b53"),
(x"38b2",x"4051",x"36da",x"3a58",x"b8de",x"0000",x"3a2d",x"3b0f",x"38b0",x"4050",x"36da",x"3bfc",x"2b27",x"0000",x"3a2d",x"3b10",x"38b2",x"4051",x"3710",x"399c",x"b9b3",x"0000",x"3a23",x"3b0f"),
(x"362c",x"4042",x"36da",x"3609",x"bb68",x"0000",x"3af0",x"39e4",x"35f7",x"403e",x"36da",x"3a6a",x"b8c7",x"0000",x"3af0",x"39d8",x"362c",x"4042",x"3710",x"3550",x"bb8b",x"0000",x"3afb",x"39e4"),
(x"35bd",x"4056",x"36da",x"2c75",x"3bfb",x"068d",x"3b11",x"39fb",x"35d3",x"4055",x"36da",x"b1d2",x"3bdd",x"0000",x"3b11",x"39f7",x"35bd",x"4056",x"3710",x"afcb",x"3bf0",x"8000",x"3b1c",x"39fb"),
(x"392f",x"4037",x"36da",x"b874",x"baa4",x"0000",x"39fd",x"3b48",x"3915",x"403e",x"36da",x"b845",x"bac3",x"0000",x"39fd",x"3b39",x"392f",x"4037",x"3710",x"b73b",x"bb22",x"0000",x"3a07",x"3b48"),
(x"38bd",x"4052",x"36da",x"35fc",x"bb6b",x"0000",x"3a88",x"3ac9",x"38b2",x"4051",x"36da",x"3a58",x"b8de",x"0000",x"3a88",x"3ac5",x"38bd",x"4052",x"3710",x"3456",x"bbb3",x"0000",x"3a93",x"3ac9"),
(x"35f7",x"403e",x"36da",x"3a6a",x"b8c7",x"0000",x"3af0",x"39d8",x"35f1",x"403d",x"36da",x"3bf9",x"2d20",x"0000",x"3af0",x"39d6",x"35f7",x"403e",x"3710",x"3a05",x"b944",x"0000",x"3afb",x"39d8"),
(x"359e",x"4054",x"36da",x"b80b",x"3ae7",x"8000",x"3b11",x"3a01",x"35bd",x"4056",x"36da",x"2c75",x"3bfb",x"068d",x"3b11",x"39fb",x"359e",x"4054",x"3710",x"b925",x"3a1f",x"0000",x"3b1c",x"3a01"),
(x"3754",x"403b",x"36da",x"3afe",x"37c4",x"0000",x"3a42",x"3b51",x"375f",x"403a",x"36da",x"3bc1",x"33d8",x"868d",x"3a42",x"3b4e",x"3754",x"403b",x"3710",x"3ba5",x"34b5",x"0000",x"3a4c",x"3b51"),
(x"38c9",x"4053",x"36da",x"3385",x"bbc6",x"0000",x"3a88",x"3ace",x"38bd",x"4052",x"36da",x"35fc",x"bb6b",x"0000",x"3a88",x"3ac9",x"38c9",x"4053",x"3710",x"34cb",x"bba1",x"0000",x"3a93",x"3ace"),
(x"35f1",x"403d",x"36da",x"3bf9",x"2d20",x"0000",x"3af0",x"39d6",x"35f3",x"403c",x"36da",x"3b36",x"36ea",x"8000",x"3af0",x"39d5",x"35f1",x"403d",x"3710",x"3bcd",x"b318",x"0000",x"3afb",x"39d6"),
(x"358a",x"4051",x"36da",x"bb1e",x"374c",x"8000",x"3b11",x"3a07",x"359e",x"4054",x"36da",x"b80b",x"3ae7",x"8000",x"3b11",x"3a01",x"358a",x"4051",x"3710",x"bbad",x"3481",x"0000",x"3b1c",x"3a07"),
(x"3915",x"403e",x"36da",x"b845",x"bac3",x"0000",x"39fd",x"3b39",x"38f6",x"4042",x"36da",x"b324",x"bbcc",x"0000",x"39fd",x"3b2b",x"3915",x"403e",x"3710",x"b90a",x"ba36",x"0000",x"3a07",x"3b39"),
(x"38d4",x"4054",x"36da",x"37f2",x"baf1",x"8000",x"3a88",x"3ad2",x"38c9",x"4053",x"36da",x"3385",x"bbc6",x"0000",x"3a88",x"3ace",x"38d4",x"4054",x"3710",x"38a8",x"ba80",x"8000",x"3a93",x"3ad2"),
(x"35f3",x"403c",x"36da",x"3b36",x"36ea",x"8000",x"3af0",x"39d5",x"35fd",x"403a",x"36da",x"3bf0",x"2ff4",x"868d",x"3af0",x"39d2",x"35f3",x"403c",x"3710",x"3b84",x"3579",x"0000",x"3afb",x"39d5"),
(x"3587",x"404f",x"36da",x"bbf7",x"adba",x"8000",x"3b11",x"3a0b",x"358a",x"4051",x"36da",x"bb1e",x"374c",x"8000",x"3b11",x"3a07",x"3587",x"404f",x"3710",x"bb8b",x"b553",x"868d",x"3b1c",x"3a0b"),
(x"38f6",x"4042",x"36da",x"b324",x"bbcc",x"0000",x"39fd",x"3b2b",x"38d5",x"4043",x"36da",x"2dde",x"bbf7",x"0000",x"39fd",x"3b1e",x"38f6",x"4042",x"3710",x"b551",x"bb8b",x"0000",x"3a07",x"3b2b"),
(x"38d9",x"4055",x"36da",x"3b88",x"b564",x"0000",x"3a88",x"3ad5",x"38d4",x"4054",x"36da",x"37f2",x"baf1",x"8000",x"3a88",x"3ad2",x"38d9",x"4055",x"3710",x"3bfc",x"ab03",x"8a8d",x"3a93",x"3ad5"),
(x"3a25",x"4041",x"36da",x"3bff",x"26b5",x"0000",x"39c6",x"33f0",x"3a26",x"4036",x"36da",x"3bff",x"26b5",x"0000",x"39b3",x"33fa",x"3a25",x"4041",x"3710",x"3bd6",x"2604",x"3256",x"39c5",x"33c0"),
(x"35fd",x"403a",x"36da",x"3bf0",x"2ff4",x"868d",x"3af0",x"39d2",x"35fd",x"4039",x"36da",x"3a08",x"b941",x"8000",x"3af0",x"39d0",x"35fd",x"403a",x"3710",x"3b91",x"3530",x"0000",x"3afb",x"39d2"),
(x"3593",x"404d",x"36da",x"bbda",x"b21b",x"0000",x"3b11",x"3a0f",x"3587",x"404f",x"36da",x"bbf7",x"adba",x"8000",x"3b11",x"3a0b",x"3593",x"404d",x"3710",x"bc00",x"15bc",x"0000",x"3b1c",x"3a0f"),
(x"38d5",x"4043",x"36da",x"2dde",x"bbf7",x"0000",x"39fd",x"3b1e",x"38bf",x"4042",x"36da",x"35f3",x"bb6c",x"0000",x"39fd",x"3b15",x"38d5",x"4043",x"3710",x"1987",x"bc00",x"0000",x"3a07",x"3b1e"),
(x"38d8",x"4055",x"36da",x"3be4",x"312f",x"8000",x"3a88",x"3ad6",x"38d9",x"4055",x"36da",x"3b88",x"b564",x"0000",x"3a88",x"3ad5",x"38d8",x"4055",x"3710",x"3b96",x"350f",x"0000",x"3a93",x"3ad6"),
(x"35fd",x"4039",x"36da",x"3a08",x"b941",x"8000",x"3af0",x"39d0",x"35f5",x"4039",x"36da",x"32d5",x"bbd0",x"0000",x"3af0",x"39ce",x"35fd",x"4039",x"3710",x"3b87",x"b567",x"868d",x"3afb",x"39d0"),
(x"3592",x"404c",x"36da",x"bba4",x"34bb",x"0000",x"3b11",x"3a11",x"3593",x"404d",x"36da",x"bbda",x"b21b",x"0000",x"3b11",x"3a0f",x"3592",x"404c",x"3710",x"ba08",x"3941",x"0000",x"3b1c",x"3a11"),
(x"38bf",x"4042",x"36da",x"35f3",x"bb6c",x"0000",x"39fd",x"3b15",x"38b2",x"4040",x"36da",x"3af2",x"b7f0",x"0000",x"39fd",x"3b10",x"38bf",x"4042",x"3710",x"3489",x"bbab",x"0000",x"3a07",x"3b15"),
(x"38c7",x"4057",x"36da",x"3653",x"3b59",x"0000",x"3a88",x"3add",x"38d8",x"4055",x"36da",x"3be4",x"312f",x"8000",x"3a88",x"3ad6",x"38c7",x"4057",x"3710",x"364a",x"3b5b",x"0000",x"3a93",x"3add"),
(x"35f5",x"4039",x"36da",x"32d5",x"bbd0",x"0000",x"3af0",x"39ce",x"35e4",x"4039",x"36da",x"b3c3",x"bbc2",x"0000",x"3af0",x"39cb",x"35f5",x"4039",x"3710",x"364b",x"bb5a",x"0000",x"3afb",x"39ce"),
(x"357d",x"404b",x"36da",x"a8c9",x"3bfe",x"0000",x"3a50",x"3b38",x"3592",x"404c",x"36da",x"bba4",x"34bb",x"0000",x"3a50",x"3b34",x"357d",x"404b",x"3710",x"26bb",x"3bff",x"0000",x"3a5a",x"3b38"),
(x"38b2",x"4040",x"36da",x"3af2",x"b7f0",x"0000",x"3b16",x"38a2",x"38b0",x"403f",x"36da",x"3ba6",x"34ac",x"0000",x"3b18",x"38a2",x"38b2",x"4040",x"3710",x"3a0a",x"b93e",x"0000",x"3b16",x"38ac"),
(x"38b7",x"4059",x"36da",x"3528",x"3b92",x"068d",x"3a88",x"3ae4",x"38c7",x"4057",x"36da",x"3653",x"3b59",x"0000",x"3a88",x"3add",x"38b7",x"4059",x"3710",x"32f7",x"3bce",x"0000",x"3a93",x"3ae4"),
(x"35e4",x"4039",x"36da",x"b3c3",x"bbc2",x"0000",x"3af0",x"39cb",x"35d3",x"403a",x"36da",x"1c81",x"bc00",x"0000",x"3af0",x"39c8",x"35e4",x"4039",x"3710",x"b0fa",x"bbe7",x"8000",x"3afb",x"39cb"),
(x"3555",x"404c",x"36da",x"345b",x"3bb2",x"0000",x"3a50",x"3b3f",x"357d",x"404b",x"36da",x"a8c9",x"3bfe",x"0000",x"3a50",x"3b38",x"3555",x"404c",x"3710",x"35eb",x"3b6e",x"0000",x"3a5a",x"3b3f"),
(x"38b0",x"403f",x"36da",x"3ba6",x"34ac",x"0000",x"3b18",x"38a2",x"38b2",x"403e",x"36da",x"399c",x"39b3",x"8000",x"3b1a",x"38a2",x"38b0",x"403f",x"3710",x"3bfc",x"ab27",x"0000",x"3b18",x"38ac"),
(x"3894",x"4059",x"36da",x"aa0a",x"3bfd",x"8000",x"3a88",x"3af1",x"38b7",x"4059",x"36da",x"3528",x"3b92",x"068d",x"3a88",x"3ae4",x"3894",x"4059",x"3710",x"b036",x"3bee",x"0000",x"3a93",x"3af1"),
(x"35d3",x"403a",x"36da",x"1c81",x"bc00",x"0000",x"3af0",x"39c8",x"35bd",x"4039",x"36da",x"afcb",x"bbf0",x"0000",x"3af0",x"39c3",x"35d3",x"403a",x"3710",x"b1d2",x"bbdd",x"0000",x"3afb",x"39c8"),
(x"353f",x"404d",x"36da",x"3746",x"3b1f",x"0000",x"3a50",x"3b44",x"3555",x"404c",x"36da",x"345b",x"3bb2",x"0000",x"3a50",x"3b3f",x"353f",x"404d",x"3710",x"379f",x"3b08",x"0000",x"3a5a",x"3b44"),
(x"38b2",x"403e",x"36da",x"399c",x"39b3",x"8000",x"3b1a",x"38a2",x"38bd",x"403d",x"36da",x"3456",x"3bb3",x"0000",x"3b1e",x"38a2",x"38b2",x"403e",x"3710",x"3a58",x"38de",x"0000",x"3b1a",x"38ac"),
(x"3877",x"4058",x"36da",x"b74e",x"3b1d",x"0000",x"3a88",x"3afc",x"3894",x"4059",x"36da",x"aa0a",x"3bfd",x"8000",x"3a88",x"3af1",x"3877",x"4058",x"3710",x"b8aa",x"3a7f",x"868d",x"3a93",x"3afc"),
(x"35bd",x"4039",x"36da",x"afcb",x"bbf0",x"0000",x"3af0",x"39c3",x"359e",x"403a",x"36da",x"b925",x"ba1f",x"0000",x"3af0",x"39bd",x"35bd",x"4039",x"3710",x"2c74",x"bbfb",x"0000",x"3afb",x"39c3"),
(x"351b",x"4050",x"36da",x"3664",x"3b55",x"0000",x"3a50",x"3b4c",x"353f",x"404d",x"36da",x"3746",x"3b1f",x"0000",x"3a50",x"3b44",x"351b",x"4050",x"3710",x"350e",x"3b96",x"0000",x"3a5a",x"3b4c"),
(x"38bd",x"403d",x"36da",x"3456",x"3bb3",x"0000",x"3a72",x"3b13",x"38c9",x"403c",x"36da",x"34cb",x"3ba1",x"8000",x"3a72",x"3b0f",x"38bd",x"403d",x"3710",x"35fc",x"3b6b",x"0000",x"3a7c",x"3b13"),
(x"386d",x"4056",x"36da",x"bac4",x"3844",x"068d",x"3a88",x"3b01",x"3877",x"4058",x"36da",x"b74e",x"3b1d",x"0000",x"3a88",x"3afc",x"386d",x"4056",x"3710",x"bba8",x"34a3",x"868d",x"3a93",x"3b01"),
(x"359e",x"403a",x"36da",x"b925",x"ba1f",x"0000",x"3af0",x"39bd",x"358a",x"403d",x"36da",x"bbad",x"b481",x"068d",x"3af0",x"39b7",x"359e",x"403a",x"3710",x"b80b",x"bae7",x"0000",x"3afb",x"39bd"),
(x"3501",x"4051",x"36da",x"2d0c",x"3bf9",x"8000",x"3a50",x"3b51",x"351b",x"4050",x"36da",x"3664",x"3b55",x"0000",x"3a50",x"3b4c",x"3501",x"4051",x"3710",x"ada8",x"3bf8",x"0000",x"3a5a",x"3b51"),
(x"38c9",x"403c",x"36da",x"34cb",x"3ba1",x"8000",x"3a72",x"3b0f",x"38d4",x"403b",x"36da",x"38a8",x"3a80",x"8000",x"3a72",x"3b0b",x"38c9",x"403c",x"3710",x"3385",x"3bc6",x"0000",x"3a7c",x"3b0f"),
(x"386c",x"4053",x"36da",x"bbdd",x"b1e1",x"8000",x"3a88",x"3b05",x"386d",x"4056",x"36da",x"bac4",x"3844",x"068d",x"3a88",x"3b01",x"386c",x"4053",x"3710",x"bb38",x"b6e2",x"868d",x"3a93",x"3b05"),
(x"358a",x"403d",x"36da",x"bbad",x"b481",x"068d",x"3af0",x"39b7",x"3587",x"4040",x"36da",x"bb8b",x"3553",x"0000",x"3af0",x"39b3",x"358a",x"403d",x"3710",x"bb1e",x"b74c",x"0000",x"3afb",x"39b7"),
(x"34e9",x"4050",x"36da",x"b50d",x"3b97",x"8000",x"3a50",x"3b56",x"3501",x"4051",x"36da",x"2d0c",x"3bf9",x"8000",x"3a50",x"3b51",x"34e9",x"4050",x"3710",x"b698",x"3b49",x"0000",x"3a5a",x"3b56"),
(x"38d4",x"403b",x"36da",x"38a8",x"3a80",x"8000",x"3a72",x"3b0b",x"38d9",x"403a",x"36da",x"3bfc",x"2b03",x"0a8d",x"3a72",x"3b08",x"38d4",x"403b",x"3710",x"37f2",x"3af1",x"8000",x"3a7c",x"3b0b"),
(x"3872",x"4051",x"36da",x"b9d1",x"b97d",x"068d",x"3a88",x"3b08",x"386c",x"4053",x"36da",x"bbdd",x"b1e1",x"8000",x"3a88",x"3b05",x"3872",x"4051",x"3710",x"b902",x"ba3c",x"0000",x"3a93",x"3b08"),
(x"3587",x"4040",x"36da",x"bb8b",x"3553",x"0000",x"3af0",x"39b3",x"3593",x"4042",x"36da",x"bc00",x"95bc",x"0000",x"3af0",x"39af",x"3587",x"4040",x"3710",x"bbf7",x"2dba",x"868d",x"3afb",x"39b3"),
(x"34cb",x"404e",x"36da",x"b64c",x"3b5a",x"0000",x"3a50",x"3b5d",x"34e9",x"4050",x"36da",x"b50d",x"3b97",x"8000",x"3a50",x"3b56",x"34cb",x"404e",x"3710",x"b501",x"3b99",x"0000",x"3a5a",x"3b5d"),
(x"38d9",x"403a",x"36da",x"3bfc",x"2b03",x"0a8d",x"3a72",x"3b08",x"38d8",x"4039",x"36da",x"3b96",x"b50f",x"0000",x"3a72",x"3b07",x"38d9",x"403a",x"3710",x"3b87",x"3565",x"0000",x"3a7c",x"3b08"),
(x"3885",x"404f",x"36da",x"b7ea",x"baf3",x"8000",x"3a88",x"3b10",x"3872",x"4051",x"36da",x"b9d1",x"b97d",x"068d",x"3a88",x"3b08",x"3885",x"404f",x"3710",x"b83d",x"bac8",x"0000",x"3a93",x"3b10"),
(x"3593",x"4042",x"36da",x"bc00",x"95bc",x"0000",x"3af0",x"39af",x"3592",x"4043",x"36da",x"ba08",x"b941",x"8000",x"3af0",x"39ae",x"3593",x"4042",x"3710",x"bbda",x"321b",x"8000",x"3afb",x"39af"),
(x"34bb",x"404d",x"36da",x"b31c",x"3bcc",x"0000",x"3a50",x"3b60",x"34cb",x"404e",x"36da",x"b64c",x"3b5a",x"0000",x"3a50",x"3b5d",x"34bb",x"404d",x"3710",x"b141",x"3be4",x"0000",x"3a5a",x"3b60"),
(x"38d8",x"4039",x"36da",x"3b96",x"b50f",x"0000",x"3a72",x"3b07",x"38c7",x"4038",x"36da",x"364a",x"bb5b",x"8000",x"3a72",x"3b00",x"38d8",x"4039",x"3710",x"3be4",x"b12f",x"868d",x"3a7c",x"3b07"),
(x"388c",x"404e",x"36da",x"bb54",x"b669",x"8000",x"3a88",x"3b13",x"3885",x"404f",x"36da",x"b7ea",x"baf3",x"8000",x"3a88",x"3b10",x"388c",x"404e",x"3710",x"bbfd",x"a9ab",x"0000",x"3a93",x"3b13"),
(x"3592",x"4043",x"36da",x"ba08",x"b941",x"8000",x"3a50",x"3bb0",x"357d",x"4043",x"36da",x"26c2",x"bbff",x"0000",x"3a50",x"3bac",x"3592",x"4043",x"3710",x"bba4",x"b4bb",x"0000",x"3a5a",x"3bb0"),
(x"349b",x"404d",x"36da",x"b221",x"3bda",x"0000",x"3a50",x"3b66",x"34bb",x"404d",x"36da",x"b31c",x"3bcc",x"0000",x"3a50",x"3b60",x"349b",x"404d",x"3710",x"b4a8",x"3ba7",x"0000",x"3a5a",x"3b66"),
(x"38c7",x"4038",x"36da",x"364a",x"bb5b",x"8000",x"3a72",x"3b00",x"38b7",x"4036",x"36da",x"32f6",x"bbce",x"0000",x"3a72",x"3af9",x"38c7",x"4038",x"3710",x"3653",x"bb59",x"0000",x"3a7c",x"3b00"),
(x"388c",x"404d",x"36da",x"bb52",x"3671",x"0000",x"3a8b",x"3b19",x"388c",x"404e",x"36da",x"bb54",x"b669",x"8000",x"3a8b",x"3b18",x"388c",x"404d",x"3710",x"b967",x"39e6",x"0000",x"3a96",x"3b19"),
(x"357d",x"4043",x"36da",x"26c2",x"bbff",x"0000",x"3a50",x"3bac",x"3555",x"4043",x"36da",x"35eb",x"bb6e",x"0000",x"3a50",x"3ba5",x"357d",x"4043",x"3710",x"a8c9",x"bbfe",x"0000",x"3a5a",x"3bac"),
(x"3485",x"404c",x"36da",x"b819",x"3ade",x"8000",x"3a50",x"3b6a",x"349b",x"404d",x"36da",x"b221",x"3bda",x"0000",x"3a50",x"3b66",x"3485",x"404c",x"3710",x"b92c",x"3a1a",x"0000",x"3a5a",x"3b6a"),
(x"38b7",x"4036",x"36da",x"32f6",x"bbce",x"0000",x"3a72",x"3af9",x"3894",x"4035",x"36da",x"b036",x"bbee",x"0000",x"3a72",x"3aec",x"38b7",x"4036",x"3710",x"3528",x"bb92",x"0000",x"3a7c",x"3af9"),
(x"3885",x"404c",x"36da",x"b305",x"3bce",x"0000",x"3a8b",x"3b1c",x"388c",x"404d",x"36da",x"bb52",x"3671",x"0000",x"3a8b",x"3b19",x"3885",x"404c",x"3710",x"b25f",x"3bd7",x"8000",x"3a96",x"3b1c"),
(x"3555",x"4043",x"36da",x"35eb",x"bb6e",x"0000",x"3a50",x"3ba5",x"353f",x"4041",x"36da",x"379f",x"bb08",x"0000",x"3a50",x"3ba0",x"3555",x"4043",x"3710",x"345a",x"bbb2",x"0000",x"3a5a",x"3ba5"),
(x"3475",x"404a",x"36da",x"baeb",x"3803",x"8000",x"3a50",x"3b6f",x"3485",x"404c",x"36da",x"b819",x"3ade",x"8000",x"3a50",x"3b6a",x"3475",x"404a",x"3710",x"bbab",x"348e",x"8000",x"3a5a",x"3b6f"),
(x"3894",x"4035",x"36da",x"b036",x"bbee",x"0000",x"3a72",x"3aec",x"3877",x"4037",x"36da",x"b8aa",x"ba7f",x"868d",x"3a72",x"3ae1",x"3894",x"4035",x"3710",x"aa0a",x"bbfd",x"8000",x"3a7c",x"3aec"),
(x"3753",x"4058",x"36da",x"38fe",x"3a3f",x"8000",x"3a8b",x"3b7d",x"3760",x"4056",x"36da",x"3bfa",x"2cac",x"868d",x"3a8b",x"3b79",x"3753",x"4058",x"3710",x"37e4",x"3af5",x"8000",x"3a96",x"3b7d"),
(x"3a2f",x"404d",x"36da",x"3bfe",x"a8f0",x"0000",x"3bfb",x"39c9",x"3a2d",x"4042",x"36da",x"3bfe",x"a8f0",x"0000",x"3bea",x"39c8",x"3a2f",x"404d",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"39bf"),
(x"353f",x"4041",x"36da",x"379f",x"bb08",x"0000",x"3a50",x"3ba0",x"351b",x"403f",x"36da",x"350e",x"bb96",x"0000",x"3a50",x"3b98",x"353f",x"4041",x"3710",x"3746",x"bb1f",x"0000",x"3a5a",x"3ba0"),
(x"39f5",x"4059",x"36da",x"a49b",x"3bff",x"8000",x"3a2d",x"3b9f",x"3a27",x"4059",x"36da",x"a3ae",x"3bff",x"0000",x"3a2d",x"3bb3",x"39f5",x"4059",x"3710",x"a4e3",x"3bff",x"1818",x"3a23",x"3b9f"),
(x"3877",x"4037",x"36da",x"b8aa",x"ba7f",x"868d",x"3a72",x"3ae1",x"386d",x"4039",x"36da",x"bba8",x"b4a3",x"8000",x"3a72",x"3adc",x"3877",x"4037",x"3710",x"b74e",x"bb1d",x"8000",x"3a7c",x"3ae1"),
(x"382a",x"404d",x"36da",x"2f40",x"3bf2",x"8000",x"3a8b",x"3b3e",x"3885",x"404c",x"36da",x"b305",x"3bce",x"0000",x"3a8b",x"3b1c",x"382a",x"404d",x"3710",x"30bd",x"3be9",x"8000",x"3a96",x"3b3e"),
(x"351b",x"403f",x"36da",x"350e",x"bb96",x"0000",x"3a50",x"3b98",x"3501",x"403e",x"36da",x"ada8",x"bbf8",x"8000",x"3a50",x"3b93",x"351b",x"403f",x"3710",x"3664",x"bb55",x"0000",x"3a5a",x"3b98"),
(x"386d",x"4039",x"36da",x"bba8",x"b4a3",x"8000",x"3a72",x"3adc",x"386c",x"403c",x"36da",x"bb38",x"36e2",x"868d",x"3a72",x"3ad8",x"386d",x"4039",x"3710",x"bac4",x"b844",x"0000",x"3a7c",x"3adc"),
(x"3813",x"404e",x"36da",x"27fc",x"3bfe",x"0000",x"3a8b",x"3b47",x"382a",x"404d",x"36da",x"2f40",x"3bf2",x"8000",x"3a8b",x"3b3e",x"3813",x"404e",x"3710",x"a8bf",x"3bfe",x"8000",x"3a96",x"3b47"),
(x"3a2d",x"4042",x"36da",x"367a",x"bb50",x"0000",x"3b1f",x"387c",x"3a25",x"4041",x"36da",x"367a",x"bb50",x"0000",x"3b21",x"387e",x"3a2d",x"4042",x"3710",x"3644",x"bb4c",x"2f83",x"3b19",x"3884"),
(x"3a1f",x"3d5c",x"3733",x"3b23",x"251e",x"3737",x"3a49",x"339f",x"3a25",x"3d5c",x"3710",x"3bd6",x"2604",x"3256",x"3a49",x"33c0",x"3a20",x"3d45",x"3732",x"3b18",x"2439",x"3763",x"3a35",x"33aa"),
(x"3a18",x"3d5c",x"3748",x"36c9",x"29dc",x"3b3c",x"3a48",x"3388",x"3a1f",x"3d5c",x"3733",x"3b23",x"251e",x"3737",x"3a49",x"339f",x"3a19",x"3d45",x"3749",x"3871",x"2587",x"3aa6",x"3a35",x"3392"),
(x"3a10",x"3d5c",x"3749",x"b4de",x"2b76",x"3b9b",x"3a48",x"337b",x"3a18",x"3d5c",x"3748",x"36c9",x"29dc",x"3b3c",x"3a48",x"3388",x"3a14",x"3d45",x"374e",x"2fa2",x"2997",x"3bef",x"3a34",x"3387"),
(x"3a09",x"3d5c",x"373b",x"b9d7",x"2404",x"3976",x"3a48",x"3369",x"3a10",x"3d5c",x"3749",x"b4de",x"2b76",x"3b9b",x"3a48",x"337b",x"3a0d",x"3d45",x"374b",x"b745",x"2966",x"3b1e",x"3a34",x"337b"),
(x"3a09",x"3d5e",x"373a",x"baf6",x"2b34",x"37d2",x"3bbc",x"39cf",x"3a09",x"3d5c",x"373b",x"b7a6",x"3a67",x"35ca",x"3bbd",x"39cf",x"3a03",x"3d5d",x"370e",x"ae5c",x"3b3a",x"36a9",x"3bc0",x"39d7"),
(x"3a09",x"3d5c",x"373b",x"b7a6",x"3a67",x"35ca",x"3bbd",x"39cf",x"3a09",x"3d5e",x"373a",x"baf6",x"2b34",x"37d2",x"3bbc",x"39cf",x"3a10",x"3d5c",x"3749",x"b3aa",x"a4b5",x"3bc3",x"3bbb",x"39cb"),
(x"3a08",x"3d73",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"3978",x"3a09",x"3d5e",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"3979",x"3a04",x"3d73",x"3727",x"bbc5",x"a8fd",x"3377",x"3bfb",x"3974"),
(x"3a03",x"3d5d",x"370e",x"bbc2",x"ab4f",x"338c",x"3bea",x"3970",x"3a04",x"3d73",x"3727",x"bbc5",x"a8fd",x"3377",x"3bfb",x"3974",x"3a09",x"3d5e",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"3979"),
(x"3a09",x"3d5e",x"373a",x"ba80",x"a874",x"38a7",x"3beb",x"3979",x"3a08",x"3d73",x"373e",x"bb1c",x"a938",x"374b",x"3bfb",x"3978",x"3a11",x"3d5e",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"397d"),
(x"3a11",x"3d5e",x"374a",x"b575",x"a7e2",x"3b83",x"3beb",x"397d",x"3a0f",x"3d72",x"374d",x"b891",x"aa52",x"3a8d",x"3bfb",x"397c",x"3a19",x"3d5e",x"374d",x"3400",x"aa73",x"3bbc",x"3beb",x"3980"),
(x"3a17",x"3d72",x"3751",x"2a2e",x"aa4f",x"3bfb",x"3bfb",x"397f",x"3a1d",x"3d72",x"374d",x"3802",x"a90b",x"3aea",x"3bfb",x"3982",x"3a19",x"3d5e",x"374d",x"3400",x"aa73",x"3bbc",x"3beb",x"3980"),
(x"3a1d",x"3d72",x"374d",x"3802",x"a90b",x"3aea",x"3bfb",x"3982",x"3a24",x"3d72",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"3986",x"3a21",x"3d5e",x"3744",x"3962",x"a91e",x"39e8",x"3beb",x"3984"),
(x"3a24",x"3d72",x"373f",x"3a93",x"a694",x"388c",x"3bfb",x"3986",x"3a2a",x"3d73",x"3725",x"3b3f",x"a65f",x"36c3",x"3bfb",x"398b",x"3a25",x"3d5e",x"3738",x"3aa3",x"a5dc",x"3875",x"3beb",x"3986"),
(x"3a1f",x"3d5c",x"3733",x"37ff",x"ba99",x"3438",x"3bba",x"39c3",x"3a25",x"3d5e",x"3738",x"36f3",x"bae7",x"3422",x"3bb7",x"39c3",x"3a25",x"3d5c",x"3710",x"3700",x"bb23",x"2f05",x"3bbd",x"39bd"),
(x"3a02",x"3d45",x"3724",x"bb1f",x"1a24",x"3747",x"3a34",x"3352",x"3a09",x"3d5c",x"373b",x"b9d7",x"2404",x"3976",x"3a48",x"3369",x"3a07",x"3d45",x"373c",x"bac4",x"2853",x"3841",x"3a34",x"336a"),
(x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e",x"3a09",x"3d5c",x"373b",x"b9d7",x"2404",x"3976",x"3a48",x"3369",x"3a02",x"3d45",x"3724",x"bb1f",x"1a24",x"3747",x"3a34",x"3352"),
(x"3a10",x"3d5c",x"3749",x"b3aa",x"a4b5",x"3bc3",x"3bbb",x"39cb",x"3a11",x"3d5e",x"374a",x"b547",x"b37e",x"3b50",x"3bb9",x"39cc",x"3a18",x"3d5c",x"3748",x"291b",x"b8de",x"3a57",x"3bba",x"39c9"),
(x"3a1f",x"3d5c",x"3733",x"37ff",x"ba99",x"3438",x"3bba",x"39c3",x"3a18",x"3d5c",x"3748",x"291b",x"b8de",x"3a57",x"3bba",x"39c9",x"3a21",x"3d5e",x"3744",x"37e0",x"ba17",x"36be",x"3bb7",x"39c5"),
(x"3a2f",x"3d73",x"3710",x"32c7",x"3bca",x"2d1d",x"3b20",x"383f",x"3a2a",x"3d73",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3843",x"3a26",x"3d74",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3842"),
(x"3a2a",x"3d73",x"3725",x"3571",x"3b76",x"2f80",x"3b22",x"3843",x"3a24",x"3d72",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3848",x"3a20",x"3d74",x"3739",x"34f2",x"3b46",x"3471",x"3b22",x"3849"),
(x"3a24",x"3d72",x"373f",x"36ad",x"3af4",x"343a",x"3b24",x"3848",x"3a1d",x"3d72",x"374d",x"3561",x"3aa0",x"372c",x"3b25",x"384c",x"3a1a",x"3d74",x"3746",x"342e",x"3adb",x"3719",x"3b22",x"384d"),
(x"3a17",x"3d72",x"3751",x"2fda",x"39a6",x"3994",x"3b24",x"384f",x"3a0f",x"3d72",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3851",x"3a15",x"3d74",x"374b",x"aaa7",x"39a6",x"39a5",x"3b22",x"384f"),
(x"3a0f",x"3d72",x"374d",x"b509",x"37b0",x"3a8c",x"3b22",x"3851",x"3a08",x"3d73",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3854",x"3a0f",x"3d74",x"3749",x"b6e3",x"3562",x"3ab3",x"3b21",x"3851"),
(x"3a08",x"3d73",x"373e",x"baca",x"3414",x"3768",x"3b1f",x"3854",x"3a04",x"3d73",x"3727",x"bada",x"b46a",x"36f8",x"3b1b",x"3857",x"3a09",x"3d74",x"373e",x"ba28",x"9dd6",x"391a",x"3b1e",x"3853"),
(x"39fb",x"3d73",x"3713",x"a9a5",x"a460",x"3bfd",x"3a5b",x"333d",x"3a02",x"3d73",x"3711",x"315a",x"2bae",x"3bdf",x"3a5b",x"3349",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e"),
(x"3a20",x"3d74",x"3739",x"3abd",x"a8b5",x"384c",x"3a5c",x"339e",x"3a24",x"3d8b",x"372b",x"3b86",x"a8a8",x"3564",x"3a6f",x"33b1",x"3a26",x"3d74",x"3710",x"3bed",x"a7ae",x"3024",x"3a5b",x"33c4"),
(x"3a21",x"3d8b",x"373a",x"3acd",x"a5ae",x"3834",x"3a6f",x"33a3",x"3a20",x"3d74",x"3739",x"3abd",x"a8b5",x"384c",x"3a5c",x"339e",x"3a1a",x"3d8a",x"3749",x"38cd",x"a812",x"3a64",x"3a6f",x"3391"),
(x"3a1a",x"3d74",x"3746",x"38a5",x"a839",x"3a81",x"3a5c",x"338e",x"3a15",x"3d74",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a5c",x"3385",x"3a1a",x"3d8a",x"3749",x"38cd",x"a812",x"3a64",x"3a6f",x"3391"),
(x"3a15",x"3d74",x"374b",x"2e56",x"a8d3",x"3bf4",x"3a5c",x"3385",x"3a0f",x"3d74",x"3749",x"b771",x"a91b",x"3b13",x"3a5c",x"3379",x"3a14",x"3d8a",x"374f",x"32be",x"a89e",x"3bd0",x"3a6f",x"3385"),
(x"3a0f",x"3d74",x"3749",x"b771",x"a91b",x"3b13",x"3a5c",x"3379",x"3a09",x"3d74",x"373e",x"ba21",x"a786",x"3921",x"3a5c",x"336a",x"3a0d",x"3d8a",x"374b",x"b6cb",x"a758",x"3b3d",x"3a6f",x"3378"),
(x"3a07",x"3d8a",x"373c",x"baa0",x"a6bb",x"3879",x"3a6f",x"3366",x"3a09",x"3d74",x"373e",x"ba21",x"a786",x"3921",x"3a5c",x"336a",x"3a00",x"3d8a",x"3722",x"ba6c",x"a860",x"38c2",x"3a6f",x"334c"),
(x"3a00",x"3d8a",x"3722",x"ba6c",x"a860",x"38c2",x"3a6f",x"334c",x"3a01",x"3d74",x"371c",x"b9f4",x"a495",x"3957",x"3a5c",x"334a",x"39fc",x"3d8a",x"3718",x"b8fc",x"a86a",x"3a40",x"3a6f",x"3340"),
(x"3475",x"3d64",x"3710",x"0000",x"0000",x"3c00",x"3a4e",x"2451",x"3475",x"3d6c",x"3710",x"0000",x"0000",x"3c00",x"3a55",x"2451",x"3485",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"24c1"),
(x"3485",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"24c1",x"3485",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"24c1",x"349b",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"255f"),
(x"34bb",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2643",x"349b",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"255f",x"34bb",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2643"),
(x"34bb",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2643",x"34bb",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2643",x"34cb",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"26b3"),
(x"34cb",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"26b3",x"34cb",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"26b3",x"34e9",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"278b"),
(x"3501",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"281a",x"34e9",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"278b",x"3501",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"281a"),
(x"3501",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"281a",x"3501",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"281a",x"351b",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2878"),
(x"353f",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"28fb",x"351b",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2878",x"353f",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"28fb"),
(x"353f",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"28fb",x"353f",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"28fb",x"3555",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2949"),
(x"3555",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2949",x"3555",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2949",x"357d",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4b",x"29d7"),
(x"3592",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2a20",x"357d",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4b",x"29d7",x"3592",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2a20"),
(x"36f7",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2d8d",x"363b",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2c3f",x"36f7",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2d8d"),
(x"363b",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2c3f",x"363b",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2c3f",x"362c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2c23"),
(x"362c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"2c23",x"362c",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2c23",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"3592",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2a20",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b",x"3592",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2a20"),
(x"35e4",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2b48",x"35f5",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2b84",x"35fd",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"2ba0"),
(x"35d3",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2b0a",x"35e4",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2b48",x"35f3",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2b7d"),
(x"35bd",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2aba",x"35d3",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2b0a",x"35f1",x"3d7d",x"3710",x"868d",x"0cea",x"3c00",x"3a63",x"2b76"),
(x"35fd",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2ba0",x"35f5",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2b84",x"35fd",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2ba0"),
(x"35fd",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2ba0",x"35e4",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2b48",x"35f3",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2b7d"),
(x"35f3",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2b7d",x"35d3",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2b0a",x"35f1",x"3d53",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2b76"),
(x"35f1",x"3d53",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2b76",x"35bd",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"2aba",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b"),
(x"359e",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a68",x"2a4d",x"35bd",x"3d85",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"2aba",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"36f7",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2d8d",x"36f7",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2d8d",x"3710",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2dbb"),
(x"380a",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2f8b",x"380a",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2f8b",x"37b8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2ee7"),
(x"37b8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2ee7",x"37b8",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2ee7",x"37a8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ec9"),
(x"37a8",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ec9",x"37a8",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2ec9",x"378c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2e97"),
(x"378c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2e97",x"378c",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2e97",x"376c",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2e5e"),
(x"3752",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2e30",x"376c",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"2e5e",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"36e3",x"3d8c",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"2d6a",x"36f7",x"3d8e",x"3710",x"0000",x"0000",x"3c00",x"3a72",x"2d8e",x"36df",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"2d63"),
(x"36df",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"2d63",x"3716",x"3d8d",x"3710",x"0000",x"0000",x"3c00",x"3a72",x"2dc4",x"36dc",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2d5e"),
(x"36e3",x"3d43",x"3710",x"0000",x"0000",x"3c00",x"3a32",x"2d6a",x"36df",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"2d63",x"36f7",x"3d41",x"3710",x"0000",x"0000",x"3c00",x"3a30",x"2d8e"),
(x"36df",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"2d63",x"36dc",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2d5e",x"3716",x"3d42",x"3710",x"0000",x"0000",x"3c00",x"3a31",x"2dc4"),
(x"3760",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2e49",x"3753",x"3d46",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"2e32",x"375f",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2e47"),
(x"375f",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"2e47",x"3742",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2e14",x"3754",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"2e33"),
(x"3742",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"2e14",x"3753",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"2e32",x"375f",x"3d83",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"2e47"),
(x"372e",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"2df0",x"3742",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"2e14",x"3754",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"2e33"),
(x"3705",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5f",x"2da6",x"36cb",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2d40",x"36c4",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2d33"),
(x"36c2",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2d2f",x"36cb",x"3d56",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2d40",x"36c4",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2d33"),
(x"36c4",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2d33",x"3705",x"3d58",x"3710",x"0000",x"0000",x"3c00",x"3a44",x"2da6",x"36dc",x"3d4a",x"3710",x"0000",x"0000",x"3c00",x"3a38",x"2d5e"),
(x"3713",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2dbf",x"3705",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5f",x"2da6",x"36dc",x"3d86",x"3710",x"0000",x"0000",x"3c00",x"3a6b",x"2d5e"),
(x"3754",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"2e33",x"3713",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2dbf",x"372e",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"2df0"),
(x"3754",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"2e33",x"372e",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"2df0",x"3713",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2dbf"),
(x"3716",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2dc5",x"3713",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"2dbf",x"3752",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"2e30"),
(x"3754",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"2e33",x"3713",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a46",x"2dbf",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"3716",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2dc5",x"3710",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"2dbb",x"3716",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2dc5"),
(x"3716",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2dc5",x"3716",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2dc5",x"3752",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"2e30"),
(x"380a",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2f8b",x"380a",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2f8b",x"3813",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2fac"),
(x"3813",x"3d74",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"2fac",x"382a",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ffc",x"3813",x"3d5c",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2fac"),
(x"382a",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"2ffc",x"382a",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2ffc",x"3885",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"30a2"),
(x"3885",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"30a2",x"388c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"30ad",x"3885",x"3d5e",x"3710",x"0000",x"0000",x"3c00",x"3a49",x"30a2"),
(x"38d5",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"3130",x"38d5",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"3130",x"38bf",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"3109"),
(x"38b2",x"3d76",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"30f1",x"38bf",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"3109",x"38b2",x"3d5a",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30f1"),
(x"38b0",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"30ed",x"38b2",x"3d76",x"3710",x"0000",x"0000",x"3c00",x"3a5d",x"30f1",x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed"),
(x"38b0",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"30ed",x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed",x"388c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"30ad"),
(x"386c",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"3075",x"3872",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"3080",x"386d",x"3d4b",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"3076"),
(x"3872",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"3080",x"3885",x"3d59",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30a2",x"3877",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a35",x"3088"),
(x"386c",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"3075",x"386d",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"3076",x"3872",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"3080"),
(x"3872",x"3d7b",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"3080",x"3877",x"3d89",x"3710",x"0000",x"0000",x"3c00",x"3a6e",x"3088",x"3885",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5e",x"30a2"),
(x"3885",x"3d77",x"3710",x"0000",x"0000",x"3c00",x"3a5e",x"30a2",x"3894",x"3d8c",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"30bc",x"388c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"30ae"),
(x"3885",x"3d59",x"3710",x"0000",x"0000",x"3c00",x"3a45",x"30a2",x"388c",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"30ae",x"3894",x"3d44",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30bc"),
(x"38d9",x"3d4d",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"3136",x"38d8",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"3135",x"38d4",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3d",x"312d"),
(x"38c7",x"3d87",x"3710",x"0000",x"0000",x"3c00",x"3a6c",x"3117",x"38d8",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"3135",x"38d4",x"3d80",x"3710",x"0000",x"0000",x"3c00",x"3a66",x"312d"),
(x"38b7",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"30f9",x"38c7",x"3d87",x"3710",x"0000",x"0000",x"3c00",x"3a6c",x"3117",x"38c9",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"311a"),
(x"38d4",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3d",x"312d",x"38c7",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3117",x"38c9",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"311a"),
(x"38b2",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"30f2",x"388c",x"3d5b",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"30ae",x"38b0",x"3d57",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"30ed"),
(x"388c",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"30ad",x"388c",x"3d75",x"3710",x"0000",x"0000",x"3c00",x"3a5c",x"30ae",x"38b0",x"3d78",x"3710",x"0000",x"0000",x"3c00",x"3a60",x"30ed"),
(x"38d5",x"3d71",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"3130",x"38f6",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"316b",x"38d5",x"3d5f",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"3130"),
(x"38f6",x"3d73",x"3710",x"0000",x"0000",x"3c00",x"3a5b",x"316b",x"3915",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"31a2",x"38f6",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a48",x"316b"),
(x"3915",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"31a2",x"392f",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"31d0",x"3915",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"31a2"),
(x"392f",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"31d0",x"393f",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"31ed",x"392f",x"3d48",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"31d0"),
(x"393f",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a70",x"31ed",x"3953",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3211",x"393f",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"31ed"),
(x"3953",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3211",x"395a",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"321d",x"3953",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3211"),
(x"395a",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a6a",x"321d",x"395d",x"3d81",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"3222",x"395a",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a39",x"321d"),
(x"395d",x"3d4f",x"3710",x"0000",x"0000",x"3c00",x"3a3c",x"3222",x"395d",x"3d81",x"3710",x"0000",x"0000",x"3c00",x"3a67",x"3222",x"3963",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"322d"),
(x"3963",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"322d",x"3972",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"3248",x"3963",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"322d"),
(x"3972",x"3d7f",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"3248",x"3985",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"3269",x"3972",x"3d50",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"3248"),
(x"3985",x"3d84",x"3710",x"0000",x"0000",x"3c00",x"3a69",x"3269",x"3994",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3284",x"3985",x"3d4c",x"3710",x"0000",x"0000",x"3c00",x"3a3a",x"3269"),
(x"3994",x"3d88",x"3710",x"0000",x"0000",x"3c00",x"3a6d",x"3284",x"3999",x"3d89",x"3710",x"935f",x"1e0a",x"3c00",x"3a6e",x"328d",x"3994",x"3d47",x"3710",x"0000",x"0000",x"3c00",x"3a36",x"3284"),
(x"3999",x"3d47",x"3710",x"96f6",x"9f93",x"3c00",x"3a35",x"328d",x"3999",x"3d89",x"3710",x"935f",x"1e0a",x"3c00",x"3a6e",x"328d",x"39fc",x"3d5d",x"3713",x"ac0e",x"a310",x"3bfb",x"3a48",x"333e"),
(x"3999",x"3d89",x"3710",x"935f",x"1e0a",x"3c00",x"3a6e",x"328d",x"39f5",x"3d8a",x"3710",x"b60a",x"25b5",x"3b67",x"3a6f",x"3331",x"39fb",x"3d73",x"3713",x"a9a5",x"a460",x"3bfd",x"3a5b",x"333d"),
(x"3a14",x"3d8a",x"374f",x"a8f4",x"3bfa",x"ac28",x"3bbf",x"3a20",x"3a0d",x"3d8a",x"374b",x"a412",x"3bfd",x"2966",x"3bc0",x"3a1e",x"3a1a",x"3d8a",x"3749",x"a2b5",x"3bfe",x"2818",x"3bc0",x"3a23"),
(x"3a1a",x"3d8a",x"3749",x"a2b5",x"3bfe",x"2818",x"3bc0",x"3a23",x"3a07",x"3d8a",x"373c",x"a752",x"3bff",x"9bfc",x"3bc3",x"3a1b",x"3a21",x"3d8b",x"373a",x"a884",x"3bfe",x"2546",x"3bc3",x"3a25"),
(x"3a21",x"3d8b",x"373a",x"a884",x"3bfe",x"2546",x"3bc3",x"3a25",x"3a00",x"3d8a",x"3722",x"23fc",x"3bf8",x"2d56",x"3bc8",x"3a19",x"3a24",x"3d8b",x"372b",x"a504",x"3bff",x"9a24",x"3bc6",x"3a27"),
(x"3a24",x"3d8b",x"372b",x"a504",x"3bff",x"9a24",x"3bc6",x"3a27",x"39fc",x"3d8a",x"3718",x"135f",x"3bfd",x"29a1",x"3bc9",x"3a17",x"3a27",x"3d8b",x"3710",x"a3ef",x"3bff",x"9818",x"3bcb",x"3a28"),
(x"3a14",x"3d45",x"374e",x"a81b",x"bbe6",x"b0f3",x"3a5b",x"3a5c",x"3a19",x"3d45",x"3749",x"209b",x"bc00",x"135f",x"3a5a",x"3a5e",x"3a0d",x"3d45",x"374b",x"1481",x"bbff",x"26a7",x"3a5a",x"3a5a"),
(x"3a19",x"3d45",x"3749",x"209b",x"bc00",x"135f",x"3a5a",x"3a5e",x"3a20",x"3d45",x"3732",x"1f93",x"bc00",x"975f",x"3a55",x"3a61",x"3a07",x"3d45",x"373c",x"0a8d",x"bbfe",x"27bb",x"3a57",x"3a57"),
(x"3a20",x"3d45",x"3732",x"1f93",x"bc00",x"975f",x"3a55",x"3a61",x"3a26",x"3d45",x"3710",x"1f5f",x"bbff",x"a032",x"3a4f",x"3a63",x"3a02",x"3d45",x"3724",x"1c81",x"bbff",x"a1d6",x"3a53",x"3a55"),
(x"3501",x"3d55",x"36da",x"ada8",x"bbf8",x"8000",x"3a5f",x"3b94",x"34e9",x"3d56",x"36da",x"b698",x"bb49",x"8000",x"3a5f",x"3b8f",x"3501",x"3d55",x"3710",x"2d0c",x"bbf9",x"0000",x"3a6a",x"3b94"),
(x"386c",x"3d51",x"36da",x"bb38",x"36e2",x"068d",x"3a33",x"39d5",x"3872",x"3d54",x"36da",x"b902",x"3a3c",x"0000",x"3a33",x"39d2",x"386c",x"3d51",x"3710",x"bbdd",x"31e1",x"0000",x"3a3e",x"39d5"),
(x"380a",x"3d74",x"36da",x"ad56",x"3bf8",x"8000",x"3a3d",x"3b7d",x"3813",x"3d74",x"36da",x"27fc",x"3bfe",x"0000",x"3a3d",x"3b80",x"380a",x"3d74",x"3710",x"ae12",x"3bf6",x"0000",x"3a32",x"3b7d"),
(x"34e9",x"3d56",x"36da",x"b698",x"bb49",x"8000",x"3a5f",x"3b8f",x"34cb",x"3d5b",x"36da",x"b501",x"bb99",x"0000",x"3a5f",x"3b88",x"34e9",x"3d56",x"3710",x"b50d",x"bb97",x"0000",x"3a6a",x"3b8f"),
(x"3a26",x"3d45",x"36da",x"1e3f",x"bc00",x"0000",x"3a44",x"3a63",x"39fc",x"3d45",x"36da",x"a111",x"bc00",x"0000",x"3a44",x"3a53",x"3a26",x"3d45",x"3710",x"1f5f",x"bbff",x"a032",x"3a4f",x"3a63"),
(x"3872",x"3d54",x"36da",x"b902",x"3a3c",x"0000",x"3a33",x"39d2",x"3885",x"3d59",x"36da",x"b83d",x"3ac8",x"0000",x"3a33",x"39ca",x"3872",x"3d54",x"3710",x"b9d1",x"397d",x"8000",x"3a3e",x"39d2"),
(x"3760",x"3d86",x"36da",x"3bfa",x"2cac",x"8000",x"3a3d",x"3b4c",x"375f",x"3d83",x"36da",x"3b14",x"b774",x"068d",x"3a3d",x"3b4e",x"3760",x"3d86",x"3710",x"3b92",x"3528",x"8000",x"3a32",x"3b4c"),
(x"34cb",x"3d5b",x"36da",x"b501",x"bb99",x"0000",x"3a5f",x"3b88",x"34bb",x"3d5c",x"36da",x"b141",x"bbe4",x"0000",x"3a5f",x"3b85",x"34cb",x"3d5b",x"3710",x"b64c",x"bb5a",x"0000",x"3a6a",x"3b88"),
(x"3885",x"3d59",x"36da",x"b83d",x"3ac8",x"0000",x"3a33",x"39ca",x"388c",x"3d5b",x"36da",x"bbfd",x"29ab",x"0000",x"3a33",x"39c7",x"3885",x"3d59",x"3710",x"b7eb",x"3af3",x"0000",x"3a3e",x"39ca"),
(x"37b8",x"3d71",x"36da",x"2df5",x"3bf7",x"8000",x"3a3d",x"3b6a",x"380a",x"3d74",x"36da",x"ad56",x"3bf8",x"8000",x"3a3d",x"3b7d",x"37b8",x"3d71",x"3710",x"30d0",x"3be8",x"0000",x"3a32",x"3b6a"),
(x"34bb",x"3d5c",x"36da",x"b141",x"bbe4",x"0000",x"3a5f",x"3b85",x"349b",x"3d5d",x"36da",x"b4a8",x"bba7",x"8000",x"3a5f",x"3b7f",x"34bb",x"3d5c",x"3710",x"b31c",x"bbcc",x"0000",x"3a6a",x"3b85"),
(x"388c",x"3d5b",x"36da",x"bbfd",x"29ab",x"0000",x"3a33",x"39c7",x"388c",x"3d5d",x"36da",x"b967",x"b9e6",x"0000",x"3a33",x"39c5",x"388c",x"3d5b",x"3710",x"bb54",x"3669",x"8000",x"3a3e",x"39c7"),
(x"37a8",x"3d71",x"36da",x"33d5",x"3bc1",x"0000",x"3a3d",x"3b67",x"37b8",x"3d71",x"36da",x"2df5",x"3bf7",x"8000",x"3a3d",x"3b6a",x"37a8",x"3d71",x"3710",x"3580",x"3b83",x"0000",x"3a32",x"3b67"),
(x"349b",x"3d5d",x"36da",x"b4a8",x"bba7",x"8000",x"3a5f",x"3b7f",x"3485",x"3d5f",x"36da",x"b92c",x"ba1a",x"8000",x"3a5f",x"3b7b",x"349b",x"3d5d",x"3710",x"b221",x"bbda",x"0000",x"3a6a",x"3b7f"),
(x"388c",x"3d5d",x"36da",x"b967",x"b9e6",x"0000",x"3a0c",x"3b9c",x"3885",x"3d5e",x"36da",x"b25f",x"bbd7",x"0000",x"3a0c",x"3b9a",x"388c",x"3d5d",x"3710",x"bb52",x"b671",x"0000",x"3a17",x"3b9c"),
(x"378c",x"3d75",x"36da",x"373a",x"3b23",x"0000",x"3a3d",x"3b60",x"37a8",x"3d71",x"36da",x"33d5",x"3bc1",x"0000",x"3a3d",x"3b67",x"378c",x"3d75",x"3710",x"3688",x"3b4d",x"8000",x"3a32",x"3b60"),
(x"3a26",x"3d74",x"36da",x"3311",x"3bcd",x"0000",x"3b16",x"383b",x"3a2f",x"3d73",x"36da",x"3311",x"3bcd",x"0000",x"3b18",x"3838",x"3a26",x"3d74",x"3710",x"3397",x"3bbb",x"2e23",x"3b1e",x"3842"),
(x"3485",x"3d5f",x"36da",x"b92c",x"ba1a",x"8000",x"3a5f",x"3b7b",x"3475",x"3d64",x"36da",x"bbab",x"b48e",x"0000",x"3a5f",x"3b76",x"3485",x"3d5f",x"3710",x"b819",x"bade",x"868d",x"3a6a",x"3b7b"),
(x"3760",x"3d4a",x"36da",x"3b92",x"b528",x"0000",x"3a0c",x"3b3c",x"3753",x"3d46",x"36da",x"37e4",x"baf5",x"8000",x"3a0c",x"3b39",x"3760",x"3d4a",x"3710",x"3bfa",x"acac",x"8000",x"3a17",x"3b3c"),
(x"376c",x"3d78",x"36da",x"3787",x"3b0e",x"0000",x"3a3d",x"3b5a",x"378c",x"3d75",x"36da",x"373a",x"3b23",x"0000",x"3a3d",x"3b60",x"376c",x"3d78",x"3710",x"3899",x"3a8b",x"0000",x"3a32",x"3b5a"),
(x"3885",x"3d5e",x"36da",x"b25f",x"bbd7",x"0000",x"3a0c",x"3b9a",x"382a",x"3d5d",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b77",x"3885",x"3d5e",x"3710",x"b305",x"bbce",x"0000",x"3a17",x"3b9a"),
(x"3752",x"3d7e",x"36da",x"3be0",x"31a3",x"8000",x"3a3d",x"3b53",x"376c",x"3d78",x"36da",x"3787",x"3b0e",x"0000",x"3a3d",x"3b5a",x"3752",x"3d7e",x"3710",x"3bfd",x"aabe",x"0000",x"3a32",x"3b53"),
(x"39fc",x"3d45",x"36da",x"a111",x"bc00",x"0000",x"3a44",x"3a53",x"3999",x"3d47",x"36da",x"b32b",x"bbcb",x"0000",x"3a44",x"3a2e",x"39fc",x"3d45",x"3710",x"9bc8",x"bc00",x"200b",x"3a4f",x"3a53"),
(x"382a",x"3d5d",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b77",x"3813",x"3d5c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a0c",x"3b6e",x"382a",x"3d5d",x"3710",x"2f41",x"bbf2",x"0000",x"3a17",x"3b77"),
(x"3742",x"3d8b",x"36da",x"342c",x"3bb9",x"8000",x"3a3d",x"3b44",x"3753",x"3d89",x"36da",x"38fe",x"3a3f",x"8000",x"3a3d",x"3b48",x"3742",x"3d8b",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b44"),
(x"3813",x"3d5c",x"36da",x"a8bf",x"bbfe",x"8000",x"3a0c",x"3b6e",x"380a",x"3d5c",x"36da",x"ae12",x"bbf6",x"0000",x"3a0c",x"3b6b",x"3813",x"3d5c",x"3710",x"27fc",x"bbfe",x"0000",x"3a17",x"3b6e"),
(x"372e",x"3d8b",x"36da",x"2fc6",x"3bf0",x"0000",x"3a3d",x"3b40",x"3742",x"3d8b",x"36da",x"342c",x"3bb9",x"8000",x"3a3d",x"3b44",x"372e",x"3d8b",x"3710",x"338a",x"3bc6",x"0000",x"3a32",x"3b40"),
(x"375f",x"3d4c",x"36da",x"3bc1",x"33d7",x"068d",x"3a0c",x"3b3e",x"3760",x"3d4a",x"36da",x"3b92",x"b528",x"0000",x"3a0c",x"3b3c",x"375f",x"3d4c",x"3710",x"3b14",x"3774",x"8000",x"3a17",x"3b3e"),
(x"3716",x"3d8d",x"36da",x"34b5",x"3ba5",x"8000",x"3a3d",x"3b3b",x"372e",x"3d8b",x"36da",x"2fc6",x"3bf0",x"0000",x"3a3d",x"3b40",x"3716",x"3d8d",x"3710",x"32c2",x"3bd1",x"8000",x"3a32",x"3b3b"),
(x"380a",x"3d5c",x"36da",x"ae12",x"bbf6",x"0000",x"3a0c",x"3b6b",x"37b8",x"3d5f",x"36da",x"30d0",x"bbe8",x"0000",x"3a0c",x"3b59",x"380a",x"3d5c",x"3710",x"ad54",x"bbf8",x"0000",x"3a17",x"3b6b"),
(x"36f7",x"3d8e",x"36da",x"ae6b",x"3bf5",x"0000",x"3a3d",x"3b35",x"3716",x"3d8d",x"36da",x"34b5",x"3ba5",x"8000",x"3a3d",x"3b3b",x"36f7",x"3d8e",x"3710",x"b463",x"3bb1",x"8000",x"3a32",x"3b35"),
(x"37b8",x"3d5f",x"36da",x"30d0",x"bbe8",x"0000",x"3a0c",x"3b59",x"37a8",x"3d5e",x"36da",x"3580",x"bb83",x"0000",x"3a0c",x"3b56",x"37b8",x"3d5f",x"3710",x"2df5",x"bbf7",x"0000",x"3a17",x"3b59"),
(x"36e3",x"3d8c",x"36da",x"b9b5",x"399a",x"0000",x"3a3d",x"3b31",x"36f7",x"3d8e",x"36da",x"ae6b",x"3bf5",x"0000",x"3a3d",x"3b35",x"36e3",x"3d8c",x"3710",x"bb17",x"3766",x"0000",x"3a32",x"3b31"),
(x"37a8",x"3d5e",x"36da",x"3580",x"bb83",x"0000",x"3a0c",x"3b56",x"378c",x"3d5a",x"36da",x"3688",x"bb4d",x"8000",x"3a0c",x"3b50",x"37a8",x"3d5e",x"3710",x"33d5",x"bbc1",x"0000",x"3a17",x"3b56"),
(x"36df",x"3d89",x"36da",x"bbbc",x"3412",x"0000",x"3a3d",x"3b2e",x"36e3",x"3d8c",x"36da",x"b9b5",x"399a",x"0000",x"3a3d",x"3b31",x"36df",x"3d89",x"3710",x"bbc6",x"338f",x"8000",x"3a32",x"3b2e"),
(x"378c",x"3d5a",x"36da",x"3688",x"bb4d",x"8000",x"3a0c",x"3b50",x"376c",x"3d57",x"36da",x"3899",x"ba8b",x"0000",x"3a0c",x"3b4a",x"378c",x"3d5a",x"3710",x"373a",x"bb23",x"0000",x"3a17",x"3b50"),
(x"36dc",x"3d86",x"36da",x"bba4",x"34ba",x"0000",x"3a3d",x"3b2c",x"36df",x"3d89",x"36da",x"bbbc",x"3412",x"0000",x"3a3d",x"3b2e",x"36dc",x"3d86",x"3710",x"bb3a",x"36d9",x"0000",x"3a32",x"3b2c"),
(x"3a27",x"3d8b",x"36da",x"3bff",x"a4d0",x"0000",x"3a6e",x"33f9",x"3a26",x"3d74",x"36da",x"3bff",x"a4d0",x"0000",x"3a5a",x"33f3",x"3a27",x"3d8b",x"3710",x"3bea",x"a4d6",x"30a2",x"3a6f",x"33c9"),
(x"3999",x"3d89",x"36da",x"b2b0",x"3bd2",x"0000",x"3bd5",x"39f0",x"39f5",x"3d8a",x"36da",x"a49b",x"3bff",x"8000",x"3bd5",x"3a14",x"3999",x"3d89",x"3710",x"b329",x"3bcb",x"8000",x"3bcb",x"39f0"),
(x"376c",x"3d57",x"36da",x"3899",x"ba8b",x"0000",x"3a0c",x"3b4a",x"3752",x"3d51",x"36da",x"3bfd",x"2ac2",x"0000",x"3a0c",x"3b43",x"376c",x"3d57",x"3710",x"3787",x"bb0e",x"0000",x"3a17",x"3b4a"),
(x"36c4",x"3d7f",x"36da",x"bb61",x"362a",x"0000",x"3a3d",x"3b25",x"36dc",x"3d86",x"36da",x"bba4",x"34ba",x"0000",x"3a3d",x"3b2c",x"36c4",x"3d7f",x"3710",x"bbc5",x"339b",x"0000",x"3a32",x"3b25"),
(x"3994",x"3d88",x"36da",x"b458",x"3bb2",x"8000",x"3bd5",x"39ee",x"3999",x"3d89",x"36da",x"b2b0",x"3bd2",x"0000",x"3bd5",x"39f0",x"3994",x"3d88",x"3710",x"b59f",x"3b7d",x"0000",x"3bcb",x"39ee"),
(x"3753",x"3d46",x"36da",x"37e4",x"baf5",x"8000",x"3a0c",x"3b39",x"3742",x"3d45",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b35",x"3753",x"3d46",x"3710",x"38fe",x"ba3f",x"0000",x"3a17",x"3b39"),
(x"36c2",x"3d7c",x"36da",x"bbe7",x"b0ec",x"0000",x"3a3d",x"3b22",x"36c4",x"3d7f",x"36da",x"bb61",x"362a",x"0000",x"3a3d",x"3b25",x"36c2",x"3d7c",x"3710",x"bafe",x"b7c2",x"868d",x"3a32",x"3b22"),
(x"3985",x"3d84",x"36da",x"b817",x"3adf",x"0000",x"3bd5",x"39e7",x"3994",x"3d88",x"36da",x"b458",x"3bb2",x"8000",x"3bd5",x"39ee",x"3985",x"3d84",x"3710",x"b796",x"3b0b",x"0000",x"3bcb",x"39e7"),
(x"3742",x"3d45",x"36da",x"30bd",x"bbe9",x"0000",x"3a0c",x"3b35",x"372e",x"3d45",x"36da",x"338a",x"bbc6",x"0000",x"3a0c",x"3b31",x"3742",x"3d45",x"3710",x"342c",x"bbb9",x"0000",x"3a17",x"3b35"),
(x"36cb",x"3d7a",x"36da",x"b922",x"ba22",x"868d",x"3a3d",x"3b20",x"36c2",x"3d7c",x"36da",x"bbe7",x"b0ec",x"0000",x"3a3d",x"3b22",x"36cb",x"3d7a",x"3710",x"b86c",x"baaa",x"0000",x"3a32",x"3b20"),
(x"3972",x"3d7f",x"36da",x"b475",x"3bae",x"0000",x"3bd5",x"39df",x"3985",x"3d84",x"36da",x"b817",x"3adf",x"0000",x"3bd5",x"39e7",x"3972",x"3d7f",x"3710",x"b0a0",x"3bea",x"0000",x"3bcb",x"39df"),
(x"372e",x"3d45",x"36da",x"338a",x"bbc6",x"0000",x"3a0c",x"3b31",x"3716",x"3d42",x"36da",x"32c2",x"bbd1",x"0000",x"3a0c",x"3b2c",x"372e",x"3d45",x"3710",x"2fc6",x"bbf0",x"0000",x"3a17",x"3b31"),
(x"3705",x"3d77",x"36da",x"b59a",x"bb7e",x"0000",x"3a3d",x"3b14",x"36cb",x"3d7a",x"36da",x"b922",x"ba22",x"868d",x"3a3d",x"3b20",x"3705",x"3d77",x"3710",x"b675",x"bb51",x"0000",x"3a32",x"3b14"),
(x"3963",x"3d7f",x"36da",x"3420",x"3bba",x"0000",x"3bd5",x"39d8",x"3972",x"3d7f",x"36da",x"b475",x"3bae",x"0000",x"3bd5",x"39df",x"3963",x"3d7f",x"3710",x"36c5",x"3b3f",x"0000",x"3bcb",x"39d8"),
(x"3716",x"3d42",x"36da",x"32c2",x"bbd1",x"0000",x"3a0c",x"3b2c",x"36f7",x"3d41",x"36da",x"b463",x"bbb1",x"8000",x"3a0c",x"3b27",x"3716",x"3d42",x"3710",x"34b5",x"bba5",x"0000",x"3a17",x"3b2c"),
(x"3713",x"3d75",x"36da",x"b972",x"b9db",x"8000",x"3a3d",x"3b11",x"3705",x"3d77",x"36da",x"b59a",x"bb7e",x"0000",x"3a3d",x"3b14",x"3713",x"3d75",x"3710",x"ba37",x"b909",x"0000",x"3a32",x"3b11"),
(x"395d",x"3d81",x"36da",x"399d",x"39b2",x"0000",x"3bd5",x"39d5",x"3963",x"3d7f",x"36da",x"3420",x"3bba",x"0000",x"3bd5",x"39d8",x"395d",x"3d81",x"3710",x"3ac1",x"3849",x"0000",x"3bcb",x"39d5"),
(x"36f7",x"3d41",x"36da",x"b463",x"bbb1",x"8000",x"3a0c",x"3b27",x"36e3",x"3d43",x"36da",x"bb17",x"b766",x"8000",x"3a0c",x"3b22",x"36f7",x"3d41",x"3710",x"ae6b",x"bbf5",x"0000",x"3a17",x"3b27"),
(x"3716",x"3d74",x"36da",x"bbb8",x"b42d",x"0000",x"3a3d",x"3b10",x"3713",x"3d75",x"36da",x"b972",x"b9db",x"8000",x"3a3d",x"3b11",x"3716",x"3d74",x"3710",x"bbad",x"3480",x"0000",x"3a32",x"3b10"),
(x"395a",x"3d84",x"36da",x"3b46",x"36a7",x"8000",x"3bd5",x"39d3",x"395d",x"3d81",x"36da",x"399d",x"39b2",x"0000",x"3bd5",x"39d5",x"395a",x"3d84",x"3710",x"3af1",x"37f3",x"0000",x"3bcb",x"39d3"),
(x"36e3",x"3d43",x"36da",x"bb17",x"b766",x"8000",x"3a0c",x"3b22",x"36df",x"3d47",x"36da",x"bbc6",x"b38f",x"8000",x"3a0c",x"3b20",x"36e3",x"3d43",x"3710",x"b9b5",x"b99a",x"868d",x"3a17",x"3b22"),
(x"3710",x"3d73",x"36da",x"b8f7",x"3a45",x"0000",x"3b06",x"39af",x"3716",x"3d74",x"36da",x"bbb8",x"b42d",x"0000",x"3b06",x"39ae",x"3710",x"3d73",x"3710",x"b80d",x"3ae5",x"0000",x"3b11",x"39af"),
(x"3953",x"3d88",x"36da",x"39a8",x"39a7",x"868d",x"3bd5",x"39ce",x"395a",x"3d84",x"36da",x"3b46",x"36a7",x"8000",x"3bd5",x"39d3",x"3953",x"3d88",x"3710",x"3857",x"3ab8",x"8000",x"3bcb",x"39ce"),
(x"36df",x"3d47",x"36da",x"bbc6",x"b38f",x"8000",x"3a0c",x"3b20",x"36dc",x"3d4a",x"36da",x"bb3a",x"b6d9",x"0000",x"3a0c",x"3b1d",x"36df",x"3d47",x"3710",x"bbbc",x"b412",x"0000",x"3a17",x"3b20"),
(x"36f7",x"3d72",x"36da",x"b12d",x"3be4",x"0000",x"3b06",x"39b4",x"3710",x"3d73",x"36da",x"b8f7",x"3a45",x"0000",x"3b06",x"39af",x"36f7",x"3d72",x"3710",x"b05b",x"3bec",x"8000",x"3b11",x"39b4"),
(x"3475",x"3d64",x"36da",x"bbab",x"b48e",x"0000",x"3a5f",x"3b76",x"3475",x"3d6c",x"36da",x"baeb",x"3803",x"868d",x"3a5f",x"3b70",x"3475",x"3d64",x"3710",x"baeb",x"b803",x"068d",x"3a6a",x"3b76"),
(x"393f",x"3d8b",x"36da",x"1cea",x"3c00",x"0000",x"3bd5",x"39c6",x"3953",x"3d88",x"36da",x"39a8",x"39a7",x"868d",x"3bd5",x"39ce",x"393f",x"3d8b",x"3710",x"b2bb",x"3bd2",x"868d",x"3bcb",x"39c6"),
(x"36dc",x"3d4a",x"36da",x"bb3a",x"b6d9",x"0000",x"3a0c",x"3b1d",x"36c4",x"3d51",x"36da",x"bbc5",x"b39b",x"0000",x"3a0c",x"3b17",x"36dc",x"3d4a",x"3710",x"bba4",x"b4ba",x"0000",x"3a17",x"3b1d"),
(x"362c",x"3d73",x"36da",x"3550",x"3b8b",x"0000",x"3b06",x"39db",x"363b",x"3d72",x"36da",x"3439",x"3bb7",x"0000",x"3b06",x"39d8",x"362c",x"3d73",x"3710",x"3609",x"3b68",x"8000",x"3b11",x"39db"),
(x"3999",x"3d47",x"36da",x"b32b",x"bbcb",x"0000",x"3a44",x"3a2e",x"3994",x"3d47",x"36da",x"b59f",x"bb7d",x"0000",x"3a44",x"3a2c",x"3999",x"3d47",x"3710",x"b2ba",x"bbd2",x"0000",x"3a4f",x"3a2e"),
(x"392f",x"3d88",x"36da",x"b73b",x"3b22",x"8000",x"3bd5",x"39bf",x"393f",x"3d8b",x"36da",x"1cea",x"3c00",x"0000",x"3bd5",x"39c6",x"392f",x"3d88",x"3710",x"b874",x"3aa4",x"0000",x"3bcb",x"39bf"),
(x"36c4",x"3d51",x"36da",x"bbc5",x"b39b",x"0000",x"3a0c",x"3b17",x"36c2",x"3d54",x"36da",x"baff",x"37c2",x"068d",x"3a0c",x"3b14",x"36c4",x"3d51",x"3710",x"bb61",x"b62a",x"0000",x"3a17",x"3b17"),
(x"363b",x"3d72",x"36da",x"3439",x"3bb7",x"0000",x"3b06",x"39d8",x"36f7",x"3d72",x"36da",x"b12d",x"3be4",x"0000",x"3b06",x"39b4",x"363b",x"3d72",x"3710",x"34bd",x"3ba4",x"0000",x"3b11",x"39d8"),
(x"3994",x"3d47",x"36da",x"b59f",x"bb7d",x"0000",x"3a44",x"3a2c",x"3985",x"3d4c",x"36da",x"b796",x"bb0b",x"0000",x"3a44",x"3a25",x"3994",x"3d47",x"3710",x"b458",x"bbb2",x"8000",x"3a4f",x"3a2c"),
(x"3754",x"3d80",x"36da",x"3ba5",x"b4b4",x"0000",x"3a3d",x"3b51",x"3752",x"3d7e",x"36da",x"3be0",x"31a3",x"8000",x"3a3d",x"3b53",x"3754",x"3d80",x"3710",x"3afe",x"b7c4",x"0000",x"3a32",x"3b51"),
(x"36c2",x"3d54",x"36da",x"baff",x"37c2",x"068d",x"3a0c",x"3b14",x"36cb",x"3d56",x"36da",x"b86c",x"3aa9",x"0000",x"3a0c",x"3b12",x"36c2",x"3d54",x"3710",x"bbe7",x"30ec",x"868d",x"3a17",x"3b14"),
(x"35f7",x"3d7a",x"36da",x"3a05",x"3944",x"868d",x"3b06",x"39e6",x"362c",x"3d73",x"36da",x"3550",x"3b8b",x"0000",x"3b06",x"39db",x"35f7",x"3d7a",x"3710",x"3a6a",x"38c7",x"0000",x"3b11",x"39e6"),
(x"3985",x"3d4c",x"36da",x"b796",x"bb0b",x"0000",x"3a44",x"3a25",x"3972",x"3d50",x"36da",x"b0a0",x"bbea",x"0000",x"3a44",x"3a1d",x"3985",x"3d4c",x"3710",x"b817",x"badf",x"0000",x"3a4f",x"3a25"),
(x"3915",x"3d7a",x"36da",x"b90a",x"3a36",x"0000",x"3bd5",x"39b0",x"392f",x"3d88",x"36da",x"b73b",x"3b22",x"8000",x"3bd5",x"39bf",x"3915",x"3d7a",x"3710",x"b845",x"3ac3",x"0000",x"3bcb",x"39b0"),
(x"36cb",x"3d56",x"36da",x"b86c",x"3aa9",x"0000",x"3a0c",x"3b12",x"3705",x"3d58",x"36da",x"b675",x"3b51",x"0000",x"3a0c",x"3b07",x"36cb",x"3d56",x"3710",x"b922",x"3a22",x"0000",x"3a17",x"3b12"),
(x"35f1",x"3d7d",x"36da",x"3bcd",x"3318",x"0000",x"3b06",x"39e8",x"35f7",x"3d7a",x"36da",x"3a05",x"3944",x"868d",x"3b06",x"39e6",x"35f1",x"3d7d",x"3710",x"3bf9",x"ad20",x"0000",x"3b11",x"39e8"),
(x"3972",x"3d50",x"36da",x"b0a0",x"bbea",x"0000",x"3a44",x"3a1d",x"3963",x"3d51",x"36da",x"36c5",x"bb3f",x"0000",x"3a44",x"3a17",x"3972",x"3d50",x"3710",x"b475",x"bbae",x"0000",x"3a4f",x"3a1d"),
(x"375f",x"3d83",x"36da",x"3b14",x"b774",x"068d",x"3a3d",x"3b4e",x"3754",x"3d80",x"36da",x"3ba5",x"b4b4",x"0000",x"3a3d",x"3b51",x"375f",x"3d83",x"3710",x"3bc1",x"b3d7",x"868d",x"3a32",x"3b4e"),
(x"3705",x"3d58",x"36da",x"b675",x"3b51",x"0000",x"3a0c",x"3b07",x"3713",x"3d5a",x"36da",x"ba37",x"3909",x"0000",x"3a0c",x"3b04",x"3705",x"3d58",x"3710",x"b599",x"3b7e",x"0000",x"3a17",x"3b07"),
(x"35f3",x"3d7e",x"36da",x"3b84",x"b57a",x"0000",x"3b06",x"39e9",x"35f1",x"3d7d",x"36da",x"3bcd",x"3318",x"0000",x"3b06",x"39e8",x"35f3",x"3d7e",x"3710",x"3b36",x"b6ea",x"8000",x"3b11",x"39e9"),
(x"3963",x"3d51",x"36da",x"36c5",x"bb3f",x"0000",x"3a44",x"3a17",x"395d",x"3d4f",x"36da",x"3ac1",x"b849",x"0000",x"3a44",x"3a15",x"3963",x"3d51",x"3710",x"3420",x"bbba",x"0000",x"3a4f",x"3a17"),
(x"38f6",x"3d73",x"36da",x"b551",x"3b8b",x"0000",x"3bd5",x"39a3",x"3915",x"3d7a",x"36da",x"b90a",x"3a36",x"0000",x"3bd5",x"39b0",x"38f6",x"3d73",x"3710",x"b324",x"3bcc",x"0000",x"3bcb",x"39a3"),
(x"3713",x"3d5a",x"36da",x"ba37",x"3909",x"0000",x"3a0c",x"3b04",x"3716",x"3d5b",x"36da",x"bbad",x"b480",x"0000",x"3a0c",x"3b03",x"3713",x"3d5a",x"3710",x"b972",x"39db",x"0000",x"3a17",x"3b04"),
(x"35fd",x"3d82",x"36da",x"3b91",x"b530",x"0000",x"3b06",x"39ed",x"35f3",x"3d7e",x"36da",x"3b84",x"b57a",x"0000",x"3b06",x"39e9",x"35fd",x"3d82",x"3710",x"3bf0",x"aff6",x"868d",x"3b11",x"39ed"),
(x"395d",x"3d4f",x"36da",x"3ac1",x"b849",x"0000",x"3a44",x"3a15",x"395a",x"3d4c",x"36da",x"3af1",x"b7f2",x"8000",x"3a44",x"3a12",x"395d",x"3d4f",x"3710",x"399d",x"b9b2",x"0000",x"3a4f",x"3a15"),
(x"38d5",x"3d71",x"36da",x"1953",x"3c00",x"0000",x"3bd5",x"3996",x"38f6",x"3d73",x"36da",x"b551",x"3b8b",x"0000",x"3bd5",x"39a3",x"38d5",x"3d71",x"3710",x"2dde",x"3bf7",x"0000",x"3bcb",x"3996"),
(x"3716",x"3d5b",x"36da",x"bbad",x"b480",x"0000",x"3a18",x"3a1b",x"3710",x"3d5d",x"36da",x"b80d",x"bae5",x"8000",x"3a18",x"3a1a",x"3716",x"3d5b",x"3710",x"bbb8",x"342d",x"0000",x"3a23",x"3a1b"),
(x"35fd",x"3d84",x"36da",x"3b87",x"3567",x"868d",x"3b06",x"39ee",x"35fd",x"3d82",x"36da",x"3b91",x"b530",x"0000",x"3b06",x"39ed",x"35fd",x"3d84",x"3710",x"3a08",x"3941",x"068d",x"3b11",x"39ee"),
(x"395a",x"3d4c",x"36da",x"3af1",x"b7f2",x"8000",x"3a44",x"3a12",x"3953",x"3d47",x"36da",x"3857",x"bab8",x"8000",x"3a44",x"3a0e",x"395a",x"3d4c",x"3710",x"3b46",x"b6a7",x"8000",x"3a4f",x"3a12"),
(x"38bf",x"3d73",x"36da",x"3489",x"3bab",x"0000",x"3bd5",x"398d",x"38d5",x"3d71",x"36da",x"1953",x"3c00",x"0000",x"3bd5",x"3996",x"38bf",x"3d73",x"3710",x"35f3",x"3b6c",x"0000",x"3bcb",x"398d"),
(x"3710",x"3d5d",x"36da",x"b80d",x"bae5",x"8000",x"3a18",x"3a1a",x"36f7",x"3d5e",x"36da",x"b05b",x"bbec",x"8000",x"3a18",x"3a15",x"3710",x"3d5d",x"3710",x"b8f7",x"ba45",x"0000",x"3a23",x"3a1a"),
(x"35f5",x"3d85",x"36da",x"364b",x"3b5a",x"068d",x"3b06",x"39f0",x"35fd",x"3d84",x"36da",x"3b87",x"3567",x"868d",x"3b06",x"39ee",x"35f5",x"3d85",x"3710",x"32d5",x"3bd0",x"0000",x"3b11",x"39f0"),
(x"3953",x"3d47",x"36da",x"3857",x"bab8",x"8000",x"3a44",x"3a0e",x"393f",x"3d45",x"36da",x"b2bb",x"bbd2",x"8000",x"3a44",x"3a06",x"3953",x"3d47",x"3710",x"39a8",x"b9a7",x"068d",x"3a4f",x"3a0e"),
(x"38b2",x"3d76",x"36da",x"3a0a",x"393e",x"8000",x"3bd5",x"3987",x"38bf",x"3d73",x"36da",x"3489",x"3bab",x"0000",x"3bd5",x"398d",x"38b2",x"3d76",x"3710",x"3af2",x"37f0",x"0000",x"3bcb",x"3987"),
(x"363b",x"3d5e",x"36da",x"34bd",x"bba4",x"0000",x"3a18",x"39f1",x"362c",x"3d5d",x"36da",x"3609",x"bb68",x"0000",x"3a18",x"39ee",x"363b",x"3d5e",x"3710",x"3439",x"bbb7",x"868d",x"3a23",x"39f1"),
(x"35e4",x"3d85",x"36da",x"b0fa",x"3be7",x"8000",x"3b06",x"39f3",x"35f5",x"3d85",x"36da",x"364b",x"3b5a",x"068d",x"3b06",x"39f0",x"35e4",x"3d85",x"3710",x"b3c3",x"3bc2",x"0000",x"3b11",x"39f3"),
(x"393f",x"3d45",x"36da",x"b2bb",x"bbd2",x"8000",x"3a44",x"3a06",x"392f",x"3d48",x"36da",x"b874",x"baa4",x"0000",x"3a44",x"39ff",x"393f",x"3d45",x"3710",x"1cea",x"bc00",x"8000",x"3a4f",x"3a06"),
(x"38b0",x"3d78",x"36da",x"3bfc",x"2b27",x"0000",x"3bd5",x"3985",x"38b2",x"3d76",x"36da",x"3a0a",x"393e",x"8000",x"3bd5",x"3987",x"38b0",x"3d78",x"3710",x"3ba6",x"b4ac",x"0000",x"3bcb",x"3985"),
(x"36f7",x"3d5e",x"36da",x"b05b",x"bbec",x"8000",x"3a18",x"3a15",x"363b",x"3d5e",x"36da",x"34bd",x"bba4",x"0000",x"3a18",x"39f1",x"36f7",x"3d5e",x"3710",x"b12d",x"bbe4",x"0000",x"3a23",x"3a15"),
(x"35d3",x"3d83",x"36da",x"b1d2",x"3bdd",x"0000",x"3b06",x"39f7",x"35e4",x"3d85",x"36da",x"b0fa",x"3be7",x"8000",x"3b06",x"39f3",x"35d3",x"3d83",x"3710",x"1c81",x"3c00",x"0000",x"3b11",x"39f7"),
(x"3752",x"3d51",x"36da",x"3bfd",x"2ac2",x"0000",x"3a0c",x"3b43",x"3754",x"3d4f",x"36da",x"3afe",x"37c4",x"0000",x"3a0c",x"3b41",x"3752",x"3d51",x"3710",x"3be0",x"b1a3",x"868d",x"3a17",x"3b43"),
(x"38b2",x"3d7a",x"36da",x"3a58",x"b8de",x"0000",x"3bd5",x"3983",x"38b0",x"3d78",x"36da",x"3bfc",x"2b27",x"0000",x"3bd5",x"3985",x"38b2",x"3d7a",x"3710",x"399c",x"b9b3",x"0000",x"3bcb",x"3983"),
(x"362c",x"3d5d",x"36da",x"3609",x"bb68",x"0000",x"3a18",x"39ee",x"35f7",x"3d55",x"36da",x"3a6a",x"b8c7",x"0000",x"3a18",x"39e3",x"362c",x"3d5d",x"3710",x"3550",x"bb8b",x"0000",x"3a23",x"39ee"),
(x"35bd",x"3d85",x"36da",x"2c75",x"3bfb",x"868d",x"3b06",x"39fb",x"35d3",x"3d83",x"36da",x"b1d2",x"3bdd",x"0000",x"3b06",x"39f7",x"35bd",x"3d85",x"3710",x"afcb",x"3bf0",x"8000",x"3b11",x"39fb"),
(x"392f",x"3d48",x"36da",x"b874",x"baa4",x"0000",x"3a44",x"39ff",x"3915",x"3d55",x"36da",x"b845",x"bac3",x"0000",x"3a44",x"39f1",x"392f",x"3d48",x"3710",x"b73b",x"bb22",x"0000",x"3a4f",x"39ff"),
(x"38bd",x"3d7d",x"36da",x"35fc",x"bb6b",x"0000",x"3a93",x"3ac9",x"38b2",x"3d7a",x"36da",x"3a58",x"b8de",x"0000",x"3a93",x"3ac5",x"38bd",x"3d7d",x"3710",x"3456",x"bbb3",x"0000",x"3a9e",x"3ac9"),
(x"35f7",x"3d55",x"36da",x"3a6a",x"b8c7",x"0000",x"3a18",x"39e3",x"35f1",x"3d53",x"36da",x"3bf9",x"2d21",x"0000",x"3a18",x"39e1",x"35f7",x"3d55",x"3710",x"3a05",x"b944",x"0000",x"3a23",x"39e3"),
(x"359e",x"3d82",x"36da",x"b80b",x"3ae7",x"8000",x"3b06",x"3a01",x"35bd",x"3d85",x"36da",x"2c75",x"3bfb",x"868d",x"3b06",x"39fb",x"359e",x"3d82",x"3710",x"b925",x"3a1f",x"0000",x"3b11",x"3a01"),
(x"3754",x"3d4f",x"36da",x"3afe",x"37c4",x"0000",x"3a0c",x"3b41",x"375f",x"3d4c",x"36da",x"3bc1",x"33d7",x"068d",x"3a0c",x"3b3e",x"3754",x"3d4f",x"3710",x"3ba5",x"34b5",x"0000",x"3a17",x"3b41"),
(x"38c9",x"3d7e",x"36da",x"3385",x"bbc6",x"0000",x"3a93",x"3ace",x"38bd",x"3d7d",x"36da",x"35fc",x"bb6b",x"0000",x"3a93",x"3ac9",x"38c9",x"3d7e",x"3710",x"34cb",x"bba1",x"0000",x"3a9e",x"3ace"),
(x"35f1",x"3d53",x"36da",x"3bf9",x"2d21",x"0000",x"3a18",x"39e1",x"35f3",x"3d51",x"36da",x"3b36",x"36ea",x"8000",x"3a18",x"39e0",x"35f1",x"3d53",x"3710",x"3bcd",x"b318",x"0000",x"3a23",x"39e1"),
(x"358a",x"3d7c",x"36da",x"bb1e",x"374c",x"8000",x"3b06",x"3a07",x"359e",x"3d82",x"36da",x"b80b",x"3ae7",x"8000",x"3b06",x"3a01",x"358a",x"3d7c",x"3710",x"bbad",x"3481",x"068d",x"3b11",x"3a07"),
(x"3915",x"3d55",x"36da",x"b845",x"bac3",x"0000",x"3a44",x"39f1",x"38f6",x"3d5d",x"36da",x"b324",x"bbcc",x"0000",x"3a44",x"39e4",x"3915",x"3d55",x"3710",x"b90a",x"ba36",x"0000",x"3a4f",x"39f1"),
(x"38d4",x"3d80",x"36da",x"37f2",x"baf1",x"8000",x"3a93",x"3ad2",x"38c9",x"3d7e",x"36da",x"3385",x"bbc6",x"0000",x"3a93",x"3ace",x"38d4",x"3d80",x"3710",x"38a8",x"ba80",x"8000",x"3a9e",x"3ad2"),
(x"35f3",x"3d51",x"36da",x"3b36",x"36ea",x"8000",x"3a18",x"39e0",x"35fd",x"3d4e",x"36da",x"3bf0",x"2ff4",x"8000",x"3a18",x"39dc",x"35f3",x"3d51",x"3710",x"3b84",x"357a",x"0000",x"3a23",x"39e0"),
(x"3587",x"3d77",x"36da",x"bbf7",x"adba",x"8000",x"3b06",x"3a0b",x"358a",x"3d7c",x"36da",x"bb1e",x"374c",x"8000",x"3b06",x"3a07",x"3587",x"3d77",x"3710",x"bb8b",x"b553",x"0000",x"3b11",x"3a0b"),
(x"38f6",x"3d5d",x"36da",x"b324",x"bbcc",x"0000",x"3a44",x"39e4",x"38d5",x"3d5f",x"36da",x"2dde",x"bbf7",x"0000",x"3a44",x"39d8",x"38f6",x"3d5d",x"3710",x"b551",x"bb8b",x"0000",x"3a4f",x"39e4"),
(x"38d9",x"3d82",x"36da",x"3b88",x"b564",x"0000",x"3a93",x"3ad5",x"38d4",x"3d80",x"36da",x"37f2",x"baf1",x"8000",x"3a93",x"3ad2",x"38d9",x"3d82",x"3710",x"3bfc",x"ab00",x"0000",x"3a9e",x"3ad5"),
(x"3a25",x"3d5c",x"36da",x"3bff",x"26b5",x"0000",x"3a4b",x"33f0",x"3a26",x"3d45",x"36da",x"3bff",x"26b5",x"0000",x"3a38",x"33fa",x"3a25",x"3d5c",x"3710",x"3bd6",x"2604",x"3256",x"3a49",x"33c0"),
(x"35fd",x"3d4e",x"36da",x"3bf0",x"2ff4",x"8000",x"3a18",x"39dc",x"35fd",x"3d4c",x"36da",x"3a08",x"b941",x"8000",x"3a18",x"39db",x"35fd",x"3d4e",x"3710",x"3b91",x"3530",x"8000",x"3a23",x"39dc"),
(x"3593",x"3d72",x"36da",x"bbda",x"b21b",x"0000",x"3b06",x"3a0f",x"3587",x"3d77",x"36da",x"bbf7",x"adba",x"8000",x"3b06",x"3a0b",x"3593",x"3d72",x"3710",x"bc00",x"15bc",x"0000",x"3b11",x"3a0f"),
(x"38d5",x"3d5f",x"36da",x"2dde",x"bbf7",x"0000",x"3a44",x"39d8",x"38bf",x"3d5d",x"36da",x"35f3",x"bb6c",x"0000",x"3a44",x"39cf",x"38d5",x"3d5f",x"3710",x"1987",x"bc00",x"0000",x"3a4f",x"39d8"),
(x"38d8",x"3d84",x"36da",x"3be4",x"312f",x"8000",x"3a93",x"3ad6",x"38d9",x"3d82",x"36da",x"3b88",x"b564",x"0000",x"3a93",x"3ad5",x"38d8",x"3d84",x"3710",x"3b96",x"350f",x"0000",x"3a9e",x"3ad6"),
(x"35fd",x"3d4c",x"36da",x"3a08",x"b941",x"8000",x"3a18",x"39db",x"35f5",x"3d4b",x"36da",x"32d5",x"bbd0",x"0000",x"3a18",x"39d9",x"35fd",x"3d4c",x"3710",x"3b87",x"b567",x"868d",x"3a23",x"39db"),
(x"3592",x"3d70",x"36da",x"bba4",x"34bb",x"0000",x"3b06",x"3a11",x"3593",x"3d72",x"36da",x"bbda",x"b21b",x"0000",x"3b06",x"3a0f",x"3592",x"3d70",x"3710",x"ba08",x"3941",x"0000",x"3b11",x"3a11"),
(x"38bf",x"3d5d",x"36da",x"35f3",x"bb6c",x"0000",x"3a44",x"39cf",x"38b2",x"3d5a",x"36da",x"3af2",x"b7f0",x"0000",x"3a44",x"39ca",x"38bf",x"3d5d",x"3710",x"3489",x"bbab",x"0000",x"3a4f",x"39cf"),
(x"38c7",x"3d87",x"36da",x"3654",x"3b58",x"8000",x"3a93",x"3add",x"38d8",x"3d84",x"36da",x"3be4",x"312f",x"8000",x"3a93",x"3ad6",x"38c7",x"3d87",x"3710",x"364a",x"3b5a",x"0000",x"3a9e",x"3add"),
(x"35f5",x"3d4b",x"36da",x"32d5",x"bbd0",x"0000",x"3a18",x"39d9",x"35e4",x"3d4b",x"36da",x"b3c3",x"bbc2",x"0000",x"3a18",x"39d6",x"35f5",x"3d4b",x"3710",x"364b",x"bb5a",x"0000",x"3a23",x"39d9"),
(x"357d",x"3d70",x"36da",x"a8c9",x"3bfe",x"0000",x"3a5f",x"3b39",x"3592",x"3d70",x"36da",x"bba4",x"34bb",x"0000",x"3a5f",x"3b35",x"357d",x"3d70",x"3710",x"26bb",x"3bff",x"0000",x"3a6a",x"3b39"),
(x"38b2",x"3d5a",x"36da",x"3af2",x"b7f0",x"0000",x"3a33",x"3a19",x"38b0",x"3d57",x"36da",x"3ba6",x"34ab",x"0000",x"3a33",x"3a17",x"38b2",x"3d5a",x"3710",x"3a0a",x"b93f",x"0000",x"3a3e",x"3a19"),
(x"38b7",x"3d8b",x"36da",x"3528",x"3b92",x"8000",x"3a93",x"3ae4",x"38c7",x"3d87",x"36da",x"3654",x"3b58",x"8000",x"3a93",x"3add",x"38b7",x"3d8b",x"3710",x"32f6",x"3bce",x"0000",x"3a9e",x"3ae4"),
(x"35e4",x"3d4b",x"36da",x"b3c3",x"bbc2",x"0000",x"3a18",x"39d6",x"35d3",x"3d4c",x"36da",x"1c81",x"bc00",x"0000",x"3a18",x"39d2",x"35e4",x"3d4b",x"3710",x"b0fa",x"bbe7",x"8000",x"3a23",x"39d6"),
(x"3555",x"3d71",x"36da",x"345a",x"3bb2",x"0000",x"3a5f",x"3b40",x"357d",x"3d70",x"36da",x"a8c9",x"3bfe",x"0000",x"3a5f",x"3b39",x"3555",x"3d71",x"3710",x"35eb",x"3b6e",x"0000",x"3a6a",x"3b40"),
(x"38b0",x"3d57",x"36da",x"3ba6",x"34ab",x"0000",x"3a33",x"3a17",x"38b2",x"3d55",x"36da",x"399c",x"39b3",x"8000",x"3a33",x"3a15",x"38b0",x"3d57",x"3710",x"3bfc",x"ab2b",x"0000",x"3a3e",x"3a17"),
(x"3894",x"3d8c",x"36da",x"aa0a",x"3bfd",x"8000",x"3a93",x"3af1",x"38b7",x"3d8b",x"36da",x"3528",x"3b92",x"8000",x"3a93",x"3ae4",x"3894",x"3d8c",x"3710",x"b036",x"3bee",x"0000",x"3a9e",x"3af1"),
(x"35d3",x"3d4c",x"36da",x"1c81",x"bc00",x"0000",x"3a18",x"39d2",x"35bd",x"3d4b",x"36da",x"afc9",x"bbf0",x"8000",x"3a18",x"39ce",x"35d3",x"3d4c",x"3710",x"b1d2",x"bbdd",x"0000",x"3a23",x"39d2"),
(x"353f",x"3d74",x"36da",x"3746",x"3b1f",x"0000",x"3a5f",x"3b45",x"3555",x"3d71",x"36da",x"345a",x"3bb2",x"0000",x"3a5f",x"3b40",x"353f",x"3d74",x"3710",x"379f",x"3b08",x"0000",x"3a6a",x"3b45"),
(x"38b2",x"3d55",x"36da",x"399c",x"39b3",x"8000",x"3a33",x"3a15",x"38bd",x"3d52",x"36da",x"3456",x"3bb3",x"0000",x"3a33",x"3a11",x"38b2",x"3d55",x"3710",x"3a58",x"38de",x"0000",x"3a3e",x"3a15"),
(x"3877",x"3d89",x"36da",x"b74e",x"3b1d",x"0000",x"3a93",x"3afc",x"3894",x"3d8c",x"36da",x"aa0a",x"3bfd",x"8000",x"3a93",x"3af1",x"3877",x"3d89",x"3710",x"b8aa",x"3a7f",x"8000",x"3a9e",x"3afc"),
(x"35bd",x"3d4b",x"36da",x"afc9",x"bbf0",x"8000",x"3a18",x"39ce",x"359e",x"3d4e",x"36da",x"b925",x"ba1f",x"8000",x"3a18",x"39c8",x"35bd",x"3d4b",x"3710",x"2c74",x"bbfb",x"068d",x"3a23",x"39ce"),
(x"351b",x"3d79",x"36da",x"3664",x"3b55",x"0000",x"3a5f",x"3b4d",x"353f",x"3d74",x"36da",x"3746",x"3b1f",x"0000",x"3a5f",x"3b45",x"351b",x"3d79",x"3710",x"350e",x"3b96",x"0000",x"3a6a",x"3b4d"),
(x"38bd",x"3d52",x"36da",x"3456",x"3bb3",x"0000",x"3a33",x"3a11",x"38c9",x"3d51",x"36da",x"34cb",x"3ba1",x"8000",x"3a33",x"3a0c",x"38bd",x"3d52",x"3710",x"35fc",x"3b6b",x"0000",x"3a3e",x"3a11"),
(x"386d",x"3d84",x"36da",x"bac4",x"3844",x"8000",x"3a93",x"3b01",x"3877",x"3d89",x"36da",x"b74e",x"3b1d",x"0000",x"3a93",x"3afc",x"386d",x"3d84",x"3710",x"bba8",x"34a3",x"0000",x"3a9e",x"3b01"),
(x"359e",x"3d4e",x"36da",x"b925",x"ba1f",x"8000",x"3a18",x"39c8",x"358a",x"3d54",x"36da",x"bbad",x"b481",x"8000",x"3a18",x"39c2",x"359e",x"3d4e",x"3710",x"b80b",x"bae7",x"0000",x"3a23",x"39c8"),
(x"3501",x"3d7b",x"36da",x"2d0c",x"3bf9",x"8000",x"3a5f",x"3b52",x"351b",x"3d79",x"36da",x"3664",x"3b55",x"0000",x"3a5f",x"3b4d",x"3501",x"3d7b",x"3710",x"ada6",x"3bf8",x"0000",x"3a6a",x"3b52"),
(x"38c9",x"3d51",x"36da",x"34cb",x"3ba1",x"8000",x"3a33",x"3a0c",x"38d4",x"3d4f",x"36da",x"38a8",x"3a80",x"8000",x"3a33",x"3a08",x"38c9",x"3d51",x"3710",x"3385",x"3bc6",x"0000",x"3a3e",x"3a0c"),
(x"386c",x"3d7f",x"36da",x"bbdd",x"b1e1",x"8000",x"3a93",x"3b05",x"386d",x"3d84",x"36da",x"bac4",x"3844",x"8000",x"3a93",x"3b01",x"386c",x"3d7f",x"3710",x"bb38",x"b6e2",x"868d",x"3a9e",x"3b05"),
(x"358a",x"3d54",x"36da",x"bbad",x"b481",x"8000",x"3a18",x"39c2",x"3587",x"3d59",x"36da",x"bb8b",x"3553",x"0000",x"3a18",x"39be",x"358a",x"3d54",x"3710",x"bb1e",x"b74c",x"0000",x"3a23",x"39c2"),
(x"34e9",x"3d79",x"36da",x"b50d",x"3b97",x"8000",x"3a5f",x"3b57",x"3501",x"3d7b",x"36da",x"2d0c",x"3bf9",x"8000",x"3a5f",x"3b52",x"34e9",x"3d79",x"3710",x"b698",x"3b49",x"0000",x"3a6a",x"3b57"),
(x"38d4",x"3d4f",x"36da",x"38a8",x"3a80",x"8000",x"3a33",x"3a08",x"38d9",x"3d4d",x"36da",x"3bfc",x"2b00",x"8000",x"3a33",x"3a06",x"38d4",x"3d4f",x"3710",x"37f2",x"3af1",x"8000",x"3a3e",x"3a08"),
(x"3872",x"3d7b",x"36da",x"b9d1",x"b97d",x"8000",x"3a93",x"3b08",x"386c",x"3d7f",x"36da",x"bbdd",x"b1e1",x"8000",x"3a93",x"3b05",x"3872",x"3d7b",x"3710",x"b902",x"ba3c",x"0000",x"3a9e",x"3b08"),
(x"3587",x"3d59",x"36da",x"bb8b",x"3553",x"0000",x"3a18",x"39be",x"3593",x"3d5d",x"36da",x"bc00",x"95bc",x"0000",x"3a18",x"39ba",x"3587",x"3d59",x"3710",x"bbf7",x"2dba",x"0000",x"3a23",x"39be"),
(x"34cb",x"3d75",x"36da",x"b64c",x"3b5a",x"0000",x"3a5f",x"3b5d",x"34e9",x"3d79",x"36da",x"b50d",x"3b97",x"8000",x"3a5f",x"3b57",x"34cb",x"3d75",x"3710",x"b501",x"3b99",x"0000",x"3a6a",x"3b5d"),
(x"38d9",x"3d4d",x"36da",x"3bfc",x"2b00",x"8000",x"3a33",x"3a06",x"38d8",x"3d4c",x"36da",x"3b96",x"b50f",x"0000",x"3a33",x"3a05",x"38d9",x"3d4d",x"3710",x"3b88",x"3564",x"0000",x"3a3e",x"3a06"),
(x"3885",x"3d77",x"36da",x"b7eb",x"baf3",x"0000",x"3a93",x"3b10",x"3872",x"3d7b",x"36da",x"b9d1",x"b97d",x"8000",x"3a93",x"3b08",x"3885",x"3d77",x"3710",x"b83d",x"bac8",x"0000",x"3a9e",x"3b10"),
(x"3593",x"3d5d",x"36da",x"bc00",x"95bc",x"0000",x"3a18",x"39ba",x"3592",x"3d60",x"36da",x"ba08",x"b941",x"8000",x"3a18",x"39b8",x"3593",x"3d5d",x"3710",x"bbda",x"321b",x"8000",x"3a23",x"39ba"),
(x"34bb",x"3d73",x"36da",x"b31c",x"3bcc",x"0000",x"3a5f",x"3b60",x"34cb",x"3d75",x"36da",x"b64c",x"3b5a",x"0000",x"3a5f",x"3b5d",x"34bb",x"3d73",x"3710",x"b13f",x"3be4",x"0000",x"3a6a",x"3b60"),
(x"38d8",x"3d4c",x"36da",x"3b96",x"b50f",x"0000",x"3a33",x"3a05",x"38c7",x"3d48",x"36da",x"364a",x"bb5b",x"8000",x"3a33",x"39fd",x"38d8",x"3d4c",x"3710",x"3be4",x"b12f",x"8a8d",x"3a3e",x"3a05"),
(x"388c",x"3d75",x"36da",x"bb54",x"b669",x"8000",x"3a93",x"3b13",x"3885",x"3d77",x"36da",x"b7eb",x"baf3",x"0000",x"3a93",x"3b10",x"388c",x"3d75",x"3710",x"bbfd",x"a9ab",x"0000",x"3a9e",x"3b13"),
(x"3592",x"3d60",x"36da",x"ba08",x"b941",x"8000",x"3a5f",x"3bb1",x"357d",x"3d60",x"36da",x"26c8",x"bbff",x"0000",x"3a5f",x"3bad",x"3592",x"3d60",x"3710",x"bba4",x"b4bb",x"0000",x"3a6a",x"3bb1"),
(x"349b",x"3d73",x"36da",x"b221",x"3bda",x"0000",x"3a5f",x"3b66",x"34bb",x"3d73",x"36da",x"b31c",x"3bcc",x"0000",x"3a5f",x"3b60",x"349b",x"3d73",x"3710",x"b4a8",x"3ba7",x"0000",x"3a6a",x"3b66"),
(x"38c7",x"3d48",x"36da",x"364a",x"bb5b",x"8000",x"3a33",x"39fd",x"38b7",x"3d45",x"36da",x"32f6",x"bbce",x"0000",x"3a33",x"39f7",x"38c7",x"3d48",x"3710",x"3653",x"bb59",x"0000",x"3a3e",x"39fd"),
(x"388c",x"3d73",x"36da",x"bb52",x"3671",x"0000",x"3a3d",x"3bb0",x"388c",x"3d75",x"36da",x"bb54",x"b669",x"8000",x"3a3d",x"3bb1",x"388c",x"3d73",x"3710",x"b967",x"39e6",x"0000",x"3a32",x"3bb0"),
(x"357d",x"3d60",x"36da",x"26c8",x"bbff",x"0000",x"3a5f",x"3bad",x"3555",x"3d5f",x"36da",x"35eb",x"bb6e",x"0000",x"3a5f",x"3ba5",x"357d",x"3d60",x"3710",x"a8c9",x"bbfe",x"0000",x"3a6a",x"3bad"),
(x"3485",x"3d71",x"36da",x"b819",x"3ade",x"8000",x"3a5f",x"3b6b",x"349b",x"3d73",x"36da",x"b221",x"3bda",x"0000",x"3a5f",x"3b66",x"3485",x"3d71",x"3710",x"b92c",x"3a1a",x"0000",x"3a6a",x"3b6b"),
(x"38b7",x"3d45",x"36da",x"32f6",x"bbce",x"0000",x"3a33",x"39f7",x"3894",x"3d44",x"36da",x"b036",x"bbee",x"0000",x"3a33",x"39ea",x"38b7",x"3d45",x"3710",x"3528",x"bb92",x"0000",x"3a3e",x"39f7"),
(x"3885",x"3d72",x"36da",x"b304",x"3bce",x"0000",x"3a3d",x"3bad",x"388c",x"3d73",x"36da",x"bb52",x"3671",x"0000",x"3a3d",x"3bb0",x"3885",x"3d72",x"3710",x"b25f",x"3bd7",x"8000",x"3a32",x"3bad"),
(x"3555",x"3d5f",x"36da",x"35eb",x"bb6e",x"0000",x"3a5f",x"3ba5",x"353f",x"3d5c",x"36da",x"379f",x"bb08",x"0000",x"3a5f",x"3ba1",x"3555",x"3d5f",x"3710",x"345a",x"bbb2",x"0000",x"3a6a",x"3ba5"),
(x"3475",x"3d6c",x"36da",x"baeb",x"3803",x"868d",x"3a5f",x"3b70",x"3485",x"3d71",x"36da",x"b819",x"3ade",x"8000",x"3a5f",x"3b6b",x"3475",x"3d6c",x"3710",x"bbab",x"348e",x"8000",x"3a6a",x"3b70"),
(x"3894",x"3d44",x"36da",x"b036",x"bbee",x"0000",x"3a33",x"39ea",x"3877",x"3d47",x"36da",x"b8aa",x"ba7f",x"8000",x"3a33",x"39de",x"3894",x"3d44",x"3710",x"aa0a",x"bbfd",x"8000",x"3a3e",x"39ea"),
(x"3753",x"3d89",x"36da",x"38fe",x"3a3f",x"8000",x"3a3d",x"3b48",x"3760",x"3d86",x"36da",x"3bfa",x"2cac",x"8000",x"3a3d",x"3b4c",x"3753",x"3d89",x"3710",x"37e4",x"3af5",x"8000",x"3a32",x"3b48"),
(x"3a2f",x"3d73",x"36da",x"3bfe",x"a8f0",x"0000",x"3bfb",x"3999",x"3a2d",x"3d5e",x"36da",x"3bfe",x"a8f0",x"0000",x"3bea",x"3999",x"3a2f",x"3d73",x"3710",x"3b78",x"a99e",x"35b0",x"3bfb",x"398f"),
(x"353f",x"3d5c",x"36da",x"379f",x"bb08",x"0000",x"3a5f",x"3ba1",x"351b",x"3d57",x"36da",x"350e",x"bb96",x"0000",x"3a5f",x"3b99",x"353f",x"3d5c",x"3710",x"3746",x"bb1f",x"0000",x"3a6a",x"3ba1"),
(x"39f5",x"3d8a",x"36da",x"a49b",x"3bff",x"8000",x"3bd5",x"3a14",x"3a27",x"3d8b",x"36da",x"a3ae",x"3bff",x"0000",x"3bd5",x"3a28",x"39f5",x"3d8a",x"3710",x"a4e3",x"3bff",x"1818",x"3bcb",x"3a14"),
(x"3877",x"3d47",x"36da",x"b8aa",x"ba7f",x"8000",x"3a33",x"39de",x"386d",x"3d4b",x"36da",x"bba8",x"b4a3",x"868d",x"3a33",x"39d9",x"3877",x"3d47",x"3710",x"b74e",x"bb1d",x"8000",x"3a3e",x"39de"),
(x"382a",x"3d72",x"36da",x"2f40",x"3bf2",x"8000",x"3a3d",x"3b89",x"3885",x"3d72",x"36da",x"b304",x"3bce",x"0000",x"3a3d",x"3bad",x"382a",x"3d72",x"3710",x"30bd",x"3be9",x"8000",x"3a32",x"3b89"),
(x"351b",x"3d57",x"36da",x"350e",x"bb96",x"0000",x"3a5f",x"3b99",x"3501",x"3d55",x"36da",x"ada8",x"bbf8",x"8000",x"3a5f",x"3b94",x"351b",x"3d57",x"3710",x"3664",x"bb55",x"0000",x"3a6a",x"3b99"),
(x"386d",x"3d4b",x"36da",x"bba8",x"b4a3",x"868d",x"3a33",x"39d9",x"386c",x"3d51",x"36da",x"bb38",x"36e2",x"068d",x"3a33",x"39d5",x"386d",x"3d4b",x"3710",x"bac4",x"b844",x"0000",x"3a3e",x"39d9"),
(x"3813",x"3d74",x"36da",x"27fc",x"3bfe",x"0000",x"3a3d",x"3b80",x"382a",x"3d72",x"36da",x"2f40",x"3bf2",x"8000",x"3a3d",x"3b89",x"3813",x"3d74",x"3710",x"a8bf",x"3bfe",x"8000",x"3a32",x"3b80"),
(x"3a2d",x"3d5e",x"36da",x"367a",x"bb50",x"0000",x"3bc0",x"39b2",x"3a25",x"3d5c",x"36da",x"367a",x"bb50",x"0000",x"3bc3",x"39b4",x"3a2d",x"3d5e",x"3710",x"3644",x"bb4c",x"2f83",x"3bba",x"39ba"),
(x"359e",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2a4d",x"35f7",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39dd",x"2b8b",x"3593",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2a24"),
(x"359e",x"403a",x"3710",x"0000",x"0000",x"3c00",x"39b7",x"2a4d",x"3593",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2a27",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b"),
(x"3592",x"3d70",x"3710",x"0000",x"0000",x"3c00",x"3a59",x"2a20",x"3593",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2a22",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"359e",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2a4d",x"358a",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2a0e",x"3593",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2a27"),
(x"359e",x"3d4e",x"3710",x"0000",x"0000",x"3c00",x"3a3b",x"2a4d",x"3593",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2a27",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b"),
(x"38b2",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"30f2",x"38b7",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"30f9",x"38bd",x"3d7d",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"3107"),
(x"38c9",x"3d51",x"3710",x"0000",x"0000",x"3c00",x"3a3e",x"311a",x"38b7",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30f9",x"38bd",x"3d52",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"3107"),
(x"2da5",x"4061",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"3ab5",x"2a34",x"4061",x"36fa",x"0000",x"8000",x"bc00",x"3557",x"3ab5",x"2da5",x"3d34",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"38f4"),
(x"2a34",x"4061",x"36fa",x"baf4",x"0000",x"37e6",x"35b0",x"3a80",x"2af5",x"405d",x"3725",x"baf4",x"0000",x"37e6",x"35bc",x"3a7b",x"2a34",x"3d34",x"36fa",x"baf4",x"0000",x"37e6",x"35b0",x"38f4"),
(x"2d44",x"3d3c",x"3725",x"0000",x"0000",x"3c00",x"3571",x"38f4",x"2af5",x"3d3c",x"3725",x"0000",x"0000",x"3c00",x"3558",x"38f4",x"2d44",x"405d",x"3725",x"0000",x"0000",x"3c00",x"3571",x"3aad"),
(x"2d44",x"405d",x"3725",x"0000",x"3a66",x"38cc",x"3b15",x"3b97",x"2af5",x"405d",x"3725",x"0000",x"3a66",x"38cc",x"3b06",x"3b97",x"2da5",x"4061",x"36fa",x"0000",x"3a66",x"38cc",x"3b19",x"3ba0"),
(x"2a34",x"3d34",x"36fa",x"0000",x"ba66",x"38cc",x"3b02",x"3ba8",x"2af5",x"3d3c",x"3725",x"0000",x"ba66",x"38cc",x"3b06",x"3bb1",x"2da5",x"3d34",x"36fa",x"0000",x"ba66",x"38cc",x"3b19",x"3ba8"),
(x"2da5",x"4061",x"36fa",x"3af5",x"0000",x"37e6",x"35a3",x"3a7f",x"2da5",x"3d34",x"36fa",x"3af4",x"0000",x"37e6",x"35a3",x"38f4",x"2d44",x"405d",x"3725",x"3af5",x"0000",x"37e6",x"3597",x"3a7c"),
(x"2a34",x"4061",x"36fa",x"0000",x"8000",x"bc00",x"3557",x"3ab5",x"2a34",x"3d34",x"36fa",x"0000",x"8000",x"bc00",x"3557",x"38f4",x"2da5",x"3d34",x"36fa",x"0000",x"8000",x"bc00",x"3533",x"38f4"),
(x"2af5",x"405d",x"3725",x"baf4",x"0000",x"37e6",x"35bc",x"3a7b",x"2af5",x"3d3c",x"3725",x"baf4",x"0000",x"37e6",x"35bc",x"38f7",x"2a34",x"3d34",x"36fa",x"baf4",x"0000",x"37e6",x"35b0",x"38f4"),
(x"2af5",x"3d3c",x"3725",x"0000",x"0000",x"3c00",x"3558",x"38f4",x"2af5",x"405d",x"3725",x"0000",x"0000",x"3c00",x"3558",x"3aad",x"2d44",x"405d",x"3725",x"0000",x"0000",x"3c00",x"3571",x"3aad"),
(x"2af5",x"405d",x"3725",x"0000",x"3a66",x"38cc",x"3b06",x"3b97",x"2a34",x"4061",x"36fa",x"0000",x"3a66",x"38cc",x"3b02",x"3ba0",x"2da5",x"4061",x"36fa",x"0000",x"3a66",x"38cc",x"3b19",x"3ba0"),
(x"2af5",x"3d3c",x"3725",x"0000",x"ba66",x"38cc",x"3b06",x"3bb1",x"2d44",x"3d3c",x"3725",x"0000",x"ba66",x"38cc",x"3b15",x"3bb1",x"2da5",x"3d34",x"36fa",x"0000",x"ba66",x"38cc",x"3b19",x"3ba8"),
(x"2da5",x"3d34",x"36fa",x"3af4",x"0000",x"37e6",x"35a3",x"38f4",x"2d44",x"3d3c",x"3725",x"3af4",x"0000",x"37e6",x"3597",x"38f8",x"2d44",x"405d",x"3725",x"3af5",x"0000",x"37e6",x"3597",x"3a7c"),
(x"2f99",x"3ef2",x"36b4",x"0000",x"0000",x"3c00",x"3a76",x"3515",x"3004",x"3eee",x"36b4",x"0000",x"0000",x"3c00",x"3a78",x"351c",x"3009",x"3eea",x"36b4",x"0000",x"0000",x"3c00",x"3a7a",x"351c"),
(x"2fe5",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7c",x"3519",x"2f19",x"3eef",x"36b4",x"0000",x"0000",x"3c00",x"3a77",x"350d",x"2f99",x"3ef2",x"36b4",x"0000",x"0000",x"3c00",x"3a76",x"3515"),
(x"2f10",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7d",x"350c",x"2ee6",x"3eea",x"36b4",x"0000",x"0000",x"3c00",x"3a7a",x"350a",x"2f19",x"3eef",x"36b4",x"0000",x"0000",x"3c00",x"3a77",x"350d"),
(x"2fda",x"3ee2",x"36b4",x"0000",x"0000",x"3c00",x"3a7e",x"3519",x"2f02",x"3ec3",x"36b4",x"0000",x"0000",x"3c00",x"3a8b",x"350b",x"2f10",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7d",x"350c"),
(x"2fda",x"3ee2",x"36b4",x"0000",x"0000",x"3c00",x"3a7e",x"3519",x"3025",x"3ec3",x"36b4",x"0000",x"0000",x"3c00",x"3a8b",x"351f",x"2f02",x"3ec3",x"36b4",x"0000",x"0000",x"3c00",x"3a8b",x"350b"),
(x"2fe5",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7c",x"3519",x"2f10",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7d",x"350c",x"2f19",x"3eef",x"36b4",x"0000",x"0000",x"3c00",x"3a77",x"350d"),
(x"2f99",x"3ef2",x"36b4",x"0000",x"0000",x"3c00",x"3a76",x"3515",x"3009",x"3eea",x"36b4",x"0000",x"0000",x"3c00",x"3a7a",x"351c",x"2fe5",x"3ee4",x"36b4",x"0000",x"0000",x"3c00",x"3a7c",x"3519"),
(x"358a",x"403d",x"3710",x"0000",x"0000",x"3c00",x"39bb",x"2a0d",x"3587",x"4040",x"3710",x"0000",x"0000",x"3c00",x"39bf",x"2a03",x"3593",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2a27"),
(x"38b7",x"4036",x"3710",x"0000",x"0000",x"3c00",x"39af",x"30f9",x"38b2",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"30f2",x"38bd",x"403d",x"3710",x"0000",x"0000",x"3c00",x"39bc",x"3107"),
(x"38b7",x"4059",x"3710",x"0000",x"0000",x"3c00",x"39eb",x"30f9",x"38c9",x"4053",x"3710",x"0000",x"0000",x"3c00",x"39e0",x"311a",x"38bd",x"4052",x"3710",x"0000",x"0000",x"3c00",x"39de",x"3107"),
(x"358a",x"3d7c",x"3710",x"0000",x"0000",x"3c00",x"3a63",x"2a04",x"359e",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a68",x"2a4d",x"3593",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2a22"),
(x"358a",x"4051",x"3710",x"0000",x"0000",x"3c00",x"39de",x"2a05",x"359e",x"4054",x"3710",x"0000",x"0000",x"3c00",x"39e3",x"2a4d",x"3593",x"404d",x"3710",x"0000",x"0000",x"3c00",x"39d6",x"2a24"),
(x"3593",x"4042",x"3710",x"0000",x"0000",x"3c00",x"39c2",x"2a27",x"3592",x"4043",x"3710",x"0000",x"0000",x"3c00",x"39c6",x"2a20",x"35f7",x"403e",x"3710",x"0000",x"0000",x"3c00",x"39bd",x"2b8b"),
(x"3593",x"3d72",x"3710",x"0000",x"0000",x"3c00",x"3a5a",x"2a22",x"359e",x"3d82",x"3710",x"0000",x"0000",x"3c00",x"3a68",x"2a4d",x"35f7",x"3d7a",x"3710",x"0000",x"0000",x"3c00",x"3a61",x"2b8b"),
(x"358a",x"3d54",x"3710",x"0000",x"0000",x"3c00",x"3a40",x"2a0e",x"3587",x"3d59",x"3710",x"0000",x"0000",x"3c00",x"3a43",x"2a04",x"3593",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2a27"),
(x"3593",x"3d5d",x"3710",x"0000",x"0000",x"3c00",x"3a47",x"2a27",x"3592",x"3d60",x"3710",x"0000",x"0000",x"3c00",x"3a4a",x"2a20",x"35f7",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"2b8b"),
(x"38b7",x"3d8b",x"3710",x"0000",x"0000",x"3c00",x"3a6f",x"30f9",x"38c9",x"3d7e",x"3710",x"0000",x"0000",x"3c00",x"3a65",x"311a",x"38bd",x"3d7d",x"3710",x"0000",x"0000",x"3c00",x"3a62",x"3107"),
(x"38b7",x"3d45",x"3710",x"0000",x"0000",x"3c00",x"3a33",x"30f9",x"38b2",x"3d55",x"3710",x"0000",x"0000",x"3c00",x"3a42",x"30f2",x"38bd",x"3d52",x"3710",x"0000",x"0000",x"3c00",x"3a41",x"3107"),
(x"b936",x"4062",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"3a68",x"b936",x"3d32",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"38f3",x"b936",x"4062",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"3a68"),
(x"2af5",x"3ee9",x"36b2",x"3c00",x"8000",x"0000",x"371d",x"30fe",x"2af5",x"3ee9",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30fe",x"2af5",x"4062",x"368e",x"3c00",x"8000",x"0000",x"3732",x"345d"),
(x"aaef",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3af7",x"3815",x"aaef",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3af7",x"3810",x"b858",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3a04",x"3815"),
(x"b936",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3a0a",x"b936",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3a0a",x"2af5",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3b6a"),
(x"2af5",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"3ada",x"b936",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"397a",x"2af5",x"4062",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"3ada"),
(x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"b86b",x"4016",x"36fb",x"0000",x"8000",x"3c00",x"39eb",x"3bb1",x"b86c",x"3dde",x"36fb",x"0000",x"8000",x"3c00",x"39eb",x"3ad5"),
(x"9da8",x"3eee",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b3b",x"9e2f",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b39",x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0"),
(x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95",x"b936",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3a95",x"aaef",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3ac4"),
(x"b858",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3bbc",x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"aaef",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3bbc"),
(x"aaef",x"3dae",x"36d0",x"0000",x"8000",x"3c00",x"3742",x"3adb",x"b858",x"3dae",x"36d0",x"0000",x"8000",x"3c00",x"35d9",x"3adb",x"aaef",x"4024",x"36d0",x"0000",x"8000",x"3c00",x"3742",x"3bfa"),
(x"aaef",x"3dae",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"3dc7",x"36e5",x"bc00",x"0000",x"0000",x"3ae4",x"3545",x"aaef",x"3dbd",x"36fb",x"bc00",x"0000",x"0000",x"3ae5",x"3546"),
(x"b858",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3a05",x"3821",x"b858",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3a05",x"3826",x"aaef",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3af8",x"3821"),
(x"a9a6",x"4015",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8",x"aaef",x"4016",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"aa60",x"401e",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1"),
(x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95",x"aaef",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3ac4",x"aa24",x"3dc9",x"36fb",x"0000",x"8000",x"3c00",x"3ab0",x"3ace"),
(x"aa60",x"401e",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1",x"aaef",x"401e",x"36e4",x"ba1e",x"b322",x"38d5",x"351b",x"38d1",x"aaef",x"4022",x"36fb",x"b9d6",x"b5ae",x"38ac",x"351f",x"38d6"),
(x"aaef",x"3dae",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"4024",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"3dd5",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545"),
(x"aaef",x"4024",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"4024",x"36fb",x"bc00",x"0000",x"0000",x"3a7f",x"3557",x"aaef",x"4022",x"36fb",x"bc00",x"0000",x"0000",x"3a83",x"3557"),
(x"a9ae",x"3dd7",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3ad3",x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95",x"aa24",x"3dc9",x"36fb",x"0000",x"8000",x"3c00",x"3ab0",x"3ace"),
(x"a9ae",x"3dd7",x"36fb",x"b993",x"1c9b",x"39bd",x"3526",x"3740",x"aaef",x"3dd5",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"a9a6",x"4015",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8"),
(x"aaef",x"3dc7",x"36e5",x"b96c",x"347c",x"396f",x"351c",x"3730",x"aaef",x"3dd5",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"aa24",x"3dc9",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"aaef",x"3dbd",x"36fb",x"b969",x"359e",x"392e",x"351f",x"3725",x"aaef",x"3dc7",x"36e5",x"b96c",x"347c",x"396f",x"351c",x"3730",x"aa24",x"3dc9",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"b857",x"401d",x"36e5",x"3bfe",x"2111",x"a780",x"3b41",x"34eb",x"b857",x"4023",x"36fb",x"3bfe",x"276c",x"a4f7",x"3b42",x"34ec",x"b858",x"4024",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9"),
(x"b858",x"3dae",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b858",x"3dae",x"36fb",x"3bff",x"a5e9",x"0000",x"3ad1",x"34ff",x"b857",x"3dbb",x"36fb",x"3bff",x"a3a0",x"a0dd",x"3ade",x"3501"),
(x"b863",x"3dc6",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0",x"b857",x"3dc6",x"36dd",x"3a1a",x"3321",x"38da",x"357e",x"38d0",x"b857",x"3dbb",x"36fb",x"39d1",x"35ef",x"389f",x"3584",x"38d6"),
(x"b857",x"4016",x"36d8",x"3bf1",x"15bc",x"afa2",x"3b3f",x"34eb",x"b858",x"4024",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b857",x"3ddc",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed"),
(x"b86c",x"3dde",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4",x"b857",x"3ddc",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b863",x"3dc6",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0"),
(x"b86b",x"4016",x"36fb",x"3935",x"9d6d",x"3a12",x"3587",x"373c",x"b857",x"4016",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b86c",x"3dde",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4"),
(x"b857",x"401d",x"36e5",x"397e",x"b36f",x"3983",x"357d",x"372e",x"b857",x"4016",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b862",x"401d",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"b857",x"4023",x"36fb",x"3958",x"b562",x"394e",x"3580",x"3722",x"b857",x"401d",x"36e5",x"397e",x"b36f",x"3983",x"357d",x"372e",x"b862",x"401d",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"2163",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b2b",x"20f3",x"3ee4",x"36fb",x"0000",x"8000",x"3c00",x"3ac6",x"3b37",x"2243",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b39"),
(x"b936",x"3d32",x"368e",x"0000",x"0000",x"bc00",x"3a79",x"30b7",x"2af5",x"3d32",x"368e",x"0000",x"0000",x"bc00",x"3b35",x"30b7",x"b936",x"4062",x"368e",x"0000",x"0000",x"bc00",x"3a79",x"290e"),
(x"9ac5",x"3ee4",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"9e2f",x"3eea",x"36fb",x"3b8f",x"3538",x"068d",x"3a18",x"3614",x"9ac5",x"3ee4",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603"),
(x"2163",x"3ec3",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a47",x"a0d7",x"3ec3",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a51",x"2163",x"3ec3",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a47"),
(x"20b0",x"3eef",x"36fb",x"b727",x"bb27",x"868d",x"3a23",x"3614",x"2243",x"3eea",x"36fb",x"bbcf",x"b2e8",x"0000",x"3a26",x"3614",x"20b0",x"3eef",x"36b4",x"b93c",x"ba0c",x"8000",x"3a23",x"3603"),
(x"9e2f",x"3eea",x"36fb",x"3b8f",x"3538",x"068d",x"3a18",x"3614",x"9da8",x"3eee",x"36fb",x"3aa7",x"b870",x"0000",x"3a1b",x"3614",x"9e2f",x"3eea",x"36b4",x"3bef",x"3011",x"8000",x"3a18",x"3603"),
(x"a0d7",x"3ec3",x"36fb",x"3bcb",x"b335",x"0000",x"3a04",x"3614",x"995f",x"3ee2",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"a0d7",x"3ec3",x"36b4",x"3bcb",x"b335",x"0000",x"3a04",x"3603"),
(x"2243",x"3eea",x"36fb",x"bbcf",x"b2e8",x"0000",x"3a26",x"3614",x"20f3",x"3ee4",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"2243",x"3eea",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603"),
(x"9da8",x"3eee",x"36fb",x"3aa7",x"b870",x"0000",x"3a1b",x"3614",x"1557",x"3ef2",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"9da8",x"3eee",x"36b4",x"38fa",x"ba42",x"8000",x"3a1b",x"3603"),
(x"995f",x"3ee2",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"9ac5",x"3ee4",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"995f",x"3ee2",x"36b4",x"3be8",x"b0e3",x"8000",x"3a14",x"3603"),
(x"20f3",x"3ee4",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"2163",x"3ec3",x"36fb",x"bbff",x"a6cf",x"0000",x"3a3b",x"3614",x"20f3",x"3ee4",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603"),
(x"1557",x"3ef2",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"20b0",x"3eef",x"36fb",x"b727",x"bb27",x"868d",x"3a23",x"3614",x"1557",x"3ef2",x"36b4",x"a8d6",x"bbfe",x"0000",x"3a1f",x"3603"),
(x"9ac5",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a18",x"20f3",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a12",x"995f",x"3ee2",x"36b4",x"0000",x"8000",x"3c00",x"3b69",x"3a18"),
(x"2af5",x"3ed3",x"36b2",x"3c00",x"8000",x"0000",x"371d",x"30d2",x"2af5",x"3ee9",x"36b2",x"3c00",x"8000",x"0000",x"371d",x"30fe",x"2af5",x"3d32",x"368e",x"3c00",x"8000",x"0000",x"3732",x"2a26"),
(x"2af5",x"3d32",x"36fb",x"3c00",x"8000",x"0000",x"36f3",x"2a26",x"2af5",x"3ed3",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30d2",x"2af5",x"3d32",x"368e",x"3c00",x"8000",x"0000",x"3732",x"2a26"),
(x"2975",x"3ed3",x"36b2",x"3c00",x"8000",x"0000",x"3b75",x"396a",x"2975",x"3ed3",x"36d6",x"3c00",x"8000",x"0000",x"3b75",x"396e",x"2975",x"3ee9",x"36b2",x"3c00",x"8000",x"0000",x"3b81",x"396a"),
(x"2af5",x"3ed3",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a4e",x"2975",x"3ed3",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a48",x"2af5",x"3ee9",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a4e"),
(x"2af5",x"3ed3",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30d2",x"2af5",x"3d32",x"36fb",x"3c00",x"8000",x"0000",x"36f3",x"2a26",x"2af5",x"3ee9",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30fe"),
(x"2af5",x"3ee9",x"36b2",x"0000",x"bc00",x"0000",x"3b98",x"396e",x"2975",x"3ee9",x"36b2",x"0000",x"bc00",x"0000",x"3b9e",x"396e",x"2af5",x"3ee9",x"36d6",x"0000",x"bc00",x"0000",x"3b98",x"396a"),
(x"2af5",x"3ed3",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"39a5",x"2975",x"3ed3",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"399f",x"2af5",x"3ed3",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"39a5"),
(x"2af5",x"3ee9",x"36d6",x"0000",x"19f0",x"bc00",x"3b81",x"3a3e",x"2975",x"3ee9",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a3e",x"2af5",x"3ed3",x"36d6",x"0000",x"19f0",x"bc00",x"3b81",x"3a33"),
(x"b936",x"3d32",x"36fb",x"bc00",x"0000",x"0000",x"35f2",x"38f3",x"b936",x"3d32",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"38f3",x"b936",x"4062",x"368e",x"bc00",x"0000",x"0000",x"35dd",x"3a68"),
(x"2af5",x"3ee9",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30fe",x"2af5",x"4062",x"36fb",x"3c00",x"8000",x"0000",x"36f3",x"345d",x"2af5",x"4062",x"368e",x"3c00",x"8000",x"0000",x"3732",x"345d"),
(x"aaef",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3af7",x"3810",x"b858",x"4024",x"36d0",x"0000",x"bc00",x"0000",x"3a04",x"3810",x"b858",x"4024",x"36fb",x"0000",x"bc00",x"0000",x"3a04",x"3815"),
(x"b936",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3a0a",x"2af5",x"3d32",x"36fb",x"0000",x"bc00",x"0000",x"3bef",x"3b6a",x"2af5",x"3d32",x"368e",x"0000",x"bc00",x"0000",x"3bfe",x"3b6a"),
(x"b936",x"4062",x"36fb",x"0000",x"3c00",x"0000",x"39c2",x"397a",x"b936",x"4062",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"397a",x"2af5",x"4062",x"368e",x"0000",x"3c00",x"0000",x"39b3",x"3ada"),
(x"b863",x"3dc6",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3acc",x"b858",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3ac4",x"b936",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3a95"),
(x"b863",x"3dc6",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3acc",x"b857",x"3dbb",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3ac8",x"b858",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3ac4"),
(x"b862",x"401d",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3bb7",x"b858",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3bbc",x"b857",x"4023",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3bbb"),
(x"b862",x"401d",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3bb7",x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"b858",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3bbc"),
(x"b86c",x"3dde",x"36fb",x"0000",x"8000",x"3c00",x"39eb",x"3ad5",x"b863",x"3dc6",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3acc",x"b936",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3a95"),
(x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"b862",x"401d",x"36fb",x"0000",x"8000",x"3c00",x"39ed",x"3bb7",x"b86b",x"4016",x"36fb",x"0000",x"8000",x"3c00",x"39eb",x"3bb1"),
(x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"b86c",x"3dde",x"36fb",x"0000",x"8000",x"3c00",x"39eb",x"3ad5",x"b936",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3a95"),
(x"aa60",x"401e",x"36fb",x"0000",x"8000",x"3c00",x"3aaf",x"3bb7",x"aaef",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3bbc",x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea"),
(x"aa60",x"401e",x"36fb",x"0000",x"8000",x"3c00",x"3aaf",x"3bb7",x"aaef",x"4022",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3bba",x"aaef",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3bbc"),
(x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea",x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95",x"2243",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b39"),
(x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea",x"2243",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b39",x"20b0",x"3eef",x"36fb",x"0000",x"8000",x"3c00",x"3ac6",x"3b3b"),
(x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0",x"aa60",x"401e",x"36fb",x"0000",x"8000",x"3c00",x"3aaf",x"3bb7",x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea"),
(x"a0d7",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3abf",x"3b2b",x"a9ae",x"3dd7",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3ad3",x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0"),
(x"9e2f",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b39",x"995f",x"3ee2",x"36fb",x"0000",x"8000",x"3c00",x"3ac2",x"3b36",x"a0d7",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3abf",x"3b2b"),
(x"9e2f",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b39",x"9ac5",x"3ee4",x"36fb",x"0000",x"8000",x"3c00",x"3ac1",x"3b37",x"995f",x"3ee2",x"36fb",x"0000",x"8000",x"3c00",x"3ac2",x"3b36"),
(x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0",x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea",x"20b0",x"3eef",x"36fb",x"0000",x"8000",x"3c00",x"3ac6",x"3b3b"),
(x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0",x"20b0",x"3eef",x"36fb",x"0000",x"8000",x"3c00",x"3ac6",x"3b3b",x"1557",x"3ef2",x"36fb",x"0000",x"8000",x"3c00",x"3ac3",x"3b3c"),
(x"9e2f",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b39",x"a0d7",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3abf",x"3b2b",x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0"),
(x"a9a6",x"4015",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3bb0",x"1557",x"3ef2",x"36fb",x"0000",x"8000",x"3c00",x"3ac3",x"3b3c",x"9da8",x"3eee",x"36fb",x"0000",x"8000",x"3c00",x"3ac0",x"3b3b"),
(x"b936",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3a95",x"b858",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"39ef",x"3ac4",x"aaef",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3ac4"),
(x"b936",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"39c5",x"3bea",x"2af5",x"4062",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3bea",x"aaef",x"4024",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3bbc"),
(x"b858",x"3dae",x"36d0",x"0000",x"8000",x"3c00",x"35d9",x"3adb",x"b858",x"4024",x"36d0",x"0000",x"8000",x"3c00",x"35d9",x"3bfa",x"aaef",x"4024",x"36d0",x"0000",x"8000",x"3c00",x"3742",x"3bfa"),
(x"aaef",x"3dbd",x"36fb",x"bc00",x"0000",x"0000",x"3ae5",x"3546",x"aaef",x"3dae",x"36fb",x"bc00",x"0000",x"0000",x"3ae8",x"3545",x"aaef",x"3dae",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542"),
(x"aaef",x"3dae",x"36d0",x"bc00",x"0000",x"0000",x"3ae7",x"3542",x"aaef",x"3dd5",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545",x"aaef",x"3dc7",x"36e5",x"bc00",x"0000",x"0000",x"3ae4",x"3545"),
(x"b858",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3a05",x"3826",x"aaef",x"3dae",x"36d0",x"0000",x"3c00",x"0000",x"3af8",x"3826",x"aaef",x"3dae",x"36fb",x"0000",x"3c00",x"0000",x"3af8",x"3821"),
(x"aaef",x"4016",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"aaef",x"401e",x"36e4",x"ba1e",x"b322",x"38d5",x"351b",x"38d1",x"aa60",x"401e",x"36fb",x"b9bc",x"b304",x"394a",x"3521",x"38d1"),
(x"aaef",x"3dae",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3ac4",x"aaef",x"3dbd",x"36fb",x"0000",x"8000",x"3c00",x"3aad",x"3ac9",x"aa24",x"3dc9",x"36fb",x"0000",x"8000",x"3c00",x"3ab0",x"3ace"),
(x"aaef",x"4024",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"4016",x"36d7",x"bc00",x"0000",x"0000",x"3a9d",x"3546",x"aaef",x"3dd5",x"36d4",x"bc00",x"0000",x"0000",x"3ae1",x"3545"),
(x"aaef",x"401e",x"36e4",x"bc00",x"0000",x"0000",x"3a8d",x"354c",x"aaef",x"4016",x"36d7",x"bc00",x"0000",x"0000",x"3a9d",x"3546",x"aaef",x"4024",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542"),
(x"aaef",x"4024",x"36d0",x"bc00",x"0000",x"0000",x"3a80",x"3542",x"aaef",x"4022",x"36fb",x"bc00",x"0000",x"0000",x"3a83",x"3557",x"aaef",x"401e",x"36e4",x"bc00",x"0000",x"0000",x"3a8d",x"354c"),
(x"aaef",x"3dd5",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"aaef",x"4016",x"36d7",x"b94c",x"a074",x"39fd",x"3519",x"38c9",x"a9a6",x"4015",x"36fb",x"b96d",x"9af6",x"39e0",x"3525",x"38c8"),
(x"aaef",x"3dd5",x"36d4",x"b96e",x"1b2b",x"39df",x"3519",x"373e",x"a9ae",x"3dd7",x"36fb",x"b993",x"1c9b",x"39bd",x"3526",x"3740",x"aa24",x"3dc9",x"36fb",x"b988",x"33a8",x"3973",x"3523",x"3732"),
(x"b858",x"4024",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b857",x"4016",x"36d8",x"3bf1",x"15bc",x"afa2",x"3b3f",x"34eb",x"b857",x"401d",x"36e5",x"3bfe",x"2111",x"a780",x"3b41",x"34eb"),
(x"b857",x"4023",x"36fb",x"3bfe",x"276c",x"a4f7",x"3b42",x"34ec",x"b858",x"4024",x"36fb",x"3bf4",x"2eb8",x"0000",x"3b42",x"34eb",x"b858",x"4024",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9"),
(x"b857",x"3dc6",x"36dd",x"3bff",x"a074",x"a611",x"3aec",x"34f3",x"b857",x"3ddc",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed",x"b858",x"3dae",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9"),
(x"b858",x"3dae",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b857",x"3dbb",x"36fb",x"3bff",x"a3a0",x"a0dd",x"3ade",x"3501",x"b857",x"3dc6",x"36dd",x"3bff",x"a074",x"a611",x"3aec",x"34f3"),
(x"b858",x"4024",x"36d0",x"3a68",x"217a",x"b8ca",x"3b42",x"34e9",x"b858",x"3dae",x"36d0",x"bb8d",x"a187",x"b543",x"3ad3",x"34e9",x"b857",x"3ddc",x"36ca",x"39ed",x"90ea",x"b95f",x"3b04",x"34ed"),
(x"b857",x"3ddc",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b857",x"3dc6",x"36dd",x"3a1a",x"3321",x"38da",x"357e",x"38d0",x"b863",x"3dc6",x"36fb",x"3a1d",x"31d2",x"38f2",x"3587",x"38d0"),
(x"b857",x"4016",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b857",x"3ddc",x"36ca",x"3a15",x"1cb5",x"3931",x"357b",x"38c5",x"b86c",x"3dde",x"36fb",x"39b6",x"128d",x"3999",x"358a",x"38c4"),
(x"b857",x"4016",x"36d8",x"39b2",x"9dbc",x"399d",x"357b",x"373c",x"b86b",x"4016",x"36fb",x"3935",x"9d6d",x"3a12",x"3587",x"373c",x"b862",x"401d",x"36fb",x"394f",x"b2e4",x"39ba",x"3584",x"372e"),
(x"2163",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b2b",x"a9ae",x"3dd7",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3ad3",x"a0d7",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3abf",x"3b2b"),
(x"2163",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b2b",x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95",x"a9ae",x"3dd7",x"36fb",x"0000",x"8000",x"3c00",x"3ab1",x"3ad3"),
(x"2163",x"3ec3",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b2b",x"2243",x"3eea",x"36fb",x"0000",x"8000",x"3c00",x"3ac7",x"3b39",x"2af5",x"3d32",x"36fb",x"0000",x"8000",x"3c00",x"3ad8",x"3a95"),
(x"2af5",x"3d32",x"368e",x"0000",x"0000",x"bc00",x"3b35",x"30b7",x"2af5",x"4062",x"368e",x"0000",x"0000",x"bc00",x"3b35",x"290e",x"b936",x"4062",x"368e",x"0000",x"0000",x"bc00",x"3a79",x"290e"),
(x"9e2f",x"3eea",x"36fb",x"3b8f",x"3538",x"068d",x"3a18",x"3614",x"9e2f",x"3eea",x"36b4",x"3bef",x"3011",x"8000",x"3a18",x"3603",x"9ac5",x"3ee4",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603"),
(x"a0d7",x"3ec3",x"36fb",x"2460",x"3bff",x"0000",x"3b6d",x"3a51",x"a0d7",x"3ec3",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a51",x"2163",x"3ec3",x"36b4",x"2460",x"3bff",x"0000",x"3b77",x"3a47"),
(x"2243",x"3eea",x"36fb",x"bbcf",x"b2e8",x"0000",x"3a26",x"3614",x"2243",x"3eea",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603",x"20b0",x"3eef",x"36b4",x"b93c",x"ba0c",x"8000",x"3a23",x"3603"),
(x"9da8",x"3eee",x"36fb",x"3aa7",x"b870",x"0000",x"3a1b",x"3614",x"9da8",x"3eee",x"36b4",x"38fa",x"ba42",x"8000",x"3a1b",x"3603",x"9e2f",x"3eea",x"36b4",x"3bef",x"3011",x"8000",x"3a18",x"3603"),
(x"995f",x"3ee2",x"36fb",x"3bd4",x"b28e",x"0000",x"3a14",x"3614",x"995f",x"3ee2",x"36b4",x"3be8",x"b0e3",x"8000",x"3a14",x"3603",x"a0d7",x"3ec3",x"36b4",x"3bcb",x"b335",x"0000",x"3a04",x"3603"),
(x"20f3",x"3ee4",x"36fb",x"bbf6",x"2e14",x"0000",x"3a2a",x"3614",x"20f3",x"3ee4",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603",x"2243",x"3eea",x"36b4",x"bbf2",x"2f67",x"868d",x"3a26",x"3603"),
(x"1557",x"3ef2",x"36fb",x"332d",x"bbcb",x"0000",x"3a1f",x"3614",x"1557",x"3ef2",x"36b4",x"a8d6",x"bbfe",x"0000",x"3a1f",x"3603",x"9da8",x"3eee",x"36b4",x"38fa",x"ba42",x"8000",x"3a1b",x"3603"),
(x"9ac5",x"3ee4",x"36fb",x"3b7d",x"359e",x"0000",x"3a15",x"3614",x"9ac5",x"3ee4",x"36b4",x"3b3f",x"36c6",x"0000",x"3a15",x"3603",x"995f",x"3ee2",x"36b4",x"3be8",x"b0e3",x"8000",x"3a14",x"3603"),
(x"2163",x"3ec3",x"36fb",x"bbff",x"a6cf",x"0000",x"3a3b",x"3614",x"2163",x"3ec3",x"36b4",x"bbff",x"a6cf",x"0000",x"3a3b",x"3603",x"20f3",x"3ee4",x"36b4",x"bbff",x"2231",x"0000",x"3a2a",x"3603"),
(x"20b0",x"3eef",x"36fb",x"b727",x"bb27",x"868d",x"3a23",x"3614",x"20b0",x"3eef",x"36b4",x"b93c",x"ba0c",x"8000",x"3a23",x"3603",x"1557",x"3ef2",x"36b4",x"a8d6",x"bbfe",x"0000",x"3a1f",x"3603"),
(x"9da8",x"3eee",x"36b4",x"0000",x"8000",x"3c00",x"3b63",x"3a1a",x"1557",x"3ef2",x"36b4",x"0000",x"8000",x"3c00",x"3b61",x"3a16",x"9e2f",x"3eea",x"36b4",x"0000",x"8000",x"3c00",x"3b65",x"3a1a"),
(x"20b0",x"3eef",x"36b4",x"0000",x"8000",x"3c00",x"3b62",x"3a12",x"9ac5",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a18",x"1557",x"3ef2",x"36b4",x"0000",x"8000",x"3c00",x"3b61",x"3a16"),
(x"2243",x"3eea",x"36b4",x"0000",x"8000",x"3c00",x"3b65",x"3a11",x"20f3",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a12",x"20b0",x"3eef",x"36b4",x"0000",x"8000",x"3c00",x"3b62",x"3a12"),
(x"2163",x"3ec3",x"36b4",x"0000",x"8000",x"3c00",x"3b79",x"3a11",x"995f",x"3ee2",x"36b4",x"0000",x"8000",x"3c00",x"3b69",x"3a18",x"20f3",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a12"),
(x"a0d7",x"3ec3",x"36b4",x"0000",x"8000",x"3c00",x"3b79",x"3a1b",x"995f",x"3ee2",x"36b4",x"0000",x"8000",x"3c00",x"3b69",x"3a18",x"2163",x"3ec3",x"36b4",x"0000",x"8000",x"3c00",x"3b79",x"3a11"),
(x"20f3",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a12",x"9ac5",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a18",x"20b0",x"3eef",x"36b4",x"0000",x"8000",x"3c00",x"3b62",x"3a12"),
(x"9e2f",x"3eea",x"36b4",x"0000",x"8000",x"3c00",x"3b65",x"3a1a",x"1557",x"3ef2",x"36b4",x"0000",x"8000",x"3c00",x"3b61",x"3a16",x"9ac5",x"3ee4",x"36b4",x"0000",x"8000",x"3c00",x"3b68",x"3a18"),
(x"2af5",x"3ee9",x"36b2",x"3c00",x"8000",x"0000",x"371d",x"30fe",x"2af5",x"4062",x"368e",x"3c00",x"8000",x"0000",x"3732",x"345d",x"2af5",x"3d32",x"368e",x"3c00",x"8000",x"0000",x"3732",x"2a26"),
(x"2af5",x"3ed3",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30d2",x"2af5",x"3ed3",x"36b2",x"3c00",x"8000",x"0000",x"371d",x"30d2",x"2af5",x"3d32",x"368e",x"3c00",x"8000",x"0000",x"3732",x"2a26"),
(x"2975",x"3ed3",x"36d6",x"3c00",x"8000",x"0000",x"3b75",x"396e",x"2975",x"3ee9",x"36d6",x"3c00",x"8000",x"0000",x"3b81",x"396e",x"2975",x"3ee9",x"36b2",x"3c00",x"8000",x"0000",x"3b81",x"396a"),
(x"2975",x"3ed3",x"36b2",x"0000",x"96f6",x"3c00",x"3b07",x"3a48",x"2975",x"3ee9",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a48",x"2af5",x"3ee9",x"36b2",x"0000",x"96f6",x"3c00",x"3afc",x"3a4e"),
(x"2af5",x"3d32",x"36fb",x"3c00",x"8000",x"0000",x"36f3",x"2a26",x"2af5",x"4062",x"36fb",x"3c00",x"8000",x"0000",x"36f3",x"345d",x"2af5",x"3ee9",x"36d6",x"3c00",x"8000",x"0000",x"3709",x"30fe"),
(x"2975",x"3ee9",x"36b2",x"0000",x"bc00",x"0000",x"3b9e",x"396e",x"2975",x"3ee9",x"36d6",x"0000",x"bc00",x"0000",x"3b9e",x"396a",x"2af5",x"3ee9",x"36d6",x"0000",x"bc00",x"0000",x"3b98",x"396a"),
(x"2975",x"3ed3",x"36d6",x"0000",x"3c00",x"0000",x"3b85",x"399f",x"2975",x"3ed3",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"399f",x"2af5",x"3ed3",x"36b2",x"0000",x"3c00",x"0000",x"3b80",x"39a5"),
(x"2975",x"3ee9",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a3e",x"2975",x"3ed3",x"36d6",x"0000",x"19f0",x"bc00",x"3b87",x"3a33",x"2af5",x"3ed3",x"36d6",x"0000",x"19f0",x"bc00",x"3b81",x"3a33"),
(x"b931",x"4036",x"3710",x"bbe9",x"26a1",x"309e",x"39b2",x"33ca",x"b930",x"4041",x"3710",x"bbeb",x"2604",x"3075",x"39c5",x"33c0",x"b92b",x"4036",x"3732",x"bb64",x"243f",x"361b",x"39b1",x"33aa"),
(x"b92b",x"4036",x"3732",x"bb64",x"243f",x"361b",x"39b1",x"33aa",x"b92a",x"4041",x"3733",x"bb1e",x"2518",x"3748",x"39c4",x"339f",x"b924",x"4036",x"3749",x"ba3b",x"2680",x"3902",x"39b0",x"3392"),
(x"b924",x"4036",x"3749",x"ba3b",x"2680",x"3902",x"39b0",x"3392",x"b922",x"4041",x"3748",x"b86c",x"29d9",x"3aa7",x"39c4",x"3388",x"b91f",x"4036",x"374e",x"ac96",x"29b2",x"3bf8",x"39b0",x"3387"),
(x"b91f",x"4036",x"374e",x"ac96",x"29b2",x"3bf8",x"39b0",x"3387",x"b91b",x"4041",x"3749",x"3594",x"2b76",x"3b7b",x"39c3",x"337b",x"b918",x"4036",x"374b",x"38f0",x"29d6",x"3a48",x"39b0",x"337b"),
(x"b907",x"4042",x"3713",x"2f5f",x"3bdb",x"30c1",x"3b21",x"38a0",x"b913",x"4041",x"373b",x"381d",x"3a67",x"34eb",x"3b1c",x"3899",x"b90e",x"4042",x"370e",x"3754",x"3ae5",x"32eb",x"3b1f",x"38a1"),
(x"b91b",x"4042",x"374a",x"3544",x"b37e",x"3b51",x"3b18",x"3896",x"b913",x"4042",x"373a",x"3ae3",x"2b4b",x"380a",x"3b1b",x"3899",x"b91b",x"4041",x"3749",x"382b",x"a439",x"3ad3",x"3b1a",x"3895"),
(x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e",x"b906",x"4036",x"3710",x"2e12",x"a673",x"3bf6",x"39b0",x"333e",x"b90c",x"4036",x"3724",x"3af5",x"1a59",x"37e2",x"39b0",x"3352"),
(x"b90f",x"404d",x"3727",x"3bc1",x"a907",x"33c0",x"3bfb",x"39a3",x"b90d",x"404d",x"3711",x"3be1",x"a6cf",x"3179",x"3bfb",x"399f",x"b90e",x"4042",x"370e",x"3bcb",x"a949",x"330f",x"3bea",x"399f"),
(x"b91a",x"404d",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"39ab",x"b913",x"404d",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"39a7",x"b91b",x"4042",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"39ac"),
(x"b922",x"404d",x"3751",x"a111",x"aa52",x"3bfd",x"3bfc",x"39af",x"b91a",x"404d",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"39ab",x"b924",x"4043",x"374d",x"af62",x"aa90",x"3bef",x"3bec",x"39af"),
(x"b92b",x"4043",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"39b3",x"b928",x"404d",x"374d",x"b867",x"a907",x"3aab",x"3bfc",x"39b1",x"b924",x"4043",x"374d",x"af62",x"aa90",x"3bef",x"3bec",x"39af"),
(x"b930",x"4043",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"39b6",x"b92f",x"404d",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"39b5",x"b92b",x"4043",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"39b3"),
(x"b938",x"4042",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"39be",x"b935",x"404d",x"3725",x"bb50",x"a63f",x"3678",x"3bfb",x"39ba",x"b930",x"4043",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"39b6"),
(x"b935",x"404d",x"3725",x"bb50",x"a63f",x"3678",x"3bfb",x"39ba",x"b938",x"4042",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"39be",x"b93a",x"404d",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3bfb",x"39bf"),
(x"b938",x"4042",x"3710",x"b678",x"bb4d",x"2af6",x"3b19",x"3884",x"b930",x"4043",x"3738",x"b75b",x"bae5",x"32d3",x"3b16",x"388d",x"b930",x"4041",x"3710",x"b700",x"bb23",x"2f0f",x"3b1b",x"3887"),
(x"b912",x"4036",x"373c",x"3aea",x"2832",x"3802",x"39b0",x"336a",x"b918",x"4036",x"374b",x"38f0",x"29d6",x"3a48",x"39b0",x"337b",x"b913",x"4041",x"373b",x"3aa1",x"2559",x"3879",x"39c3",x"3369"),
(x"b924",x"4043",x"374d",x"b1ce",x"b808",x"3ac1",x"3b16",x"3893",x"b91b",x"4042",x"374a",x"3544",x"b37e",x"3b51",x"3b18",x"3896",x"b922",x"4041",x"3748",x"b511",x"b92e",x"398b",x"3b18",x"3893"),
(x"b924",x"4043",x"374d",x"b1ce",x"b808",x"3ac1",x"3b16",x"3893",x"b922",x"4041",x"3748",x"b511",x"b92e",x"398b",x"3b18",x"3893",x"b92b",x"4043",x"3744",x"b779",x"ba1b",x"3724",x"3b16",x"388f"),
(x"b92a",x"4041",x"3733",x"b800",x"ba99",x"3435",x"3b19",x"388d",x"b930",x"4043",x"3738",x"b75b",x"bae5",x"32d3",x"3b16",x"388d",x"b92b",x"4043",x"3744",x"b779",x"ba1b",x"3724",x"3b16",x"388f"),
(x"b92a",x"404d",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3827",x"b935",x"404d",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3821",x"b931",x"404d",x"3710",x"b3e2",x"3bbf",x"28bf",x"3b1e",x"3820"),
(x"b925",x"404d",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"382b",x"b92f",x"404d",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3826",x"b92a",x"404d",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3827"),
(x"b920",x"404d",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"382d",x"b928",x"404d",x"374d",x"b4d8",x"3aa1",x"3784",x"3b25",x"382a",x"b925",x"404d",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"382b"),
(x"b920",x"404d",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"382d",x"b922",x"404d",x"3751",x"9ac2",x"39ac",x"39a3",x"3b24",x"382d",x"b928",x"404d",x"374d",x"b4d8",x"3aa1",x"3784",x"3b25",x"382a"),
(x"b919",x"404e",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"382f",x"b91a",x"404d",x"374d",x"35fb",x"37c0",x"3a53",x"3b22",x"3830",x"b920",x"404d",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"382d"),
(x"b913",x"404e",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3831",x"b913",x"404d",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3832",x"b919",x"404e",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"382f"),
(x"b90b",x"404d",x"371c",x"391d",x"b988",x"3561",x"3b19",x"3835",x"b90f",x"404d",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3835",x"b913",x"404e",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3831"),
(x"b90b",x"404d",x"371c",x"391d",x"b988",x"3561",x"3b19",x"3835",x"b90d",x"404d",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"3838",x"b90f",x"404d",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3835"),
(x"b906",x"404d",x"3713",x"2edc",x"bb7b",x"3565",x"3b16",x"3836",x"b90d",x"404d",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"3838",x"b90b",x"404d",x"371c",x"391d",x"b988",x"3561",x"3b19",x"3835"),
(x"b90e",x"4042",x"370e",x"b4eb",x"a6e9",x"3b9c",x"39c4",x"334b",x"b90d",x"404d",x"3711",x"b36d",x"a40b",x"3bc7",x"39d6",x"3349",x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e"),
(x"b931",x"4059",x"3710",x"bbfe",x"a4d0",x"28c6",x"39ea",x"33c9",x"b92f",x"4059",x"372b",x"bbac",x"a891",x"347c",x"39eb",x"33b1",x"b931",x"404d",x"3710",x"bbea",x"a7ae",x"307d",x"39d7",x"33c4"),
(x"b92a",x"404d",x"3739",x"bb13",x"a8dd",x"3771",x"39d7",x"339e",x"b92f",x"4059",x"372b",x"bbac",x"a891",x"347c",x"39eb",x"33b1",x"b92c",x"4059",x"373a",x"baa5",x"a5fd",x"3872",x"39eb",x"33a3"),
(x"b925",x"404d",x"3746",x"b918",x"a84d",x"3a28",x"39d8",x"338e",x"b92a",x"404d",x"3739",x"bb13",x"a8dd",x"3771",x"39d7",x"339e",x"b925",x"4059",x"3749",x"b926",x"a7c8",x"3a1d",x"39eb",x"3391"),
(x"b91f",x"4059",x"374f",x"a812",x"a959",x"3bfd",x"39eb",x"3384",x"b920",x"404d",x"374b",x"b451",x"a960",x"3bb2",x"39d8",x"3385",x"b925",x"4059",x"3749",x"b926",x"a7c8",x"3a1d",x"39eb",x"3391"),
(x"b918",x"4059",x"374b",x"38ec",x"a7f6",x"3a4c",x"39eb",x"3378",x"b919",x"404e",x"3749",x"3647",x"a97a",x"3b59",x"39d8",x"3379",x"b91f",x"4059",x"374f",x"a812",x"a959",x"3bfd",x"39eb",x"3384"),
(x"b911",x"4059",x"373c",x"3ac9",x"a6b5",x"383a",x"39eb",x"3366",x"b913",x"404e",x"373e",x"3ac8",x"a7bb",x"383c",x"39d8",x"336a",x"b918",x"4059",x"374b",x"38ec",x"a7f6",x"3a4c",x"39eb",x"3378"),
(x"b90b",x"404d",x"371c",x"3aa9",x"a818",x"386b",x"39d7",x"334a",x"b913",x"404e",x"373e",x"3ac8",x"a7bb",x"383c",x"39d8",x"336a",x"b90b",x"4059",x"3722",x"3b0f",x"a82c",x"3781",x"39ea",x"334c"),
(x"b906",x"404d",x"3713",x"29ab",x"208e",x"3bfd",x"39d7",x"333d",x"b90b",x"404d",x"371c",x"3aa9",x"a818",x"386b",x"39d7",x"334a",x"b907",x"4059",x"3718",x"38f7",x"a86d",x"3a44",x"39eb",x"3340"),
(x"b135",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"24c1",x"b116",x"404a",x"3710",x"0000",x"8000",x"3c00",x"39d1",x"2450",x"b135",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"24c1"),
(x"b135",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"24c1",x"b135",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"24c1",x"b161",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"255f"),
(x"b161",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"255f",x"b161",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"255f",x"b1a1",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2642"),
(x"b1c1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"26b3",x"b1a1",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2642",x"b1c1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"26b3"),
(x"b1c1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"26b3",x"b1c1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"26b3",x"b1fd",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"278b"),
(x"b22d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"281a",x"b1fd",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"278b",x"b22d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"281a"),
(x"b261",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"2878",x"b22d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"281a",x"b261",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39be",x"2878"),
(x"b2aa",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"28fa",x"b261",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"2878",x"b2aa",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"28fa"),
(x"b2aa",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"28fa",x"b2aa",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"28fa",x"b2d6",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2949"),
(x"b326",x"404b",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"29d7",x"b2d6",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2949",x"b326",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"29d7"),
(x"b34f",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"2a20",x"b326",x"404b",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"29d7",x"b34f",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2a20"),
(x"b451",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2c3f",x"b50c",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2d8d",x"b451",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2c3f"),
(x"b451",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2c3f",x"b451",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2c3f",x"b441",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2c23"),
(x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b",x"b441",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2c23",x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b"),
(x"b34f",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2a20",x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b",x"b34f",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"2a20"),
(x"b413",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"2ba0",x"b40b",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2b83",x"b413",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2ba0"),
(x"b413",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2ba0",x"b3f4",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2b47",x"b409",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2b7d"),
(x"b409",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2b7d",x"b3d2",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"2b0a",x"b407",x"4052",x"3710",x"0000",x"8000",x"3c00",x"39df",x"2b76"),
(x"b3f4",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2b47",x"b40b",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2b83",x"b413",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2ba0"),
(x"b3d2",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2b0a",x"b3f4",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2b47",x"b409",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2b7d"),
(x"b3a5",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"2ab9",x"b3d2",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2b0a",x"b407",x"403d",x"3710",x"8000",x"0cea",x"3c00",x"39bb",x"2b76"),
(x"b368",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2a4d",x"b3a5",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"2ab9",x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b"),
(x"b407",x"4052",x"3710",x"0000",x"8000",x"3c00",x"39df",x"2b76",x"b3a5",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2ab9",x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b"),
(x"b368",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2a4d",x"b351",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2a27",x"b340",x"403d",x"3710",x"0000",x"8000",x"3c00",x"39bb",x"2a0d"),
(x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b",x"b351",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2a24",x"b34f",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"2a20"),
(x"b50c",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2d8d",x"b50c",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2d8d",x"b526",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2dbb"),
(x"b5ce",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2ee7",x"b62a",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2f8b",x"b5ce",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ee7"),
(x"b5ce",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2ee7",x"b5ce",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ee7",x"b5bd",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2ec9"),
(x"b5a1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2e97",x"b5bd",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2ec9",x"b5a1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2e97"),
(x"b5a1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2e97",x"b5a1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2e97",x"b581",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"2e5e"),
(x"b568",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2e30",x"b581",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"2e5e",x"b568",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2e30"),
(x"b52b",x"405a",x"3710",x"0000",x"8000",x"3c00",x"39ed",x"2dc4",x"b50d",x"405b",x"3710",x"0000",x"8000",x"3c00",x"39ee",x"2d8e",x"b4f5",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"2d63"),
(x"b544",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2df0",x"b52b",x"405a",x"3710",x"0000",x"8000",x"3c00",x"39ed",x"2dc4",x"b4f2",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2d5e"),
(x"b52b",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ad",x"2dc4",x"b4f5",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"2d63",x"b50d",x"4034",x"3710",x"0000",x"8000",x"3c00",x"39ac",x"2d8e"),
(x"b544",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2df0",x"b4f2",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2d5e",x"b52b",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ad",x"2dc4"),
(x"b558",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2e14",x"b568",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b0",x"2e32",x"b575",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2e47"),
(x"b544",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2df0",x"b558",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2e14",x"b569",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"2e33"),
(x"b575",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e7",x"2e49",x"b568",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39ea",x"2e32",x"b575",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e4",x"2e47"),
(x"b575",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e4",x"2e47",x"b558",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2e14",x"b569",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"2e33"),
(x"b4d8",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"2d2f",x"b4e1",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2d3f",x"b4da",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"2d33"),
(x"b51a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"2da6",x"b4e1",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39be",x"2d3f",x"b4da",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"2d33"),
(x"b528",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"2dbf",x"b51a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"2da6",x"b4f2",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2d5e"),
(x"b4da",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"2d33",x"b51a",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"2da6",x"b4f2",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2d5e"),
(x"b4f2",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2d5e",x"b528",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2dbf",x"b544",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2df0"),
(x"b4f2",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2d5e",x"b544",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2df0",x"b528",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"2dbf"),
(x"b569",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"2e33",x"b528",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2dbf",x"b568",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2e30"),
(x"b52c",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2dc5",x"b528",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"2dbf",x"b568",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2e30"),
(x"b526",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2dbb",x"b526",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2dbb",x"b52c",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2dc5"),
(x"b568",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2e30",x"b52c",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2dc5",x"b568",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2e30"),
(x"b63d",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2fac",x"b63d",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2fac",x"b62a",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2f8b"),
(x"b669",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2ffc",x"b669",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2ffc",x"b63d",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2fac"),
(x"b721",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30a2",x"b721",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30a2",x"b669",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2ffc"),
(x"b72d",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30ad",x"b721",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30a2",x"b72d",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30ad"),
(x"b794",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"3109",x"b794",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"3109",x"b7c0",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"3130"),
(x"b77a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"30f1",x"b794",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"3109",x"b77a",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"30f1"),
(x"b776",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"30ed",x"b77a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"30f1",x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed"),
(x"b776",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"30ed",x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed",x"b72d",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30ad"),
(x"b705",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3088",x"b6fb",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"3080",x"b6f1",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3076"),
(x"b73e",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ae",x"30bc",x"b721",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"30a2",x"b705",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3088"),
(x"b705",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3088",x"b6f1",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3076",x"b6fb",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"3080"),
(x"b73e",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39ec",x"30bc",x"b705",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3088",x"b721",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"30a2"),
(x"b783",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"30f9",x"b73e",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39ec",x"30bc",x"b72e",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"30ae"),
(x"b783",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"30f9",x"b72e",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"30ae",x"b73e",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ae",x"30bc"),
(x"b7a4",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"3117",x"b7c7",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3135",x"b7bd",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"312d"),
(x"b7c7",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e4",x"3136",x"b7c7",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3135",x"b7bd",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"312d"),
(x"b7bd",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"312d",x"b7a4",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"3117",x"b7a8",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"311a"),
(x"b783",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"30f9",x"b7a4",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"3117",x"b7a8",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"311a"),
(x"b72d",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30ad",x"b72e",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"30ae",x"b776",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"30ed"),
(x"b77b",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"30f2",x"b72e",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"30ae",x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed"),
(x"b783",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"30f9",x"b77b",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"30f2",x"b72e",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"30ae"),
(x"b77b",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"30f2",x"b783",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"30f9",x"b72e",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"30ae"),
(x"b77b",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"30f2",x"b783",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"30f9",x"b790",x"403d",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"3107"),
(x"b7a8",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"311a",x"b783",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"30f9",x"b790",x"4052",x"3710",x"0000",x"8000",x"3c00",x"39de",x"3107"),
(x"b801",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"316b",x"b801",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"316b",x"b7c0",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"3130"),
(x"b820",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"31a2",x"b801",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"316b",x"b820",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"31a2"),
(x"b83a",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"31d0",x"b83a",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"31d0",x"b820",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"31a2"),
(x"b84a",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"31ed",x"b84a",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"31ed",x"b83a",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"31d0"),
(x"b85e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3211",x"b85e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3211",x"b84a",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"31ed"),
(x"b865",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"321d",x"b85e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3211",x"b865",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"321d"),
(x"b867",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"3222",x"b867",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"3222",x"b865",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"321d"),
(x"b86e",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"322d",x"b867",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"3222",x"b86e",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"322d"),
(x"b87d",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"3248",x"b87d",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"3248",x"b86e",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"322d"),
(x"b88f",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3269",x"b88f",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3269",x"b87d",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"3248"),
(x"b89e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3284",x"b88f",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3269",x"b89e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3284"),
(x"b8a3",x"4037",x"3710",x"2081",x"9ea7",x"3bff",x"39b1",x"328d",x"b8a3",x"4058",x"3710",x"2160",x"1cd0",x"3bff",x"39e9",x"328d",x"b89e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3284"),
(x"b906",x"404d",x"3713",x"29ab",x"208e",x"3bfd",x"39d7",x"333d",x"b8a3",x"4058",x"3710",x"2160",x"1cd0",x"3bff",x"39e9",x"328d",x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e"),
(x"b907",x"4059",x"3718",x"38f7",x"a86d",x"3a44",x"39eb",x"3340",x"b8ff",x"4059",x"3710",x"2904",x"26d5",x"3bfd",x"39eb",x"3331",x"b906",x"404d",x"3713",x"29ab",x"208e",x"3bfd",x"39d7",x"333d"),
(x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e",x"b8a3",x"4037",x"3710",x"2081",x"9ea7",x"3bff",x"39b1",x"328d",x"b906",x"4036",x"3710",x"2e12",x"a673",x"3bf6",x"39b0",x"333e"),
(x"b911",x"4059",x"373c",x"2504",x"3bff",x"2111",x"3a1b",x"3ba6",x"b918",x"4059",x"374b",x"270a",x"3bfd",x"287a",x"3a18",x"3ba9",x"b925",x"4059",x"3749",x"257a",x"3bfd",x"28f7",x"3a18",x"3bae"),
(x"b90b",x"4059",x"3722",x"2773",x"3bfe",x"22dc",x"3a1f",x"3ba4",x"b911",x"4059",x"373c",x"2504",x"3bff",x"2111",x"3a1b",x"3ba6",x"b92c",x"4059",x"373a",x"25e9",x"3bff",x"17c8",x"3a1b",x"3bb1"),
(x"b907",x"4059",x"3718",x"25bc",x"3bfe",x"2673",x"3a21",x"3ba2",x"b90b",x"4059",x"3722",x"2773",x"3bfe",x"22dc",x"3a1f",x"3ba4",x"b92f",x"4059",x"372b",x"26c2",x"3bfe",x"24a2",x"3a1e",x"3bb2"),
(x"b8ff",x"4059",x"3710",x"257a",x"3bff",x"15bc",x"3a23",x"3b9f",x"b907",x"4059",x"3718",x"25bc",x"3bfe",x"2673",x"3a21",x"3ba2",x"b931",x"4059",x"3710",x"2418",x"3bff",x"1a24",x"3a23",x"3bb3"),
(x"b912",x"4036",x"373c",x"184d",x"bbff",x"26c8",x"3a0f",x"3ba4",x"b924",x"4036",x"3749",x"1ef6",x"bbff",x"23ef",x"3a12",x"3bab",x"b918",x"4036",x"374b",x"2511",x"bbff",x"224c",x"3a12",x"3ba6"),
(x"b90c",x"4036",x"3724",x"9e3f",x"bbff",x"a025",x"3a0b",x"3ba2",x"b92b",x"4036",x"3732",x"9cd0",x"bc00",x"1bc8",x"3a0d",x"3bae",x"b912",x"4036",x"373c",x"184d",x"bbff",x"26c8",x"3a0f",x"3ba4"),
(x"b906",x"4036",x"3710",x"2546",x"bbff",x"9624",x"3a07",x"3b9f",x"b931",x"4036",x"3710",x"9ec2",x"bc00",x"9da1",x"3a07",x"3bb0",x"b90c",x"4036",x"3724",x"9e3f",x"bbff",x"a025",x"3a0b",x"3ba2"),
(x"b1fd",x"403f",x"3710",x"375d",x"bb1a",x"0000",x"3a5a",x"3b8e",x"b1fd",x"403f",x"36da",x"35da",x"bb72",x"0000",x"3a50",x"3b8e",x"b22d",x"403e",x"3710",x"2c28",x"bbfb",x"0000",x"3a5a",x"3b93"),
(x"b6fb",x"403e",x"3710",x"37ed",x"3af2",x"0000",x"3a7c",x"3ad4",x"b6fb",x"403e",x"36da",x"38e1",x"3a57",x"0000",x"3a72",x"3ad4",x"b6ef",x"403c",x"3710",x"3b57",x"3658",x"8000",x"3a7c",x"3ad8"),
(x"b63d",x"404e",x"3710",x"affc",x"3bf0",x"0000",x"3a96",x"3b47",x"b63d",x"404e",x"36da",x"ab45",x"3bfc",x"0000",x"3a8b",x"3b47",x"b62a",x"404d",x"3710",x"2fbb",x"3bf1",x"0000",x"3a96",x"3b4a"),
(x"b1c1",x"4041",x"3710",x"367f",x"bb4f",x"0000",x"3a5a",x"3b87",x"b1c1",x"4041",x"36da",x"37bc",x"bb00",x"0000",x"3a50",x"3b87",x"b1fd",x"403f",x"3710",x"375d",x"bb1a",x"0000",x"3a5a",x"3b8e"),
(x"b906",x"4036",x"3710",x"2546",x"bbff",x"9624",x"3a07",x"3b9f",x"b906",x"4036",x"36da",x"2273",x"bbff",x"0000",x"39fd",x"3b9f",x"b931",x"4036",x"3710",x"9ec2",x"bc00",x"9da1",x"3a07",x"3bb0"),
(x"b721",x"4040",x"3710",x"37a6",x"3b06",x"8000",x"3a7c",x"3acc",x"b721",x"4040",x"36da",x"3711",x"3b2d",x"0000",x"3a72",x"3acc",x"b6fb",x"403e",x"3710",x"37ed",x"3af2",x"0000",x"3a7c",x"3ad4"),
(x"b575",x"4055",x"3710",x"ba67",x"b8cb",x"0000",x"3a96",x"3b77",x"b575",x"4055",x"36da",x"bb59",x"b650",x"8000",x"3a8b",x"3b77",x"b575",x"4056",x"3710",x"bb97",x"350c",x"8000",x"3a96",x"3b79"),
(x"b1a1",x"4042",x"3710",x"2ede",x"bbf4",x"0000",x"3a5a",x"3b84",x"b1a1",x"4042",x"36da",x"314f",x"bbe3",x"0000",x"3a50",x"3b84",x"b1c1",x"4041",x"3710",x"367f",x"bb4f",x"0000",x"3a5a",x"3b87"),
(x"b72e",x"4041",x"3710",x"3b4f",x"367e",x"8000",x"3a7c",x"3ac9",x"b72e",x"4041",x"36da",x"39a7",x"39a9",x"0000",x"3a72",x"3ac9",x"b721",x"4040",x"3710",x"37a6",x"3b06",x"8000",x"3a7c",x"3acc"),
(x"b62a",x"404d",x"3710",x"2fbb",x"3bf1",x"0000",x"3a96",x"3b4a",x"b62a",x"404d",x"36da",x"303b",x"3bed",x"8000",x"3a8b",x"3b4a",x"b5ce",x"404c",x"3710",x"2f26",x"3bf3",x"0000",x"3a96",x"3b5c"),
(x"b161",x"4042",x"3710",x"3407",x"bbbd",x"8000",x"3a5a",x"3b7e",x"b161",x"4042",x"36da",x"30d8",x"bbe8",x"8000",x"3a50",x"3b7e",x"b1a1",x"4042",x"3710",x"2ede",x"bbf4",x"0000",x"3a5a",x"3b84"),
(x"b72d",x"4042",x"3710",x"3778",x"bb13",x"0000",x"3a7c",x"3ac8",x"b72d",x"4042",x"36da",x"3a45",x"b8f8",x"0000",x"3a72",x"3ac8",x"b72e",x"4041",x"3710",x"3b4f",x"367e",x"8000",x"3a7c",x"3ac9"),
(x"b5ce",x"404c",x"3710",x"2f26",x"3bf3",x"0000",x"3a96",x"3b5c",x"b5ce",x"404c",x"36da",x"2ae9",x"3bfc",x"8000",x"3a8b",x"3b5c",x"b5bd",x"404c",x"3710",x"b559",x"3b8a",x"0000",x"3a96",x"3b5f"),
(x"b135",x"4043",x"3710",x"3934",x"ba13",x"0000",x"3a5a",x"3b7a",x"b135",x"4043",x"36da",x"3822",x"bad9",x"8000",x"3a50",x"3b7a",x"b161",x"4042",x"3710",x"3407",x"bbbd",x"8000",x"3a5a",x"3b7e"),
(x"b721",x"4042",x"3710",x"0cea",x"bc00",x"0000",x"3a4c",x"3bad",x"b721",x"4042",x"36da",x"2560",x"bbff",x"8000",x"3a42",x"3bad",x"b72d",x"4042",x"3710",x"3778",x"bb13",x"0000",x"3a4c",x"3bb0"),
(x"b5bd",x"404c",x"3710",x"b559",x"3b8a",x"0000",x"3a96",x"3b5f",x"b5bd",x"404c",x"36da",x"b6e1",x"3b38",x"0000",x"3a8b",x"3b5f",x"b5a1",x"404e",x"3710",x"b72d",x"3b26",x"8000",x"3a96",x"3b65"),
(x"b93a",x"404d",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"381d",x"b93a",x"404d",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"3816",x"b931",x"404d",x"3710",x"b3e2",x"3bbf",x"28bf",x"3b1e",x"3820"),
(x"b116",x"4045",x"3710",x"3bdf",x"b1b0",x"0000",x"3a5a",x"3b75",x"b116",x"4045",x"36da",x"3b51",x"b675",x"8000",x"3a50",x"3b75",x"b135",x"4043",x"3710",x"3934",x"ba13",x"0000",x"3a5a",x"3b7a"),
(x"b568",x"4037",x"3710",x"b810",x"bae4",x"0000",x"3a4c",x"3b48",x"b568",x"4037",x"36da",x"b919",x"ba29",x"0000",x"3a42",x"3b48",x"b575",x"4038",x"3710",x"bab5",x"b85c",x"8000",x"3a4c",x"3b4c"),
(x"b5a1",x"404e",x"3710",x"b72d",x"3b26",x"8000",x"3a96",x"3b65",x"b5a1",x"404e",x"36da",x"b67b",x"3b50",x"0000",x"3a8b",x"3b65",x"b581",x"4050",x"3710",x"b794",x"3b0b",x"0000",x"3a96",x"3b6c"),
(x"b669",x"4042",x"3710",x"abae",x"bbfc",x"0000",x"3a4c",x"3b89",x"b669",x"4042",x"36da",x"a65f",x"bbff",x"0000",x"3a42",x"3b89",x"b721",x"4042",x"3710",x"0cea",x"bc00",x"0000",x"3a4c",x"3bad"),
(x"b581",x"4050",x"3710",x"b794",x"3b0b",x"0000",x"3a96",x"3b6c",x"b581",x"4050",x"36da",x"b89f",x"3a87",x"0000",x"3a8b",x"3b6c",x"b568",x"4053",x"3710",x"b9f3",x"3958",x"0000",x"3a96",x"3b72"),
(x"b8a3",x"4037",x"3710",x"2a1e",x"bbfd",x"0000",x"3a07",x"3b78",x"b8a3",x"4037",x"36da",x"2850",x"bbfe",x"8000",x"39fd",x"3b78",x"b906",x"4036",x"3710",x"2546",x"bbff",x"9624",x"3a07",x"3b9f"),
(x"b63d",x"4041",x"3710",x"ab45",x"bbfc",x"0000",x"3a4c",x"3b80",x"b63d",x"4041",x"36da",x"affc",x"bbf0",x"8000",x"3a42",x"3b80",x"b669",x"4042",x"3710",x"abae",x"bbfc",x"0000",x"3a4c",x"3b89"),
(x"b568",x"4058",x"3710",x"b919",x"3a29",x"0000",x"3a96",x"3b7d",x"b568",x"4058",x"36da",x"b810",x"3ae4",x"8000",x"3a8b",x"3b7d",x"b558",x"4059",x"3710",x"b3cc",x"3bc2",x"8000",x"3a96",x"3b80"),
(x"b62a",x"4041",x"3710",x"303a",x"bbed",x"0000",x"3a4c",x"3b7c",x"b62a",x"4041",x"36da",x"2fb9",x"bbf1",x"0000",x"3a42",x"3b7c",x"b63d",x"4041",x"3710",x"ab45",x"bbfc",x"0000",x"3a4c",x"3b80"),
(x"b558",x"4059",x"3710",x"b3cc",x"3bc2",x"8000",x"3a96",x"3b80",x"b558",x"4059",x"36da",x"b02d",x"3bee",x"0000",x"3a8b",x"3b80",x"b544",x"4059",x"3710",x"b138",x"3be4",x"0000",x"3a96",x"3b84"),
(x"b575",x"4038",x"3710",x"bab5",x"b85c",x"8000",x"3a4c",x"3b4c",x"b575",x"4038",x"36da",x"bb97",x"b50d",x"0000",x"3a42",x"3b4c",x"b575",x"403a",x"3710",x"bb59",x"3650",x"8000",x"3a4c",x"3b4e"),
(x"b544",x"4059",x"3710",x"b138",x"3be4",x"0000",x"3a96",x"3b84",x"b544",x"4059",x"36da",x"b46b",x"3bb0",x"0000",x"3a8b",x"3b84",x"b52b",x"405a",x"3710",x"b472",x"3baf",x"0000",x"3a96",x"3b89"),
(x"b5ce",x"4043",x"3710",x"2ae9",x"bbfc",x"0000",x"3a4c",x"3b6a",x"b5ce",x"4043",x"36da",x"2f26",x"bbf3",x"0000",x"3a42",x"3b6a",x"b62a",x"4041",x"3710",x"303a",x"bbed",x"0000",x"3a4c",x"3b7c"),
(x"b52b",x"405a",x"3710",x"b472",x"3baf",x"0000",x"3a96",x"3b89",x"b52b",x"405a",x"36da",x"b237",x"3bd8",x"0000",x"3a8b",x"3b89",x"b50d",x"405b",x"3710",x"253f",x"3bff",x"0000",x"3a96",x"3b8f"),
(x"b5bd",x"4043",x"3710",x"b6e1",x"bb38",x"0000",x"3a4c",x"3b66",x"b5bd",x"4043",x"36da",x"b559",x"bb8a",x"0000",x"3a42",x"3b66",x"b5ce",x"4043",x"3710",x"2ae9",x"bbfc",x"0000",x"3a4c",x"3b6a"),
(x"b50d",x"405b",x"3710",x"253f",x"3bff",x"0000",x"3a96",x"3b8f",x"b50d",x"405b",x"36da",x"324a",x"3bd8",x"8000",x"3a8b",x"3b8f",x"b4f9",x"405a",x"3710",x"38a5",x"3a82",x"068d",x"3a96",x"3b93"),
(x"b5a1",x"4041",x"3710",x"b67b",x"bb50",x"8000",x"3a4c",x"3b60",x"b5a1",x"4041",x"36da",x"b72c",x"bb26",x"8000",x"3a42",x"3b60",x"b5bd",x"4043",x"3710",x"b6e1",x"bb38",x"0000",x"3a4c",x"3b66"),
(x"b4f9",x"405a",x"3710",x"38a5",x"3a82",x"068d",x"3a96",x"3b93",x"b4f9",x"405a",x"36da",x"3a57",x"38e0",x"8000",x"3a8b",x"3b93",x"b4f5",x"4058",x"3710",x"3bbb",x"341b",x"8000",x"3a96",x"3b96"),
(x"b581",x"403f",x"3710",x"b89f",x"ba87",x"0000",x"3a4c",x"3b59",x"b581",x"403f",x"36da",x"b794",x"bb0b",x"0000",x"3a42",x"3b59",x"b5a1",x"4041",x"3710",x"b67b",x"bb50",x"8000",x"3a4c",x"3b60"),
(x"b4f5",x"4058",x"3710",x"3bbb",x"341b",x"8000",x"3a96",x"3b96",x"b4f5",x"4058",x"36da",x"3bc4",x"33a2",x"0000",x"3a8b",x"3b96",x"b4f2",x"4056",x"3710",x"3aea",x"3805",x"8000",x"3a96",x"3b98"),
(x"b931",x"404d",x"3710",x"bbea",x"a7ae",x"307d",x"39d7",x"33c4",x"b931",x"404d",x"36da",x"bbff",x"a4d0",x"0000",x"39d6",x"33f3",x"b931",x"4059",x"3710",x"bbfe",x"a4d0",x"28c6",x"39ea",x"33c9"),
(x"b8ff",x"4059",x"3710",x"2581",x"3bff",x"15bc",x"3a23",x"3b9f",x"b8ff",x"4059",x"36da",x"26a7",x"3bff",x"8000",x"3a2d",x"3b9f",x"b8a3",x"4058",x"3710",x"286a",x"3bfe",x"8000",x"3a23",x"3b7b"),
(x"b568",x"403c",x"3710",x"bb03",x"b7b1",x"868d",x"3a4c",x"3b53",x"b568",x"403c",x"36da",x"b9f3",x"b958",x"0000",x"3a42",x"3b53",x"b581",x"403f",x"3710",x"b89f",x"ba87",x"0000",x"3a4c",x"3b59"),
(x"b4f2",x"4056",x"3710",x"3aea",x"3805",x"8000",x"3a96",x"3b98",x"b4f2",x"4056",x"36da",x"3a46",x"38f6",x"0000",x"3a8b",x"3b98",x"b4da",x"4053",x"3710",x"3a4b",x"38ef",x"0000",x"3a96",x"3b9f"),
(x"b8a3",x"4058",x"3710",x"286a",x"3bfe",x"8000",x"3a23",x"3b7b",x"b8a3",x"4058",x"36da",x"2a59",x"3bfd",x"0000",x"3a2d",x"3b7b",x"b89e",x"4058",x"3710",x"36f0",x"3b35",x"0000",x"3a23",x"3b79"),
(x"b558",x"4036",x"3710",x"b02d",x"bbee",x"0000",x"3a4c",x"3b44",x"b558",x"4036",x"36da",x"b3cc",x"bbc2",x"8000",x"3a42",x"3b44",x"b568",x"4037",x"3710",x"b810",x"bae4",x"0000",x"3a4c",x"3b48"),
(x"b4da",x"4053",x"3710",x"3a4b",x"38ef",x"0000",x"3a96",x"3b9f",x"b4da",x"4053",x"36da",x"3afc",x"37cc",x"0000",x"3a8b",x"3b9f",x"b4d8",x"4051",x"3710",x"3be5",x"b11d",x"868d",x"3a96",x"3ba1"),
(x"b89e",x"4058",x"3710",x"36f0",x"3b35",x"0000",x"3a23",x"3b79",x"b89e",x"4058",x"36da",x"380f",x"3ae4",x"068d",x"3a2d",x"3b79",x"b88f",x"4055",x"3710",x"380a",x"3ae7",x"0000",x"3a23",x"3b72"),
(x"b544",x"4036",x"3710",x"b46b",x"bbb0",x"0000",x"3a4c",x"3b40",x"b544",x"4036",x"36da",x"b138",x"bbe4",x"0000",x"3a42",x"3b40",x"b558",x"4036",x"3710",x"b02d",x"bbee",x"0000",x"3a4c",x"3b44"),
(x"b4d8",x"4051",x"3710",x"3be5",x"b11d",x"868d",x"3a96",x"3ba1",x"b4d8",x"4051",x"36da",x"3af9",x"b7d8",x"8000",x"3a8b",x"3ba1",x"b4e1",x"4050",x"3710",x"3599",x"bb7e",x"0000",x"3a96",x"3ba3"),
(x"b88f",x"4055",x"3710",x"380a",x"3ae7",x"0000",x"3a23",x"3b72",x"b88f",x"4055",x"36da",x"377a",x"3b12",x"0000",x"3a2d",x"3b72",x"b87d",x"4053",x"3710",x"3541",x"3b8e",x"0000",x"3a23",x"3b6a"),
(x"b52b",x"4035",x"3710",x"b237",x"bbd8",x"0000",x"3a4c",x"3b3b",x"b52b",x"4035",x"36da",x"b472",x"bbaf",x"0000",x"3a42",x"3b3b",x"b544",x"4036",x"3710",x"b46b",x"bbb0",x"0000",x"3a4c",x"3b40"),
(x"b4e1",x"4050",x"3710",x"3599",x"bb7e",x"0000",x"3a96",x"3ba3",x"b4e1",x"4050",x"36da",x"33d2",x"bbc1",x"8000",x"3a8b",x"3ba3",x"b51a",x"404f",x"3710",x"332b",x"bbcb",x"0000",x"3a96",x"3bae"),
(x"b87d",x"4053",x"3710",x"3541",x"3b8e",x"0000",x"3a23",x"3b6a",x"b87d",x"4053",x"36da",x"3244",x"3bd8",x"0000",x"3a2d",x"3b6a",x"b86e",x"4053",x"3710",x"ad02",x"3bf9",x"0000",x"3a23",x"3b64"),
(x"b50d",x"4034",x"3710",x"324a",x"bbd8",x"8000",x"3a4c",x"3b35",x"b50d",x"4034",x"36da",x"253f",x"bbff",x"8000",x"3a42",x"3b35",x"b52b",x"4035",x"3710",x"b237",x"bbd8",x"0000",x"3a4c",x"3b3b"),
(x"b51a",x"404f",x"3710",x"332b",x"bbcb",x"0000",x"3a96",x"3bae",x"b51a",x"404f",x"36da",x"347c",x"bbad",x"0000",x"3a8b",x"3bae",x"b528",x"404e",x"3710",x"37ff",x"baed",x"0000",x"3a96",x"3bb1"),
(x"b86e",x"4053",x"3710",x"ad02",x"3bf9",x"0000",x"3a23",x"3b64",x"b86e",x"4053",x"36da",x"b407",x"3bbe",x"8000",x"3a2d",x"3b64",x"b867",x"4054",x"3710",x"b975",x"39d8",x"0000",x"3a23",x"3b61"),
(x"b4f9",x"4035",x"3710",x"3a57",x"b8e0",x"0000",x"3a4c",x"3b31",x"b4f9",x"4035",x"36da",x"38a5",x"ba82",x"8000",x"3a42",x"3b31",x"b50d",x"4034",x"3710",x"324a",x"bbd8",x"8000",x"3a4c",x"3b35"),
(x"b528",x"404e",x"3710",x"37ff",x"baed",x"0000",x"3a96",x"3bb1",x"b528",x"404e",x"36da",x"38ed",x"ba4d",x"8000",x"3a8b",x"3bb1",x"b52c",x"404e",x"3710",x"3bfc",x"ab69",x"0000",x"3a96",x"3bb2"),
(x"b867",x"4054",x"3710",x"b975",x"39d8",x"0000",x"3a23",x"3b61",x"b867",x"4054",x"36da",x"baa2",x"3877",x"0000",x"3a2d",x"3b61",x"b865",x"4055",x"3710",x"bb0e",x"378a",x"0000",x"3a23",x"3b5e"),
(x"b4f5",x"4037",x"3710",x"3bc4",x"b3a1",x"8000",x"3a4c",x"3b2e",x"b4f5",x"4037",x"36da",x"3bbb",x"b41b",x"8000",x"3a42",x"3b2e",x"b4f9",x"4035",x"3710",x"3a57",x"b8e0",x"0000",x"3a4c",x"3b31"),
(x"b52c",x"404e",x"3710",x"3bfc",x"ab69",x"0000",x"3b1c",x"39ae",x"b52c",x"404e",x"36da",x"3b0d",x"378c",x"0000",x"3b11",x"39ae",x"b526",x"404d",x"3710",x"35f8",x"3b6b",x"0000",x"3b1c",x"39af"),
(x"b865",x"4055",x"3710",x"bb0e",x"378a",x"0000",x"3a23",x"3b5e",x"b865",x"4055",x"36da",x"baaf",x"3865",x"8000",x"3a2d",x"3b5e",x"b85e",x"4058",x"3710",x"b878",x"3aa2",x"0000",x"3a23",x"3b5a"),
(x"b4f2",x"4038",x"3710",x"3a46",x"b8f6",x"0000",x"3a4c",x"3b2b",x"b4f2",x"4038",x"36da",x"3aea",x"b805",x"8000",x"3a42",x"3b2b",x"b4f5",x"4037",x"3710",x"3bc4",x"b3a1",x"8000",x"3a4c",x"3b2e"),
(x"b526",x"404d",x"3710",x"35f8",x"3b6b",x"0000",x"3b1c",x"39af",x"b526",x"404d",x"36da",x"33bb",x"3bc3",x"0000",x"3b11",x"39af",x"b50c",x"404c",x"3710",x"292b",x"3bfe",x"8000",x"3b1c",x"39b4"),
(x"b116",x"404a",x"3710",x"3b51",x"3675",x"0000",x"3a5a",x"3b6f",x"b116",x"404a",x"36da",x"3bdf",x"31b0",x"868d",x"3a50",x"3b6f",x"b116",x"4045",x"3710",x"3bdf",x"b1b0",x"0000",x"3a5a",x"3b75"),
(x"b85e",x"4058",x"3710",x"b878",x"3aa2",x"0000",x"3a23",x"3b5a",x"b85e",x"4058",x"36da",x"b5f3",x"3b6d",x"8000",x"3a2d",x"3b5a",x"b84a",x"4059",x"3710",x"ac15",x"3bfb",x"868d",x"3a23",x"3b51"),
(x"b4da",x"403c",x"3710",x"3afc",x"b7cc",x"8000",x"3a4c",x"3b24",x"b4da",x"403c",x"36da",x"3a4b",x"b8ef",x"068d",x"3a42",x"3b24",x"b4f2",x"4038",x"3710",x"3a46",x"b8f6",x"0000",x"3a4c",x"3b2b"),
(x"b451",x"404c",x"3710",x"a0dd",x"3c00",x"0000",x"3b1c",x"39d8",x"b451",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3b11",x"39d8",x"b441",x"404d",x"3710",x"b6f3",x"3b34",x"0000",x"3b1c",x"39db"),
(x"b89e",x"4037",x"3710",x"380f",x"bae4",x"068d",x"3a07",x"3b76",x"b89e",x"4037",x"36da",x"36f0",x"bb35",x"0000",x"39fd",x"3b76",x"b8a3",x"4037",x"3710",x"2a1e",x"bbfd",x"0000",x"3a07",x"3b78"),
(x"b84a",x"4059",x"3710",x"ac15",x"3bfb",x"868d",x"3a23",x"3b51",x"b84a",x"4059",x"36da",x"30e0",x"3be8",x"8000",x"3a2d",x"3b51",x"b83a",x"4057",x"3710",x"3890",x"3a92",x"0000",x"3a23",x"3b4b"),
(x"b4d8",x"403d",x"3710",x"3af9",x"37d7",x"868d",x"3a4c",x"3b22",x"b4d8",x"403d",x"36da",x"3be5",x"311d",x"0000",x"3a42",x"3b22",x"b4da",x"403c",x"3710",x"3afc",x"b7cc",x"8000",x"3a4c",x"3b24"),
(x"b50c",x"404c",x"3710",x"292b",x"3bfe",x"8000",x"3b1c",x"39b4",x"b50c",x"404c",x"36da",x"236c",x"3bff",x"0000",x"3b11",x"39b4",x"b451",x"404c",x"3710",x"a0dd",x"3c00",x"0000",x"3b1c",x"39d8"),
(x"b88f",x"403a",x"3710",x"377a",x"bb12",x"8000",x"3a07",x"3b6f",x"b88f",x"403a",x"36da",x"380a",x"bae7",x"0000",x"39fd",x"3b6f",x"b89e",x"4037",x"3710",x"380f",x"bae4",x"068d",x"3a07",x"3b76"),
(x"b568",x"4053",x"3710",x"b9f3",x"3958",x"0000",x"3a96",x"3b72",x"b568",x"4053",x"36da",x"bb03",x"37b2",x"868d",x"3a8b",x"3b72",x"b569",x"4054",x"3710",x"bb2d",x"b70f",x"0000",x"3a96",x"3b74"),
(x"b4e1",x"403e",x"3710",x"33d2",x"3bc1",x"868d",x"3a4c",x"3b1f",x"b4e1",x"403e",x"36da",x"3599",x"3b7e",x"0000",x"3a42",x"3b1f",x"b4d8",x"403d",x"3710",x"3af9",x"37d7",x"868d",x"3a4c",x"3b22"),
(x"b441",x"404d",x"3710",x"b6f3",x"3b34",x"0000",x"3b1c",x"39db",x"b441",x"404d",x"36da",x"b7a3",x"3b07",x"0000",x"3b11",x"39db",x"b40d",x"4051",x"3710",x"b83a",x"3aca",x"0000",x"3b1c",x"39e6"),
(x"b87d",x"403c",x"3710",x"3244",x"bbd8",x"0000",x"3a07",x"3b67",x"b87d",x"403c",x"36da",x"3541",x"bb8e",x"0000",x"39fd",x"3b67",x"b88f",x"403a",x"3710",x"377a",x"bb12",x"8000",x"3a07",x"3b6f"),
(x"b83a",x"4057",x"3710",x"3890",x"3a92",x"0000",x"3a23",x"3b4b",x"b83a",x"4057",x"36da",x"3953",x"39f7",x"8000",x"3a2d",x"3b4b",x"b820",x"4051",x"3710",x"391f",x"3a25",x"0000",x"3a23",x"3b3c"),
(x"b51a",x"4040",x"3710",x"347c",x"3bad",x"8000",x"3a4c",x"3b14",x"b51a",x"4040",x"36da",x"332b",x"3bcb",x"0000",x"3a42",x"3b14",x"b4e1",x"403e",x"3710",x"33d2",x"3bc1",x"868d",x"3a4c",x"3b1f"),
(x"b40d",x"4051",x"3710",x"b83a",x"3aca",x"0000",x"3b1c",x"39e6",x"b40d",x"4051",x"36da",x"b8bf",x"3a70",x"068d",x"3b11",x"39e6",x"b407",x"4052",x"3710",x"bb61",x"362a",x"0000",x"3b1c",x"39e8"),
(x"b86e",x"403c",x"3710",x"b406",x"bbbe",x"0000",x"3a07",x"3b61",x"b86e",x"403c",x"36da",x"ad01",x"bbf9",x"0000",x"39fd",x"3b61",x"b87d",x"403c",x"3710",x"3244",x"bbd8",x"0000",x"3a07",x"3b67"),
(x"b569",x"4054",x"3710",x"bb2d",x"b70f",x"0000",x"3a96",x"3b74",x"b569",x"4054",x"36da",x"ba4b",x"b8f0",x"0000",x"3a8b",x"3b74",x"b575",x"4055",x"3710",x"ba67",x"b8cb",x"0000",x"3a96",x"3b77"),
(x"b528",x"4041",x"3710",x"38ed",x"3a4d",x"8000",x"3a4c",x"3b11",x"b528",x"4041",x"36da",x"37fe",x"3aed",x"0000",x"3a42",x"3b11",x"b51a",x"4040",x"3710",x"347c",x"3bad",x"8000",x"3a4c",x"3b14"),
(x"b407",x"4052",x"3710",x"bb61",x"362a",x"0000",x"3b1c",x"39e8",x"b407",x"4052",x"36da",x"bbf7",x"2ddc",x"0000",x"3b11",x"39e8",x"b409",x"4053",x"3710",x"bb1a",x"b75c",x"8000",x"3b1c",x"39e9"),
(x"b867",x"403b",x"3710",x"baa2",x"b877",x"0000",x"3a07",x"3b5e",x"b867",x"403b",x"36da",x"b975",x"b9d8",x"0000",x"39fd",x"3b5e",x"b86e",x"403c",x"3710",x"b406",x"bbbe",x"0000",x"3a07",x"3b61"),
(x"b820",x"4051",x"3710",x"391f",x"3a25",x"0000",x"3a23",x"3b3c",x"b820",x"4051",x"36da",x"385c",x"3ab4",x"0000",x"3a2d",x"3b3c",x"b801",x"404d",x"3710",x"3561",x"3b88",x"0000",x"3a23",x"3b2e"),
(x"b52c",x"4041",x"3710",x"3b0d",x"b78c",x"0000",x"3a4c",x"3b10",x"b52c",x"4041",x"36da",x"3bfc",x"2b6f",x"0000",x"3a42",x"3b10",x"b528",x"4041",x"3710",x"38ed",x"3a4d",x"8000",x"3a4c",x"3b11"),
(x"b409",x"4053",x"3710",x"bb1a",x"b75c",x"8000",x"3b1c",x"39e9",x"b409",x"4053",x"36da",x"bab5",x"b85b",x"0000",x"3b11",x"39e9",x"b413",x"4054",x"3710",x"bb08",x"b7a1",x"868d",x"3b1c",x"39ed"),
(x"b865",x"4039",x"3710",x"baaf",x"b865",x"8000",x"3a07",x"3b5b",x"b865",x"4039",x"36da",x"bb0e",x"b78a",x"0000",x"39fd",x"3b5b",x"b867",x"403b",x"3710",x"baa2",x"b877",x"0000",x"3a07",x"3b5e"),
(x"b801",x"404d",x"3710",x"3561",x"3b88",x"0000",x"3a23",x"3b2e",x"b801",x"404d",x"36da",x"3346",x"3bca",x"0000",x"3a2d",x"3b2e",x"b7c0",x"404c",x"3710",x"29e3",x"3bfd",x"0000",x"3a23",x"3b21"),
(x"b526",x"4042",x"3710",x"33bc",x"bbc3",x"0000",x"3afb",x"3a0f",x"b526",x"4042",x"36da",x"35f9",x"bb6b",x"0000",x"3af0",x"3a0f",x"b52c",x"4041",x"3710",x"3b0d",x"b78c",x"0000",x"3afb",x"3a11"),
(x"b413",x"4054",x"3710",x"bb08",x"b7a1",x"868d",x"3b1c",x"39ed",x"b413",x"4054",x"36da",x"bba9",x"b499",x"0000",x"3b11",x"39ed",x"b413",x"4055",x"3710",x"bb8c",x"354a",x"868d",x"3b1c",x"39ee"),
(x"b85e",x"4037",x"3710",x"b5f3",x"bb6d",x"8000",x"3a07",x"3b57",x"b85e",x"4037",x"36da",x"b878",x"baa2",x"0000",x"39fd",x"3b57",x"b865",x"4039",x"3710",x"baaf",x"b865",x"8000",x"3a07",x"3b5b"),
(x"b7c0",x"404c",x"3710",x"29e3",x"3bfd",x"0000",x"3a23",x"3b21",x"b7c0",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3a2d",x"3b21",x"b794",x"404d",x"3710",x"b357",x"3bc9",x"0000",x"3a23",x"3b18"),
(x"b50c",x"4042",x"3710",x"236c",x"bbff",x"0000",x"3afb",x"3a0a",x"b50c",x"4042",x"36da",x"292b",x"bbfe",x"8000",x"3af0",x"3a0a",x"b526",x"4042",x"3710",x"33bc",x"bbc3",x"0000",x"3afb",x"3a0f"),
(x"b413",x"4055",x"3710",x"bb8c",x"354a",x"868d",x"3b1c",x"39ee",x"b413",x"4055",x"36da",x"ba12",x"3935",x"8000",x"3b11",x"39ee",x"b40b",x"4056",x"3710",x"b3aa",x"3bc4",x"8000",x"3b1c",x"39f0"),
(x"b84a",x"4036",x"3710",x"30e0",x"bbe8",x"8000",x"3a07",x"3b4e",x"b84a",x"4036",x"36da",x"ac15",x"bbfb",x"068d",x"39fd",x"3b4e",x"b85e",x"4037",x"3710",x"b5f3",x"bb6d",x"8000",x"3a07",x"3b57"),
(x"b794",x"404d",x"3710",x"b357",x"3bc9",x"0000",x"3a23",x"3b18",x"b794",x"404d",x"36da",x"b51c",x"3b94",x"0000",x"3a2d",x"3b18",x"b77a",x"404e",x"3710",x"b83f",x"3ac7",x"0000",x"3a23",x"3b13"),
(x"b441",x"4042",x"3710",x"b7a4",x"bb07",x"0000",x"3afb",x"39e4",x"b441",x"4042",x"36da",x"b6f3",x"bb34",x"0000",x"3af0",x"39e4",x"b451",x"4042",x"3710",x"a987",x"bbfe",x"8000",x"3afb",x"39e7"),
(x"b40b",x"4056",x"3710",x"b3aa",x"3bc4",x"8000",x"3b1c",x"39f0",x"b40b",x"4056",x"36da",x"aabe",x"3bfd",x"868d",x"3b11",x"39f0",x"b3f4",x"4056",x"3710",x"3148",x"3be3",x"8000",x"3b1c",x"39f3"),
(x"b83a",x"4037",x"3710",x"3953",x"b9f7",x"068d",x"3a07",x"3b48",x"b83a",x"4037",x"36da",x"3890",x"ba92",x"0000",x"39fd",x"3b48",x"b84a",x"4036",x"3710",x"30e0",x"bbe8",x"8000",x"3a07",x"3b4e"),
(x"b77a",x"404e",x"3710",x"b83f",x"3ac7",x"0000",x"3a23",x"3b13",x"b77a",x"404e",x"36da",x"b97c",x"39d2",x"0000",x"3a2d",x"3b13",x"b776",x"4050",x"3710",x"bbee",x"3037",x"0000",x"3a23",x"3b10"),
(x"b451",x"4042",x"3710",x"a987",x"bbfe",x"8000",x"3afb",x"39e7",x"b451",x"4042",x"36da",x"a0ea",x"bc00",x"0000",x"3af0",x"39e7",x"b50c",x"4042",x"3710",x"236c",x"bbff",x"0000",x"3afb",x"3a0a"),
(x"b3f4",x"4056",x"3710",x"3148",x"3be3",x"8000",x"3b1c",x"39f3",x"b3f4",x"4056",x"36da",x"3408",x"3bbd",x"0000",x"3b11",x"39f3",x"b3d2",x"4055",x"3710",x"2ffb",x"3bf0",x"0000",x"3b1c",x"39f7"),
(x"b569",x"403b",x"3710",x"ba4b",x"38f0",x"0000",x"3a4c",x"3b51",x"b569",x"403b",x"36da",x"bb2d",x"370f",x"0000",x"3a42",x"3b51",x"b568",x"403c",x"3710",x"bb03",x"b7b1",x"868d",x"3a4c",x"3b53"),
(x"b776",x"4050",x"3710",x"bbee",x"3037",x"0000",x"3a23",x"3b10",x"b776",x"4050",x"36da",x"bbce",x"b2fb",x"0000",x"3a2d",x"3b10",x"b77b",x"4051",x"3710",x"b937",x"ba10",x"0000",x"3a23",x"3b0f"),
(x"b40d",x"403e",x"3710",x"b8bf",x"ba70",x"8000",x"3afb",x"39d8",x"b40d",x"403e",x"36da",x"b83a",x"baca",x"0000",x"3af0",x"39d8",x"b441",x"4042",x"3710",x"b7a4",x"bb07",x"0000",x"3afb",x"39e4"),
(x"b3d2",x"4055",x"3710",x"2ffb",x"3bf0",x"0000",x"3b1c",x"39f7",x"b3d2",x"4055",x"36da",x"abf9",x"3bfc",x"0000",x"3b11",x"39f7",x"b3a5",x"4056",x"3710",x"24fd",x"3bff",x"0000",x"3b1c",x"39fb"),
(x"b820",x"403e",x"3710",x"385c",x"bab4",x"8000",x"3a07",x"3b39",x"b820",x"403e",x"36da",x"391f",x"ba25",x"0000",x"39fd",x"3b39",x"b83a",x"4037",x"3710",x"3953",x"b9f7",x"068d",x"3a07",x"3b48"),
(x"b77b",x"4051",x"3710",x"b937",x"ba10",x"0000",x"3a93",x"3ac5",x"b77b",x"4051",x"36da",x"b853",x"baba",x"0000",x"3a88",x"3ac5",x"b790",x"4052",x"3710",x"b606",x"bb69",x"0000",x"3a93",x"3ac9"),
(x"b407",x"403d",x"3710",x"bbf7",x"addb",x"0000",x"3afb",x"39d6",x"b407",x"403d",x"36da",x"bb61",x"b629",x"0000",x"3af0",x"39d6",x"b40d",x"403e",x"3710",x"b8bf",x"ba70",x"8000",x"3afb",x"39d8"),
(x"b3a5",x"4056",x"3710",x"24fd",x"3bff",x"0000",x"3b1c",x"39fb",x"b3a5",x"4056",x"36da",x"32b6",x"3bd2",x"068d",x"3b11",x"39fb",x"b368",x"4054",x"3710",x"37ea",x"3af3",x"8000",x"3b1c",x"3a01"),
(x"b575",x"403a",x"3710",x"bb59",x"3650",x"8000",x"3a4c",x"3b4e",x"b575",x"403a",x"36da",x"ba67",x"38cb",x"868d",x"3a42",x"3b4e",x"b569",x"403b",x"3710",x"ba4b",x"38f0",x"0000",x"3a4c",x"3b51"),
(x"b790",x"4052",x"3710",x"b606",x"bb69",x"0000",x"3a93",x"3ac9",x"b790",x"4052",x"36da",x"b461",x"bbb1",x"0000",x"3a88",x"3ac9",x"b7a8",x"4053",x"3710",x"b360",x"bbc8",x"0000",x"3a93",x"3ace"),
(x"b409",x"403c",x"3710",x"bab5",x"385b",x"0000",x"3afb",x"39d5",x"b409",x"403c",x"36da",x"bb1a",x"375d",x"0000",x"3af0",x"39d5",x"b407",x"403d",x"3710",x"bbf7",x"addb",x"0000",x"3afb",x"39d6"),
(x"b368",x"4054",x"3710",x"37ea",x"3af3",x"8000",x"3b1c",x"3a01",x"b368",x"4054",x"36da",x"3912",x"3a2f",x"8000",x"3b11",x"3a01",x"b340",x"4051",x"3710",x"3aba",x"3853",x"0000",x"3b1c",x"3a07"),
(x"b801",x"4042",x"3710",x"3346",x"bbca",x"0000",x"3a07",x"3b2b",x"b801",x"4042",x"36da",x"3561",x"bb88",x"0000",x"39fd",x"3b2b",x"b820",x"403e",x"3710",x"385c",x"bab4",x"8000",x"3a07",x"3b39"),
(x"b7a8",x"4053",x"3710",x"b360",x"bbc8",x"0000",x"3a93",x"3ace",x"b7a8",x"4053",x"36da",x"b4b8",x"bba4",x"8000",x"3a88",x"3ace",x"b7bd",x"4054",x"3710",x"b6d2",x"bb3c",x"0000",x"3a93",x"3ad2"),
(x"b413",x"403a",x"3710",x"bba9",x"3499",x"8000",x"3afb",x"39d2",x"b413",x"403a",x"36da",x"bb07",x"37a1",x"8000",x"3af0",x"39d2",x"b409",x"403c",x"3710",x"bab5",x"385b",x"0000",x"3afb",x"39d5"),
(x"b340",x"4051",x"3710",x"3aba",x"3853",x"0000",x"3b1c",x"3a07",x"b340",x"4051",x"36da",x"3b6b",x"35fb",x"8000",x"3b11",x"3a07",x"b33a",x"404f",x"3710",x"3bf6",x"ae02",x"8000",x"3b1c",x"3a0b"),
(x"b7c0",x"4043",x"3710",x"a984",x"bbfe",x"0000",x"3a07",x"3b1e",x"b7c0",x"4043",x"36da",x"29e3",x"bbfd",x"0000",x"39fd",x"3b1e",x"b801",x"4042",x"3710",x"3346",x"bbca",x"0000",x"3a07",x"3b2b"),
(x"b7bd",x"4054",x"3710",x"b6d2",x"bb3c",x"0000",x"3a93",x"3ad2",x"b7bd",x"4054",x"36da",x"b821",x"bada",x"8000",x"3a88",x"3ad2",x"b7c7",x"4055",x"3710",x"ba01",x"b948",x"0000",x"3a93",x"3ad5"),
(x"b931",x"4036",x"3710",x"bbe9",x"26a1",x"309e",x"39b2",x"33ca",x"b931",x"4036",x"36da",x"bbff",x"26b5",x"0000",x"39b3",x"33fa",x"b930",x"4041",x"3710",x"bbeb",x"2604",x"3075",x"39c5",x"33c0"),
(x"b413",x"4039",x"3710",x"ba12",x"b935",x"068d",x"3afb",x"39d0",x"b413",x"4039",x"36da",x"bb8c",x"b54a",x"868d",x"3af0",x"39d0",x"b413",x"403a",x"3710",x"bba9",x"3499",x"8000",x"3afb",x"39d2"),
(x"b33a",x"404f",x"3710",x"3bf6",x"ae02",x"8000",x"3b1c",x"3a0b",x"b33a",x"404f",x"36da",x"3b88",x"b564",x"068d",x"3b11",x"3a0b",x"b351",x"404d",x"3710",x"3b23",x"b738",x"0000",x"3b1c",x"3a0f"),
(x"b794",x"4042",x"3710",x"b51c",x"bb94",x"0000",x"3a07",x"3b15",x"b794",x"4042",x"36da",x"b357",x"bbc9",x"0000",x"39fd",x"3b15",x"b7c0",x"4043",x"3710",x"a984",x"bbfe",x"0000",x"3a07",x"3b1e"),
(x"b7c7",x"4055",x"3710",x"ba01",x"b948",x"0000",x"3a93",x"3ad5",x"b7c7",x"4055",x"36da",x"bb43",x"b6b4",x"0000",x"3a88",x"3ad5",x"b7c7",x"4055",x"3710",x"b8b7",x"3a76",x"0000",x"3a93",x"3ad6"),
(x"b40b",x"4039",x"3710",x"aabe",x"bbfd",x"8000",x"3afb",x"39ce",x"b40b",x"4039",x"36da",x"b3aa",x"bbc4",x"0000",x"3af0",x"39ce",x"b413",x"4039",x"3710",x"ba12",x"b935",x"068d",x"3afb",x"39d0"),
(x"b351",x"404d",x"3710",x"3b23",x"b738",x"0000",x"3b1c",x"3a0f",x"b351",x"404d",x"36da",x"3bb2",x"b458",x"0000",x"3b11",x"3a0f",x"b34f",x"404c",x"3710",x"3913",x"3a2e",x"8000",x"3b1c",x"3a11"),
(x"b77a",x"4040",x"3710",x"b97c",x"b9d2",x"8000",x"3a07",x"3b10",x"b77a",x"4040",x"36da",x"b83f",x"bac7",x"0000",x"39fd",x"3b10",x"b794",x"4042",x"3710",x"b51c",x"bb94",x"0000",x"3a07",x"3b15"),
(x"b7c7",x"4055",x"3710",x"b8b7",x"3a76",x"0000",x"3a93",x"3ad6",x"b7c7",x"4055",x"36da",x"b744",x"3b20",x"0cea",x"3a88",x"3ad6",x"b7a4",x"4057",x"3710",x"b654",x"3b58",x"0000",x"3a93",x"3add"),
(x"b3f4",x"4039",x"3710",x"3408",x"bbbd",x"0000",x"3afb",x"39cb",x"b3f4",x"4039",x"36da",x"3148",x"bbe3",x"0000",x"3af0",x"39cb",x"b40b",x"4039",x"3710",x"aabe",x"bbfd",x"8000",x"3afb",x"39ce"),
(x"b34f",x"404c",x"3710",x"3913",x"3a2e",x"8000",x"3a5a",x"3b34",x"b34f",x"404c",x"36da",x"3448",x"3bb5",x"0000",x"3a50",x"3b34",x"b326",x"404b",x"3710",x"a5e9",x"3bff",x"0000",x"3a5a",x"3b38"),
(x"b776",x"403f",x"3710",x"bbce",x"32fb",x"0000",x"3b18",x"38ac",x"b776",x"403f",x"36da",x"bbee",x"b037",x"0000",x"3b18",x"38a2",x"b77a",x"4040",x"3710",x"b97c",x"b9d2",x"8000",x"3b16",x"38ac"),
(x"b7a4",x"4057",x"3710",x"b654",x"3b58",x"0000",x"3a93",x"3add",x"b7a4",x"4057",x"36da",x"b64b",x"3b5a",x"8000",x"3a88",x"3add",x"b783",x"4059",x"3710",x"b33d",x"3bca",x"0000",x"3a93",x"3ae4"),
(x"b3d2",x"403a",x"3710",x"abf9",x"bbfc",x"8000",x"3afb",x"39c8",x"b3d2",x"403a",x"36da",x"2ffb",x"bbf0",x"0000",x"3af0",x"39c8",x"b3f4",x"4039",x"3710",x"3408",x"bbbd",x"0000",x"3afb",x"39cb"),
(x"b326",x"404b",x"3710",x"a5e9",x"3bff",x"0000",x"3a5a",x"3b38",x"b326",x"404b",x"36da",x"ad8e",x"3bf8",x"0000",x"3a50",x"3b38",x"b2d6",x"404c",x"3710",x"b287",x"3bd4",x"0000",x"3a5a",x"3b3f"),
(x"b77b",x"403e",x"3710",x"b853",x"3aba",x"0000",x"3b1a",x"38ac",x"b77b",x"403e",x"36da",x"b937",x"3a10",x"8000",x"3b1a",x"38a2",x"b776",x"403f",x"3710",x"bbce",x"32fb",x"0000",x"3b18",x"38ac"),
(x"b783",x"4059",x"3710",x"b33d",x"3bca",x"0000",x"3a93",x"3ae4",x"b783",x"4059",x"36da",x"afa0",x"3bf1",x"0000",x"3a88",x"3ae4",x"b73e",x"4059",x"3710",x"27ae",x"3bfe",x"0000",x"3a93",x"3af1"),
(x"b3a5",x"4039",x"3710",x"32b6",x"bbd2",x"0000",x"3afb",x"39c3",x"b3a5",x"4039",x"36da",x"2504",x"bbff",x"0000",x"3af0",x"39c3",x"b3d2",x"403a",x"3710",x"abf9",x"bbfc",x"8000",x"3afb",x"39c8"),
(x"b2d6",x"404c",x"3710",x"b287",x"3bd4",x"0000",x"3a5a",x"3b3f",x"b2d6",x"404c",x"36da",x"b4dd",x"3b9f",x"0000",x"3a50",x"3b3f",x"b2aa",x"404d",x"3710",x"b78b",x"3b0e",x"0000",x"3a5a",x"3b44"),
(x"b790",x"403d",x"3710",x"b461",x"3bb1",x"0000",x"3b1e",x"38ac",x"b790",x"403d",x"36da",x"b606",x"3b69",x"0000",x"3b1e",x"38a2",x"b77b",x"403e",x"3710",x"b853",x"3aba",x"0000",x"3b1a",x"38ac"),
(x"b73e",x"4059",x"3710",x"27ae",x"3bfe",x"0000",x"3a93",x"3af1",x"b73e",x"4059",x"36da",x"2f57",x"3bf2",x"8000",x"3a88",x"3af1",x"b705",x"4058",x"3710",x"34b8",x"3ba4",x"0000",x"3a93",x"3afc"),
(x"b368",x"403a",x"3710",x"3912",x"ba2f",x"0000",x"3afb",x"39bd",x"b368",x"403a",x"36da",x"37ea",x"baf3",x"8000",x"3af0",x"39bd",x"b3a5",x"4039",x"3710",x"32b6",x"bbd2",x"0000",x"3afb",x"39c3"),
(x"b2aa",x"404d",x"3710",x"b78b",x"3b0e",x"0000",x"3a5a",x"3b44",x"b2aa",x"404d",x"36da",x"b7e2",x"3af5",x"0000",x"3a50",x"3b44",x"b261",x"4050",x"3710",x"b72e",x"3b26",x"8000",x"3a5a",x"3b4c"),
(x"b7a8",x"403c",x"3710",x"b4b8",x"3ba4",x"8000",x"3a7c",x"3b0f",x"b7a8",x"403c",x"36da",x"b360",x"3bc8",x"8000",x"3a72",x"3b0f",x"b790",x"403d",x"3710",x"b461",x"3bb1",x"0000",x"3a7c",x"3b13"),
(x"b705",x"4058",x"3710",x"34b8",x"3ba4",x"0000",x"3a93",x"3afc",x"b705",x"4058",x"36da",x"36ee",x"3b35",x"0000",x"3a88",x"3afc",x"b6f1",x"4056",x"3710",x"3a69",x"38c9",x"068d",x"3a93",x"3b01"),
(x"b340",x"403d",x"3710",x"3b6b",x"b5fb",x"0000",x"3afb",x"39b7",x"b340",x"403d",x"36da",x"3aba",x"b853",x"8000",x"3af0",x"39b7",x"b368",x"403a",x"3710",x"3912",x"ba2f",x"0000",x"3afb",x"39bd"),
(x"b261",x"4050",x"3710",x"b72e",x"3b26",x"8000",x"3a5a",x"3b4c",x"b261",x"4050",x"36da",x"b5e0",x"3b70",x"8000",x"3a50",x"3b4c",x"b22d",x"4051",x"3710",x"ae8a",x"3bf5",x"8000",x"3a5a",x"3b51"),
(x"b7bd",x"403b",x"3710",x"b821",x"3ada",x"8000",x"3a7c",x"3b0b",x"b7bd",x"403b",x"36da",x"b6d2",x"3b3c",x"0000",x"3a72",x"3b0b",x"b7a8",x"403c",x"3710",x"b4b8",x"3ba4",x"8000",x"3a7c",x"3b0f"),
(x"b6f1",x"4056",x"3710",x"3a69",x"38c9",x"068d",x"3a93",x"3b01",x"b6f1",x"4056",x"36da",x"3b73",x"35d3",x"8000",x"3a88",x"3b01",x"b6ef",x"4053",x"3710",x"3be9",x"b0b7",x"0000",x"3a93",x"3b05"),
(x"b33a",x"4040",x"3710",x"3b88",x"3564",x"0000",x"3afb",x"39b3",x"b33a",x"4040",x"36da",x"3bf6",x"2e02",x"8000",x"3af0",x"39b3",x"b340",x"403d",x"3710",x"3b6b",x"b5fb",x"0000",x"3afb",x"39b7"),
(x"b22d",x"4051",x"3710",x"ae8a",x"3bf5",x"8000",x"3a5a",x"3b51",x"b22d",x"4051",x"36da",x"2c28",x"3bfb",x"0000",x"3a50",x"3b51",x"b1fd",x"4050",x"3710",x"35da",x"3b72",x"0000",x"3a5a",x"3b56"),
(x"b7c7",x"403a",x"3710",x"bb43",x"36b4",x"0000",x"3a7c",x"3b08",x"b7c7",x"403a",x"36da",x"ba01",x"3948",x"8000",x"3a72",x"3b08",x"b7bd",x"403b",x"3710",x"b821",x"3ada",x"8000",x"3a7c",x"3b0b"),
(x"b6ef",x"4053",x"3710",x"3be9",x"b0b7",x"0000",x"3a93",x"3b05",x"b6ef",x"4053",x"36da",x"3b57",x"b659",x"8000",x"3a88",x"3b05",x"b6fb",x"4051",x"3710",x"38e1",x"ba57",x"0000",x"3a93",x"3b08"),
(x"b351",x"4042",x"3710",x"3bb3",x"3458",x"0000",x"3afb",x"39af",x"b351",x"4042",x"36da",x"3b23",x"3738",x"0000",x"3af0",x"39af",x"b33a",x"4040",x"3710",x"3b88",x"3564",x"0000",x"3afb",x"39b3"),
(x"b1fd",x"4050",x"3710",x"35da",x"3b72",x"0000",x"3a5a",x"3b56",x"b1fd",x"4050",x"36da",x"375d",x"3b1a",x"8000",x"3a50",x"3b56",x"b1c1",x"404e",x"3710",x"37bd",x"3b00",x"0000",x"3a5a",x"3b5d"),
(x"b7c7",x"4039",x"3710",x"b744",x"bb20",x"868d",x"3a7c",x"3b07",x"b7c7",x"4039",x"36da",x"b8b7",x"ba76",x"0000",x"3a72",x"3b07",x"b7c7",x"403a",x"3710",x"bb43",x"36b4",x"0000",x"3a7c",x"3b08"),
(x"b6fb",x"4051",x"3710",x"38e1",x"ba57",x"0000",x"3a93",x"3b08",x"b6fb",x"4051",x"36da",x"37ed",x"baf2",x"068d",x"3a88",x"3b08",x"b721",x"404f",x"3710",x"3711",x"bb2d",x"0000",x"3a93",x"3b10"),
(x"b34f",x"4043",x"3710",x"3448",x"bbb5",x"0000",x"3afb",x"39ae",x"b34f",x"4043",x"36da",x"3913",x"ba2f",x"8000",x"3af0",x"39ae",x"b351",x"4042",x"3710",x"3bb3",x"3458",x"0000",x"3afb",x"39af"),
(x"b1c1",x"404e",x"3710",x"37bd",x"3b00",x"0000",x"3a5a",x"3b5d",x"b1c1",x"404e",x"36da",x"3680",x"3b4f",x"8000",x"3a50",x"3b5d",x"b1a1",x"404d",x"3710",x"314c",x"3be3",x"0000",x"3a5a",x"3b60"),
(x"b7a4",x"4038",x"3710",x"b64a",x"bb5a",x"8000",x"3a7c",x"3b00",x"b7a4",x"4038",x"36da",x"b654",x"bb58",x"8000",x"3a72",x"3b00",x"b7c7",x"4039",x"3710",x"b744",x"bb20",x"868d",x"3a7c",x"3b07"),
(x"b721",x"404f",x"3710",x"3711",x"bb2d",x"0000",x"3a93",x"3b10",x"b721",x"404f",x"36da",x"37a6",x"bb06",x"0000",x"3a88",x"3b10",x"b72e",x"404e",x"3710",x"39a7",x"b9a8",x"0000",x"3a93",x"3b13"),
(x"b326",x"4043",x"3710",x"ad8e",x"bbf8",x"0000",x"3a5a",x"3bac",x"b326",x"4043",x"36da",x"a5e9",x"bbff",x"0000",x"3a50",x"3bac",x"b34f",x"4043",x"3710",x"3448",x"bbb5",x"0000",x"3a5a",x"3bb0"),
(x"b1a1",x"404d",x"3710",x"314c",x"3be3",x"0000",x"3a5a",x"3b60",x"b1a1",x"404d",x"36da",x"2ede",x"3bf4",x"0000",x"3a50",x"3b60",x"b161",x"404d",x"3710",x"30d8",x"3be8",x"8000",x"3a5a",x"3b66"),
(x"b783",x"4036",x"3710",x"afa0",x"bbf1",x"0000",x"3a7c",x"3af9",x"b783",x"4036",x"36da",x"b33d",x"bbca",x"8000",x"3a72",x"3af9",x"b7a4",x"4038",x"3710",x"b64a",x"bb5a",x"8000",x"3a7c",x"3b00"),
(x"b72e",x"404e",x"3710",x"39a7",x"b9a8",x"0000",x"3a96",x"3b18",x"b72e",x"404e",x"36da",x"3b4f",x"b67e",x"8000",x"3a8b",x"3b18",x"b72d",x"404d",x"3710",x"3a45",x"38f8",x"0000",x"3a96",x"3b19"),
(x"b2d6",x"4043",x"3710",x"b4dc",x"bb9f",x"0000",x"3a5a",x"3ba5",x"b2d6",x"4043",x"36da",x"b287",x"bbd4",x"0000",x"3a50",x"3ba5",x"b326",x"4043",x"3710",x"ad8e",x"bbf8",x"0000",x"3a5a",x"3bac"),
(x"b161",x"404d",x"3710",x"30d8",x"3be8",x"8000",x"3a5a",x"3b66",x"b161",x"404d",x"36da",x"3407",x"3bbe",x"0000",x"3a50",x"3b66",x"b135",x"404c",x"3710",x"3822",x"3ad9",x"0000",x"3a5a",x"3b6a"),
(x"b73e",x"4035",x"3710",x"2f55",x"bbf2",x"0000",x"3a7c",x"3aec",x"b73e",x"4035",x"36da",x"27ae",x"bbff",x"0000",x"3a72",x"3aec",x"b783",x"4036",x"3710",x"afa0",x"bbf1",x"0000",x"3a7c",x"3af9"),
(x"b72d",x"404d",x"3710",x"3a45",x"38f8",x"0000",x"3a96",x"3b19",x"b72d",x"404d",x"36da",x"3778",x"3b13",x"0000",x"3a8b",x"3b19",x"b721",x"404c",x"3710",x"2560",x"3bff",x"0000",x"3a96",x"3b1c"),
(x"b2aa",x"4041",x"3710",x"b7e2",x"baf5",x"0000",x"3a5a",x"3ba0",x"b2aa",x"4041",x"36da",x"b78b",x"bb0e",x"0000",x"3a50",x"3ba0",x"b2d6",x"4043",x"3710",x"b4dc",x"bb9f",x"0000",x"3a5a",x"3ba5"),
(x"b135",x"404c",x"3710",x"3822",x"3ad9",x"0000",x"3a5a",x"3b6a",x"b135",x"404c",x"36da",x"3934",x"3a13",x"8000",x"3a50",x"3b6a",x"b116",x"404a",x"3710",x"3b51",x"3675",x"0000",x"3a5a",x"3b6f"),
(x"b705",x"4037",x"3710",x"36ee",x"bb35",x"0000",x"3a7c",x"3ae1",x"b705",x"4037",x"36da",x"34b8",x"bba4",x"8000",x"3a72",x"3ae1",x"b73e",x"4035",x"3710",x"2f55",x"bbf2",x"0000",x"3a7c",x"3aec"),
(x"b575",x"4056",x"3710",x"bb97",x"350c",x"8000",x"3a96",x"3b79",x"b575",x"4056",x"36da",x"bab5",x"385c",x"8000",x"3a8b",x"3b79",x"b568",x"4058",x"3710",x"b919",x"3a29",x"0000",x"3a96",x"3b7d"),
(x"b938",x"4042",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"39be",x"b938",x"4042",x"36da",x"bbfe",x"a8f0",x"0000",x"3bea",x"39c8",x"b93a",x"404d",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3bfb",x"39bf"),
(x"b261",x"403f",x"3710",x"b5e0",x"bb70",x"8000",x"3a5a",x"3b98",x"b261",x"403f",x"36da",x"b72e",x"bb26",x"0000",x"3a50",x"3b98",x"b2aa",x"4041",x"3710",x"b7e2",x"baf5",x"0000",x"3a5a",x"3ba0"),
(x"b931",x"4059",x"3710",x"2418",x"3bff",x"1a24",x"3a23",x"3bb3",x"b931",x"4059",x"36da",x"23ae",x"3bff",x"0000",x"3a2d",x"3bb3",x"b8ff",x"4059",x"3710",x"257a",x"3bff",x"15bc",x"3a23",x"3b9f"),
(x"b6f1",x"4039",x"3710",x"3b73",x"b5d3",x"0000",x"3a7c",x"3adc",x"b6f1",x"4039",x"36da",x"3a69",x"b8c9",x"868d",x"3a72",x"3adc",x"b705",x"4037",x"3710",x"36ee",x"bb35",x"0000",x"3a7c",x"3ae1"),
(x"b721",x"404c",x"3710",x"2560",x"3bff",x"0000",x"3a96",x"3b1c",x"b721",x"404c",x"36da",x"0cea",x"3c00",x"0000",x"3a8b",x"3b1c",x"b669",x"404d",x"3710",x"a666",x"3bff",x"0000",x"3a96",x"3b3e"),
(x"b22d",x"403e",x"3710",x"2c28",x"bbfb",x"0000",x"3a5a",x"3b93",x"b22d",x"403e",x"36da",x"ae8a",x"bbf5",x"8000",x"3a50",x"3b93",x"b261",x"403f",x"3710",x"b5e0",x"bb70",x"8000",x"3a5a",x"3b98"),
(x"b6ef",x"403c",x"3710",x"3b57",x"3658",x"8000",x"3a7c",x"3ad8",x"b6ef",x"403c",x"36da",x"3be9",x"30b7",x"868d",x"3a72",x"3ad8",x"b6f1",x"4039",x"3710",x"3b73",x"b5d3",x"0000",x"3a7c",x"3adc"),
(x"b669",x"404d",x"3710",x"a666",x"3bff",x"0000",x"3a96",x"3b3e",x"b669",x"404d",x"36da",x"abae",x"3bfc",x"8000",x"3a8b",x"3b3e",x"b63d",x"404e",x"3710",x"affc",x"3bf0",x"0000",x"3a96",x"3b47"),
(x"b930",x"4041",x"3710",x"b700",x"bb23",x"2f0f",x"3b1b",x"3887",x"b930",x"4041",x"36da",x"b67a",x"bb50",x"0000",x"3b21",x"387e",x"b938",x"4042",x"3710",x"b678",x"bb4d",x"2af6",x"3b19",x"3884"),
(x"a165",x"3ee0",x"36eb",x"bbf4",x"2d6d",x"ac2c",x"3917",x"3210",x"a379",x"3ee5",x"36eb",x"bba3",x"b453",x"2fdf",x"3919",x"31f6",x"a1bd",x"3ee0",x"3715",x"bbf4",x"2da3",x"2b3e",x"390d",x"31fc"),
(x"a271",x"3ee5",x"3718",x"bbb8",x"b22d",x"31b0",x"390e",x"31e7",x"a379",x"3ee5",x"36eb",x"bba3",x"b453",x"2fdf",x"3919",x"31f6",x"a303",x"3eed",x"3715",x"bbda",x"2e4f",x"312f",x"3911",x"31c8"),
(x"a303",x"3eed",x"3715",x"bbda",x"2e4f",x"312f",x"3911",x"31c8",x"a3d0",x"3eed",x"36eb",x"bb7a",x"3531",x"30a8",x"391c",x"31d5",x"a0f3",x"3ef4",x"3714",x"ba0a",x"3915",x"3126",x"3914",x"31a4"),
(x"a0f3",x"3ef4",x"3714",x"ba0a",x"3915",x"3126",x"3914",x"31a4",x"a133",x"3ef6",x"36eb",x"b8c7",x"3a49",x"310c",x"391e",x"31a8",x"96c5",x"3ef8",x"3714",x"b236",x"3bc0",x"30e1",x"3915",x"317d"),
(x"96c5",x"3ef8",x"3714",x"b236",x"3bc0",x"30e1",x"3915",x"317d",x"9725",x"3efa",x"36eb",x"a3ae",x"3bec",x"3065",x"391f",x"3181",x"21e6",x"3ef7",x"3714",x"335f",x"3baf",x"30fd",x"3916",x"3143"),
(x"21e6",x"3ef7",x"3714",x"335f",x"3baf",x"30fd",x"3916",x"3143",x"22b9",x"3ef8",x"36eb",x"36e0",x"3b1c",x"3118",x"3920",x"313f",x"24a4",x"3ef1",x"3715",x"3a37",x"38de",x"311d",x"3915",x"311d"),
(x"24a4",x"3ef1",x"3715",x"3a37",x"38de",x"311d",x"3915",x"311d",x"2505",x"3ef2",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3920",x"3117",x"252e",x"3eea",x"3715",x"3bf2",x"2495",x"2f43",x"3914",x"30fc"),
(x"256c",x"3eea",x"36eb",x"3bf7",x"2138",x"2dcf",x"391f",x"30f5",x"250e",x"3ee3",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"391d",x"30d7",x"252e",x"3eea",x"3715",x"3bf2",x"2495",x"2f43",x"3914",x"30fc"),
(x"250e",x"3ee3",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"391d",x"30d7",x"2470",x"3ede",x"36eb",x"3bfd",x"212b",x"29e6",x"391c",x"30c1",x"24bc",x"3ee3",x"3715",x"3b87",x"b537",x"2d81",x"3913",x"30de"),
(x"24de",x"3ec4",x"3717",x"3be8",x"30a2",x"2973",x"390d",x"305d",x"250d",x"3ec4",x"36eb",x"3b9b",x"34d2",x"2ca7",x"3917",x"3054",x"25c0",x"3ec2",x"3714",x"3b74",x"35a6",x"2d5e",x"390d",x"304b"),
(x"20e0",x"3edf",x"3718",x"bbf1",x"95bc",x"2fb4",x"392d",x"2d20",x"2066",x"3edf",x"36eb",x"bbf7",x"9e73",x"2dbc",x"392c",x"2cc6",x"20c8",x"3ee4",x"3716",x"bbad",x"3434",x"2e8a",x"3928",x"2d1c"),
(x"2116",x"3ec2",x"3718",x"ba6d",x"3838",x"3468",x"394c",x"2d1c",x"2029",x"3ec5",x"36eb",x"ba79",x"3840",x"3401",x"3948",x"2cc1",x"20e0",x"3edf",x"3718",x"bbf1",x"95bc",x"2fb4",x"392d",x"2d20"),
(x"a4d5",x"3eb8",x"3715",x"b3c8",x"bbc2",x"235f",x"38fc",x"32a0",x"a50e",x"3eb9",x"36eb",x"b409",x"bbbc",x"27db",x"3905",x"32b4",x"a4b5",x"3ec3",x"3715",x"bbb4",x"33e8",x"2ed7",x"3900",x"3276"),
(x"25ec",x"3ec3",x"36eb",x"3b76",x"3593",x"2dee",x"3917",x"3044",x"262b",x"3eb8",x"36eb",x"36d0",x"bb39",x"2aae",x"3914",x"3017",x"25c0",x"3ec2",x"3714",x"3b74",x"35a6",x"2d5e",x"390d",x"304b"),
(x"993e",x"3edf",x"3716",x"3bce",x"b2bb",x"2b41",x"38fa",x"2d2d",x"9909",x"3ee3",x"3715",x"3b88",x"3531",x"2dc2",x"38ff",x"2d27",x"9651",x"3ee0",x"36eb",x"3bd3",x"b208",x"2da6",x"38fa",x"2cd5"),
(x"9db7",x"3ee9",x"3717",x"3bd6",x"323b",x"2a8a",x"3905",x"2d2c",x"9caa",x"3ee8",x"36ee",x"3b20",x"3725",x"2d51",x"3904",x"2cda",x"9909",x"3ee3",x"3715",x"3b88",x"3531",x"2dc2",x"38ff",x"2d27"),
(x"9cfd",x"3eed",x"3716",x"3aa6",x"b86c",x"2baa",x"390a",x"2d29",x"9cff",x"3eec",x"36ee",x"3b1d",x"b747",x"2911",x"3909",x"2cda",x"9db7",x"3ee9",x"3717",x"3bd6",x"323b",x"2a8a",x"3905",x"2d2c"),
(x"21f4",x"3eec",x"3714",x"bb34",x"b6e6",x"2b2e",x"391f",x"2d20",x"219c",x"3eec",x"36ee",x"ba30",x"b90f",x"2921",x"391e",x"2cd4",x"1f52",x"3ef0",x"3715",x"b638",x"bb5e",x"243f",x"3918",x"2d23"),
(x"9651",x"3ee0",x"36eb",x"3bd3",x"b208",x"2da6",x"38fa",x"2cd5",x"9fcf",x"3ec6",x"36eb",x"3be6",x"2cac",x"3077",x"38de",x"2ce5",x"993e",x"3edf",x"3716",x"3bce",x"b2bb",x"2b41",x"38fa",x"2d2d"),
(x"25f4",x"3eb9",x"3714",x"2745",x"ad9b",x"3bf7",x"3997",x"3194",x"24de",x"3ec4",x"3717",x"2984",x"a0c2",x"3bfd",x"3995",x"31ae",x"25c0",x"3ec2",x"3714",x"33e6",x"2587",x"3bc0",x"3997",x"31a9"),
(x"a4b5",x"3ec3",x"3715",x"b3f3",x"1d38",x"3bbf",x"397f",x"31ac",x"a3f1",x"3ec4",x"3718",x"a6a1",x"97c8",x"3bff",x"3981",x"31ad",x"a4d5",x"3eb8",x"3715",x"a081",x"ad9e",x"3bf8",x"397f",x"3194"),
(x"a271",x"3ee5",x"3718",x"28fa",x"a4f7",x"3bfe",x"3983",x"31f6",x"9909",x"3ee3",x"3715",x"28d3",x"a80e",x"3bfd",x"3988",x"31f3",x"a1bd",x"3ee0",x"3715",x"a1a1",x"23fc",x"3bff",x"3983",x"31eb"),
(x"a303",x"3eed",x"3715",x"9ec2",x"2bd5",x"3bfc",x"3982",x"3208",x"9db7",x"3ee9",x"3717",x"250b",x"281b",x"3bfe",x"3987",x"31ff",x"a271",x"3ee5",x"3718",x"28fa",x"a4f7",x"3bfe",x"3983",x"31f6"),
(x"a0f3",x"3ef4",x"3714",x"263f",x"27c8",x"3bfe",x"3984",x"3218",x"9cfd",x"3eed",x"3716",x"252b",x"2c96",x"3bfa",x"3987",x"3208",x"a303",x"3eed",x"3715",x"9ec2",x"2bd5",x"3bfc",x"3982",x"3208"),
(x"96c5",x"3ef8",x"3714",x"a194",x"a0dd",x"3bff",x"3989",x"3221",x"94d9",x"3eef",x"3713",x"184d",x"9cd0",x"3c00",x"3989",x"320d",x"a0f3",x"3ef4",x"3714",x"263f",x"27c8",x"3bfe",x"3984",x"3218"),
(x"21e6",x"3ef7",x"3714",x"1df0",x"2487",x"3bff",x"3990",x"321e",x"1f52",x"3ef0",x"3715",x"9cb5",x"191e",x"3c00",x"398e",x"320f",x"96c5",x"3ef8",x"3714",x"a194",x"a0dd",x"3bff",x"3989",x"3221"),
(x"24a4",x"3ef1",x"3715",x"a793",x"184d",x"3bff",x"3994",x"3211",x"21f4",x"3eec",x"3714",x"9da1",x"252b",x"3bff",x"3991",x"3205",x"21e6",x"3ef7",x"3714",x"1df0",x"2487",x"3bff",x"3990",x"321e"),
(x"2211",x"3ee8",x"3716",x"2338",x"267a",x"3bff",x"3991",x"31fe",x"21f4",x"3eec",x"3714",x"9da1",x"252b",x"3bff",x"3991",x"3205",x"252e",x"3eea",x"3715",x"9818",x"26bb",x"3bff",x"3995",x"3201"),
(x"20c8",x"3ee4",x"3716",x"24bc",x"2b17",x"3bfc",x"398f",x"31f4",x"2211",x"3ee8",x"3716",x"2338",x"267a",x"3bff",x"3991",x"31fe",x"24bc",x"3ee3",x"3715",x"2645",x"29e0",x"3bfd",x"3994",x"31f1"),
(x"2464",x"3ede",x"3717",x"27d5",x"236c",x"3bfe",x"3994",x"31e7",x"20e0",x"3edf",x"3718",x"2793",x"243f",x"3bfe",x"398f",x"31ea",x"24bc",x"3ee3",x"3715",x"2645",x"29e0",x"3bfd",x"3994",x"31f1"),
(x"2464",x"3ede",x"3717",x"27d5",x"236c",x"3bfe",x"3994",x"31e7",x"24de",x"3ec4",x"3717",x"2984",x"a0c2",x"3bfd",x"3995",x"31ae",x"20e0",x"3edf",x"3718",x"2793",x"243f",x"3bfe",x"398f",x"31ea"),
(x"2211",x"3ee8",x"3716",x"bba5",x"34a4",x"2a11",x"3922",x"2d21",x"21cf",x"3ee8",x"36ee",x"bb7c",x"357c",x"2d58",x"3921",x"2cd1",x"21f4",x"3eec",x"3714",x"bb34",x"b6e6",x"2b2e",x"391f",x"2d20"),
(x"a3f1",x"3ec4",x"3718",x"bba4",x"33dc",x"313e",x"3900",x"3269",x"a46c",x"3ec5",x"36eb",x"bbaa",x"3475",x"2c25",x"390b",x"327d",x"a1bd",x"3ee0",x"3715",x"bbf4",x"2da3",x"2b3e",x"390d",x"31fc"),
(x"a4fc",x"3ec4",x"36eb",x"bbc6",x"328d",x"2f71",x"390a",x"3287",x"a46c",x"3ec5",x"36eb",x"bbaa",x"3475",x"2c25",x"390b",x"327d",x"a4b5",x"3ec3",x"3715",x"bbb4",x"33e8",x"2ed7",x"3900",x"3276"),
(x"25f4",x"3eb9",x"3714",x"2745",x"ad9b",x"3bf7",x"3997",x"3194",x"2116",x"3ec2",x"3718",x"23ae",x"ac2f",x"3bfb",x"398f",x"31a9",x"24de",x"3ec4",x"3717",x"2984",x"a0c2",x"3bfd",x"3995",x"31ae"),
(x"a069",x"3ec3",x"3718",x"a24c",x"a379",x"3bff",x"3985",x"31ab",x"2116",x"3ec2",x"3718",x"23ae",x"ac2f",x"3bfb",x"398f",x"31a9",x"a4d5",x"3eb8",x"3715",x"a081",x"ad9e",x"3bf8",x"397f",x"3194"),
(x"a3f1",x"3ec4",x"3718",x"a6a1",x"97c8",x"3bff",x"3981",x"31ad",x"a069",x"3ec3",x"3718",x"a24c",x"a379",x"3bff",x"3985",x"31ab",x"a4d5",x"3eb8",x"3715",x"a081",x"ad9e",x"3bf8",x"397f",x"3194"),
(x"9cfd",x"3eed",x"3716",x"3aa6",x"b86c",x"2baa",x"390a",x"2d29",x"94d9",x"3eef",x"3713",x"3405",x"bbbe",x"a393",x"390f",x"2d21",x"9cff",x"3eec",x"36ee",x"3b1d",x"b747",x"2911",x"3909",x"2cda"),
(x"2464",x"3ede",x"3717",x"3bff",x"2481",x"2487",x"3911",x"30ca",x"2470",x"3ede",x"36eb",x"3bfd",x"212b",x"29e6",x"391c",x"30c1",x"24de",x"3ec4",x"3717",x"3be8",x"30a2",x"2973",x"390d",x"305d"),
(x"1f52",x"3ef0",x"3715",x"b638",x"bb5e",x"243f",x"3918",x"2d23",x"1f13",x"3ef0",x"36ee",x"b188",x"bbe0",x"a53f",x"3917",x"2cd5",x"94d9",x"3eef",x"3713",x"3405",x"bbbe",x"a393",x"390f",x"2d21"),
(x"9fcf",x"3ec6",x"36eb",x"3be6",x"2cac",x"3077",x"38de",x"2ce5",x"2029",x"3ec5",x"36eb",x"ba79",x"3840",x"3401",x"38cd",x"2cc1",x"a069",x"3ec3",x"3718",x"398b",x"396b",x"33db",x"38db",x"2d41"),
(x"262b",x"3eb8",x"36eb",x"36d0",x"bb39",x"2aae",x"3914",x"3017",x"a50e",x"3eb9",x"36eb",x"b409",x"bbbc",x"27db",x"3905",x"2ec4",x"25f4",x"3eb9",x"3714",x"2f03",x"bbf3",x"23ef",x"390b",x"3022"),
(x"2211",x"3ee8",x"3716",x"bba5",x"34a4",x"2a11",x"3922",x"2d21",x"20c8",x"3ee4",x"3716",x"bbad",x"3434",x"2e8a",x"3928",x"2d1c",x"21cf",x"3ee8",x"36ee",x"bb7c",x"357c",x"2d58",x"3921",x"2cd1"),
(x"9df1",x"3fc7",x"3715",x"2d56",x"20d0",x"3bf8",x"3bad",x"3b15",x"91f4",x"3fd4",x"3716",x"30f9",x"a8af",x"3be5",x"3ba8",x"3b0a",x"20f7",x"3fcc",x"370e",x"2fd2",x"2717",x"3bef",x"3ba1",x"3b12"),
(x"9df1",x"3fc7",x"3715",x"bbc5",x"2b9a",x"3358",x"3b3e",x"38e9",x"a03c",x"3fc7",x"36eb",x"bb99",x"3315",x"330d",x"3b44",x"38e9",x"91f4",x"3fd4",x"3716",x"badd",x"375a",x"334d",x"3b3f",x"38e1"),
(x"9a85",x"3f8f",x"3713",x"ada3",x"2f15",x"3beb",x"3baf",x"3b45",x"8010",x"3f87",x"3714",x"ac39",x"29a5",x"3bf9",x"3bad",x"3b4b",x"9d28",x"3f8f",x"3712",x"aa69",x"287e",x"3bfc",x"3bb1",x"3b44"),
(x"a273",x"3f87",x"3712",x"aa73",x"2a97",x"3bfa",x"3bb7",x"3b4a",x"a34c",x"3f8d",x"3711",x"a481",x"2546",x"3bff",x"3bb8",x"3b46",x"9ff6",x"3f91",x"3711",x"a994",x"2977",x"3bfc",x"3bb3",x"3b42"),
(x"9ff6",x"3f91",x"3711",x"a994",x"2977",x"3bfc",x"3bb3",x"3b42",x"9d28",x"3f8f",x"3712",x"aa69",x"287e",x"3bfc",x"3bb1",x"3b44",x"a273",x"3f87",x"3712",x"aa73",x"2a97",x"3bfa",x"3bb7",x"3b4a"),
(x"9e8d",x"3f84",x"3716",x"af14",x"329b",x"3bc7",x"3bb2",x"3b4e",x"9c36",x"3f82",x"3718",x"ae36",x"a160",x"3bf6",x"3bb0",x"3b4f",x"a17b",x"3f81",x"3711",x"afec",x"ac2c",x"3beb",x"3bb6",x"3b4f"),
(x"9c14",x"3f6f",x"370f",x"2b8a",x"30ae",x"3be6",x"3bb1",x"3b60",x"a035",x"3f6a",x"3713",x"ae9c",x"3366",x"3bbd",x"3bb5",x"3b64",x"9c56",x"3f71",x"370e",x"26d5",x"25c2",x"3bfe",x"3bb1",x"3b5e"),
(x"a425",x"3f70",x"370f",x"acd8",x"a71d",x"3bf9",x"3bbb",x"3b5e",x"9f72",x"3f76",x"3713",x"a538",x"ac79",x"3bfa",x"3bb4",x"3b59",x"a289",x"3f6b",x"370f",x"9df0",x"a631",x"3bff",x"3bb9",x"3b62"),
(x"a425",x"3f70",x"370f",x"acd8",x"a71d",x"3bf9",x"3bbb",x"3b5e",x"a407",x"3f79",x"370f",x"aec5",x"1a59",x"3bf4",x"3bba",x"3b56",x"9f72",x"3f76",x"3713",x"a538",x"ac79",x"3bfa",x"3bb4",x"3b59"),
(x"a17b",x"3f81",x"3711",x"afec",x"ac2c",x"3beb",x"3bb6",x"3b4f",x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53",x"9d1a",x"3f7a",x"3710",x"ac5b",x"b0a5",x"3be5",x"3bb1",x"3b56"),
(x"1d4c",x"3f53",x"3717",x"97c8",x"9f79",x"3c00",x"3ba9",x"3b76",x"1e77",x"3f4b",x"3715",x"a6c2",x"ac63",x"3bfa",x"3ba8",x"3b7e",x"19fe",x"3f52",x"3717",x"aff2",x"aa7d",x"3bed",x"3bab",x"3b78"),
(x"a2cb",x"3f51",x"3714",x"1553",x"ab62",x"3bfc",x"3bb8",x"3b78",x"a38f",x"3f55",x"3712",x"b163",x"a345",x"3be2",x"3bb9",x"3b75",x"a13d",x"3f5b",x"3716",x"acd8",x"a7e2",x"3bf9",x"3bb5",x"3b70"),
(x"a13d",x"3f5b",x"3716",x"acd8",x"a7e2",x"3bf9",x"3bb5",x"3b70",x"9e62",x"3f5a",x"3716",x"2818",x"ad04",x"3bf8",x"3bb2",x"3b71",x"a2cb",x"3f51",x"3714",x"1553",x"ab62",x"3bfc",x"3bb8",x"3b78"),
(x"987a",x"3f57",x"3714",x"a4fd",x"ada9",x"3bf7",x"3baf",x"3b74",x"9d1e",x"3f4e",x"3711",x"240b",x"ad5c",x"3bf8",x"3bb1",x"3b7b",x"9e62",x"3f5a",x"3716",x"2818",x"ad04",x"3bf8",x"3bb2",x"3b71"),
(x"0e53",x"3f54",x"3714",x"b036",x"a73e",x"3bed",x"3bad",x"3b76",x"19fe",x"3f52",x"3717",x"aff2",x"aa7d",x"3bed",x"3bab",x"3b78",x"9a71",x"3f4c",x"3711",x"b27d",x"16f6",x"3bd5",x"3bb0",x"3b7c"),
(x"a16d",x"3f34",x"3711",x"b115",x"27d5",x"3be4",x"3bb6",x"3b90",x"9ae8",x"3f45",x"3712",x"b146",x"2c91",x"3bde",x"3bb0",x"3b82",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f"),
(x"1e3f",x"3f34",x"3715",x"28bf",x"afdb",x"3bef",x"3ba9",x"3b91",x"1f1f",x"3f39",x"3718",x"2138",x"ae95",x"3bf4",x"3ba8",x"3b8c",x"21e0",x"3f38",x"3719",x"a90e",x"af00",x"3bf2",x"3ba5",x"3b8d"),
(x"1e3f",x"3f34",x"3715",x"28bf",x"afdb",x"3bef",x"3ba9",x"3b91",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f",x"1f1f",x"3f39",x"3718",x"2138",x"ae95",x"3bf4",x"3ba8",x"3b8c"),
(x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"1e5a",x"3f3a",x"3718",x"2b4f",x"2525",x"3bfc",x"3ba9",x"3b8b",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f"),
(x"20ca",x"3f3e",x"3715",x"2d65",x"ac5a",x"3bf3",x"3ba6",x"3b89",x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"2288",x"3f43",x"3718",x"2cf2",x"18ea",x"3bf9",x"3ba3",x"3b85"),
(x"2257",x"3f49",x"3712",x"3542",x"30b9",x"3b76",x"3ba4",x"3b7f",x"22dc",x"3f47",x"3712",x"359c",x"336a",x"3b42",x"3ba3",x"3b81",x"2091",x"3f49",x"3717",x"2d2f",x"2ecb",x"3bed",x"3ba6",x"3b80"),
(x"2091",x"3f49",x"3717",x"2d2f",x"2ecb",x"3bed",x"3ba6",x"3b80",x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"1f4b",x"3f49",x"3716",x"b009",x"2da6",x"3be7",x"3ba8",x"3b7f"),
(x"1e77",x"3f4b",x"3715",x"a6c2",x"ac63",x"3bfa",x"3ba8",x"3b7e",x"1f4b",x"3f49",x"3716",x"b009",x"2da6",x"3be7",x"3ba8",x"3b7f",x"990c",x"3f4b",x"3712",x"af67",x"a981",x"3bf0",x"3baf",x"3b7e"),
(x"1f29",x"3f4d",x"3714",x"a57a",x"ae8a",x"3bf4",x"3ba8",x"3b7c",x"1e77",x"3f4b",x"3715",x"a6c2",x"ac63",x"3bfa",x"3ba8",x"3b7e",x"1d4c",x"3f53",x"3717",x"97c8",x"9f79",x"3c00",x"3ba9",x"3b76"),
(x"2147",x"3f51",x"3718",x"ac00",x"290e",x"3bfa",x"3ba5",x"3b79",x"20ef",x"3f58",x"3715",x"a51e",x"2d06",x"3bf9",x"3ba6",x"3b73",x"2442",x"3f5d",x"3714",x"175f",x"2c2c",x"3bfb",x"3ba0",x"3b6f"),
(x"2442",x"3f5d",x"3714",x"175f",x"2c2c",x"3bfb",x"3ba0",x"3b6f",x"2308",x"3f60",x"3714",x"2dba",x"2266",x"3bf7",x"3ba3",x"3b6c",x"24cc",x"3f69",x"3712",x"3106",x"273e",x"3be5",x"3b9f",x"3b64"),
(x"24cc",x"3f69",x"3712",x"3106",x"273e",x"3be5",x"3b9f",x"3b64",x"2365",x"3f6b",x"3715",x"3468",x"247a",x"3bb0",x"3ba2",x"3b63",x"243c",x"3f75",x"3710",x"3550",x"2e33",x"3b81",x"3ba0",x"3b5a"),
(x"243c",x"3f75",x"3710",x"3550",x"2e33",x"3b81",x"3ba0",x"3b5a",x"22bc",x"3f73",x"3717",x"3273",x"2f43",x"3bc8",x"3ba3",x"3b5c",x"21ba",x"3f7d",x"3712",x"2b5c",x"2345",x"3bfc",x"3ba5",x"3b54"),
(x"21ba",x"3f7d",x"3712",x"2b5c",x"2345",x"3bfc",x"3ba5",x"3b54",x"1f35",x"3f7a",x"3711",x"ae24",x"2a2b",x"3bf4",x"3ba8",x"3b56",x"1a19",x"3f7b",x"3712",x"2dd2",x"b04b",x"3be4",x"3bab",x"3b55"),
(x"9588",x"3f84",x"3716",x"a559",x"32c7",x"3bd1",x"3bae",x"3b4d",x"08f2",x"3f83",x"3716",x"2f4b",x"aa5f",x"3bf0",x"3bad",x"3b4f",x"9c36",x"3f82",x"3718",x"ae36",x"a160",x"3bf6",x"3bb0",x"3b4f"),
(x"9588",x"3f84",x"3716",x"a559",x"32c7",x"3bd1",x"3bae",x"3b4d",x"9c36",x"3f82",x"3718",x"ae36",x"a160",x"3bf6",x"3bb0",x"3b4f",x"9e8d",x"3f84",x"3716",x"af14",x"329b",x"3bc7",x"3bb2",x"3b4e"),
(x"8010",x"3f87",x"3714",x"ac39",x"29a5",x"3bf9",x"3bad",x"3b4b",x"9a85",x"3f8f",x"3713",x"ada3",x"2f15",x"3beb",x"3baf",x"3b45",x"1f40",x"3f8e",x"3717",x"b0e7",x"3057",x"3bd4",x"3ba7",x"3b45"),
(x"1f40",x"3f8e",x"3717",x"b0e7",x"3057",x"3bd4",x"3ba7",x"3b45",x"1820",x"3f93",x"370f",x"aedc",x"2cd0",x"3bee",x"3bab",x"3b41",x"221f",x"3f9c",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3ba3",x"3b3a"),
(x"221f",x"3f9c",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3ba3",x"3b3a",x"1d56",x"3f9e",x"3716",x"aadf",x"a6b5",x"3bfc",x"3ba8",x"3b38",x"2273",x"3faa",x"3717",x"abf6",x"25ae",x"3bfb",x"3ba1",x"3b2f"),
(x"2273",x"3faa",x"3717",x"abf6",x"25ae",x"3bfb",x"3ba1",x"3b2f",x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21",x"2386",x"3fb5",x"370f",x"36ca",x"2fac",x"3b2e",x"3b9e",x"3b26"),
(x"2243",x"3fba",x"3713",x"2f9d",x"b907",x"3a26",x"3ba0",x"3b21",x"2312",x"3fb8",x"370d",x"3809",x"2e09",x"3add",x"3b9f",x"3b23",x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21"),
(x"20f7",x"3fcc",x"370e",x"2fd2",x"2717",x"3bef",x"3ba1",x"3b12",x"21a5",x"3fc1",x"3712",x"29f0",x"2b1d",x"3bfa",x"3ba1",x"3b1b",x"9df1",x"3fc7",x"3715",x"2d56",x"20d0",x"3bf8",x"3bad",x"3b15"),
(x"9cbb",x"3fba",x"3715",x"bb81",x"b440",x"330f",x"3b3e",x"38ef",x"1882",x"3fa8",x"370e",x"bb5f",x"b5f1",x"2f4f",x"3b3c",x"38f9",x"9f02",x"3fb9",x"36eb",x"bb89",x"b473",x"31fc",x"3b43",x"38f0"),
(x"a122",x"3f23",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3b85",x"39fe",x"a167",x"3f14",x"36eb",x"3bf5",x"2e59",x"2467",x"3b86",x"3a06",x"a175",x"3f1a",x"3710",x"3bfd",x"a997",x"a0a8",x"3b8a",x"3a03"),
(x"8dee",x"3f36",x"36eb",x"b469",x"bb91",x"316a",x"3b85",x"39f3",x"a122",x"3f23",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3b85",x"39fe",x"9c3a",x"3f30",x"3714",x"3b1c",x"b754",x"223f",x"3b8a",x"39f7"),
(x"a167",x"3f14",x"36eb",x"3bf5",x"2e59",x"2467",x"3b86",x"3a06",x"a051",x"3f0c",x"36eb",x"3ab1",x"3862",x"21e3",x"3b86",x"3a0a",x"a099",x"3f0e",x"3712",x"3b76",x"35c5",x"204d",x"3b8a",x"3a09"),
(x"a051",x"3f0c",x"36eb",x"3ab1",x"3862",x"21e3",x"3b86",x"3a0a",x"9b3f",x"3f08",x"36eb",x"37e1",x"3af5",x"269a",x"3b86",x"3a0d",x"9ecc",x"3f0b",x"3714",x"395a",x"39f1",x"2025",x"3b8b",x"3a0b"),
(x"9b3f",x"3f08",x"36eb",x"37e1",x"3af5",x"269a",x"3b86",x"3a0d",x"197e",x"3f07",x"36eb",x"303c",x"3beb",x"299e",x"3b86",x"3a11",x"9aa8",x"3f08",x"3714",x"35bf",x"3b76",x"27db",x"3b8b",x"3a0d"),
(x"197e",x"3f07",x"36eb",x"303c",x"3beb",x"299e",x"3b86",x"3a11",x"20a0",x"3f08",x"36eb",x"b868",x"3aab",x"296a",x"3b86",x"3a14",x"1a1e",x"3f06",x"3715",x"a836",x"3bfd",x"294f",x"3b8b",x"3a11"),
(x"20b2",x"3f08",x"3716",x"b86f",x"3aa7",x"2604",x"3b8b",x"3a14",x"20a0",x"3f08",x"36eb",x"b868",x"3aab",x"296a",x"3b86",x"3a14",x"2335",x"3f0e",x"3714",x"bb01",x"37b5",x"2839",x"3b8b",x"3a18"),
(x"2300",x"3f0e",x"36eb",x"baf3",x"37df",x"2b38",x"3b86",x"3a18",x"23d0",x"3f13",x"36eb",x"bbf9",x"2d11",x"2511",x"3b85",x"3a1b",x"2335",x"3f0e",x"3714",x"bb01",x"37b5",x"2839",x"3b8b",x"3a18"),
(x"23d0",x"3f13",x"36eb",x"bbf9",x"2d11",x"2511",x"3b85",x"3a1b",x"2300",x"3f18",x"36eb",x"b90c",x"ba34",x"2532",x"3b85",x"3a1e",x"23d3",x"3f13",x"3714",x"bbe6",x"b10f",x"9bfc",x"3b8b",x"3a1b"),
(x"22d3",x"3f18",x"3715",x"b928",x"ba1d",x"1553",x"3a62",x"3a41",x"2300",x"3f18",x"36eb",x"b90c",x"ba34",x"2532",x"3a68",x"3a42",x"20d5",x"3f18",x"3714",x"2fe4",x"bbee",x"2901",x"3a63",x"3a3f"),
(x"20d5",x"3f18",x"3714",x"2fe4",x"bbee",x"2901",x"3a63",x"3a3f",x"20b2",x"3f18",x"36eb",x"35dd",x"bb6d",x"2be9",x"3a68",x"3a3f",x"1e4f",x"3f16",x"3711",x"364f",x"bb52",x"2d1b",x"3a64",x"3a3d"),
(x"865b",x"3f23",x"36eb",x"b9db",x"396c",x"2c1a",x"3a69",x"3a32",x"13e1",x"3f25",x"36eb",x"bbf6",x"2a70",x"2d61",x"3a69",x"3a31",x"3d81",x"3f23",x"3711",x"ba7a",x"38b0",x"2839",x"3a64",x"3a33"),
(x"1e4f",x"3f16",x"3711",x"364f",x"bb52",x"2d1b",x"3a64",x"3a3d",x"1ead",x"3f15",x"36eb",x"32b1",x"bbc8",x"2e54",x"3a68",x"3a3d",x"14bb",x"3f16",x"3710",x"b416",x"bbad",x"2f8d",x"3a64",x"3a3b"),
(x"998f",x"3f6e",x"36eb",x"3b7d",x"b521",x"3095",x"3b28",x"3928",x"9f83",x"3f68",x"36eb",x"35e4",x"bb4d",x"31a2",x"3b2b",x"3927",x"9c14",x"3f6f",x"370f",x"3a9b",x"b854",x"30fa",x"3b26",x"3924"),
(x"9cbb",x"3fba",x"3715",x"bb81",x"b440",x"330f",x"3b3e",x"38ef",x"9f02",x"3fb9",x"36eb",x"bb89",x"b473",x"31fc",x"3b43",x"38f0",x"9df1",x"3fc7",x"3715",x"bbc5",x"2b9a",x"3358",x"3b3e",x"38e9"),
(x"2375",x"3f22",x"3711",x"a8d9",x"a52b",x"3bfe",x"3ba2",x"3ba0",x"983c",x"3f20",x"3710",x"a856",x"a9ab",x"3bfc",x"3bb0",x"3ba1",x"1f0f",x"3f25",x"3718",x"ab65",x"b528",x"3b8f",x"3ba8",x"3b9d"),
(x"210e",x"3fbb",x"36eb",x"3be3",x"2ce8",x"30c3",x"3b3c",x"38cf",x"20f8",x"3fba",x"3716",x"38de",x"3a57",x"297d",x"3b38",x"38d2",x"20d5",x"3fbc",x"3715",x"3bd7",x"b1f9",x"2c2a",x"3b38",x"38d3"),
(x"21ba",x"3f7d",x"3712",x"384e",x"3ab0",x"2ec8",x"3b30",x"3b43",x"2267",x"3f7e",x"36eb",x"3958",x"39de",x"2fdf",x"3b35",x"3b43",x"243c",x"3f75",x"3710",x"3b6a",x"35bb",x"2efe",x"3b31",x"3b3e"),
(x"0f13",x"3f15",x"36eb",x"b37e",x"bbba",x"2ef6",x"3a69",x"3a3a",x"9889",x"3f18",x"36eb",x"baa4",x"b859",x"2fe5",x"3a69",x"3a38",x"14bb",x"3f16",x"3710",x"b416",x"bbad",x"2f8d",x"3a64",x"3a3b"),
(x"1e18",x"3f31",x"36eb",x"3bfa",x"a0b5",x"2cb4",x"3a30",x"3a63",x"1e52",x"3f28",x"36eb",x"3be6",x"308f",x"2c41",x"3a31",x"3a5e",x"1d4f",x"3f31",x"3715",x"3bfa",x"a710",x"2c48",x"3a2b",x"3a61"),
(x"951c",x"3f19",x"3711",x"ba7e",x"b887",x"3089",x"3a64",x"3a39",x"9889",x"3f18",x"36eb",x"baa4",x"b859",x"2fe5",x"3a69",x"3a38",x"99ac",x"3f1c",x"3710",x"bbcc",x"b228",x"2f2f",x"3a64",x"3a37"),
(x"9aca",x"3f71",x"36eb",x"3b19",x"3744",x"2cf7",x"3b27",x"3929",x"998f",x"3f6e",x"36eb",x"3b7d",x"b521",x"3095",x"3b28",x"3928",x"9c56",x"3f71",x"370e",x"3b25",x"370d",x"2d68",x"3b25",x"3924"),
(x"9c70",x"3f4d",x"36eb",x"b7d8",x"baf6",x"2a35",x"3b1d",x"3b24",x"a30f",x"3f4f",x"36eb",x"b6fe",x"bb25",x"2ea4",x"3b1f",x"3b1f",x"9d1e",x"3f4e",x"3711",x"b4dc",x"bb97",x"2d61",x"3b19",x"3b22"),
(x"9a2a",x"3f21",x"36eb",x"bb02",x"3776",x"2fc8",x"3a69",x"3a34",x"865b",x"3f23",x"36eb",x"b9db",x"396c",x"2c1a",x"3a69",x"3a32",x"983c",x"3f20",x"3710",x"bb2f",x"36d9",x"2e52",x"3a64",x"3a35"),
(x"08f2",x"3f83",x"3716",x"37e9",x"3af1",x"2aa7",x"3b2f",x"3b4a",x"8d14",x"3f84",x"36eb",x"3776",x"3b0b",x"2d41",x"3b34",x"3b4b",x"21ba",x"3f7d",x"3712",x"384e",x"3ab0",x"2ec8",x"3b30",x"3b43"),
(x"1e3f",x"3f34",x"3715",x"395d",x"b9e3",x"2de3",x"3a2a",x"3a62",x"1e6c",x"3f33",x"36eb",x"39df",x"b964",x"2d28",x"3a2f",x"3a63",x"1d4f",x"3f31",x"3715",x"3bfa",x"a710",x"2c48",x"3a2b",x"3a61"),
(x"9f72",x"3f76",x"3713",x"3b5b",x"3634",x"2c03",x"3b22",x"3925",x"9f02",x"3f76",x"36eb",x"3ad3",x"3822",x"2c4d",x"3b24",x"392a",x"9c56",x"3f71",x"370e",x"3b25",x"370d",x"2d68",x"3b25",x"3924"),
(x"1d56",x"3f9e",x"3716",x"bbff",x"20c2",x"2138",x"3b3a",x"38ff",x"1d3a",x"3f9d",x"36eb",x"bbfe",x"1e8d",x"2828",x"3b3f",x"3900",x"1882",x"3fa8",x"370e",x"bb5f",x"b5f1",x"2f4f",x"3b3c",x"38f9"),
(x"9427",x"3f84",x"36eb",x"3b23",x"b71d",x"2cde",x"3b34",x"3b4b",x"8d14",x"3f84",x"36eb",x"3776",x"3b0b",x"2d41",x"3b34",x"3b4b",x"9588",x"3f84",x"3716",x"3bde",x"31b5",x"2825",x"3b2e",x"3b4b"),
(x"21e0",x"3f38",x"3719",x"39a6",x"b994",x"2fc6",x"3a29",x"3a66",x"22d4",x"3f38",x"36eb",x"39ed",x"b94b",x"2f45",x"3a2e",x"3a68",x"1e3f",x"3f34",x"3715",x"395d",x"b9e3",x"2de3",x"3a2a",x"3a62"),
(x"9acb",x"3f4a",x"36eb",x"bbf8",x"a379",x"2d44",x"3a2d",x"3a14",x"9c70",x"3f4d",x"36eb",x"b7d8",x"baf6",x"2a35",x"3a2c",x"3a12",x"9a71",x"3f4c",x"3711",x"bb12",x"b763",x"2ca3",x"3a28",x"3a14"),
(x"9f87",x"3f78",x"3713",x"3b09",x"b791",x"2ab8",x"3b21",x"3925",x"9f11",x"3f77",x"36eb",x"39e9",x"b955",x"2e31",x"3b23",x"392a",x"9f72",x"3f76",x"3713",x"3b5b",x"3634",x"2c03",x"3b22",x"3925"),
(x"173f",x"3f94",x"36eb",x"bab4",x"3859",x"2a66",x"3b3e",x"3905",x"1d3a",x"3f9d",x"36eb",x"bbfe",x"1e8d",x"2828",x"3b3f",x"3900",x"1820",x"3f93",x"370f",x"bad7",x"3821",x"29e6",x"3b3a",x"3904"),
(x"141e",x"3f86",x"36eb",x"397a",x"b9b6",x"309a",x"3b26",x"38b9",x"9427",x"3f84",x"36eb",x"3b23",x"b71d",x"2cde",x"3b25",x"38b9",x"8010",x"3f87",x"3714",x"39e8",x"b951",x"2f27",x"3b23",x"38be"),
(x"2283",x"3f3b",x"36eb",x"32cb",x"3bc1",x"2fc5",x"3a2e",x"3a69",x"22d4",x"3f38",x"36eb",x"39ed",x"b94b",x"2f45",x"3a2e",x"3a68",x"21d8",x"3f39",x"3719",x"3250",x"3bca",x"2f22",x"3a29",x"3a66"),
(x"9bea",x"3f46",x"36eb",x"bb57",x"3625",x"2e99",x"3a2d",x"3a16",x"9acb",x"3f4a",x"36eb",x"bbf8",x"a379",x"2d44",x"3a2d",x"3a14",x"9ae8",x"3f45",x"3712",x"bb92",x"3509",x"2cb0",x"3a29",x"3a18"),
(x"9096",x"3f7b",x"36eb",x"3046",x"bbe8",x"2cb7",x"3b1f",x"3af2",x"9f11",x"3f77",x"36eb",x"39e9",x"b955",x"2e31",x"3b1f",x"3aee",x"9d1a",x"3f7a",x"3710",x"3833",x"bac7",x"2d1d",x"3b1b",x"3aef"),
(x"9a85",x"3f8f",x"3713",x"b7c3",x"3af3",x"2e28",x"3b39",x"3908",x"9bdf",x"3f8f",x"36eb",x"b73f",x"3b1a",x"2d3c",x"3b3e",x"3909",x"1820",x"3f93",x"370f",x"bad7",x"3821",x"29e6",x"3b3a",x"3904"),
(x"2078",x"3f8e",x"36eb",x"3aff",x"b73c",x"3197",x"3b2a",x"38bd",x"141e",x"3f86",x"36eb",x"397a",x"b9b6",x"309a",x"3b26",x"38b9",x"1f40",x"3f8e",x"3717",x"3a77",x"b889",x"310e",x"3b27",x"38c1"),
(x"1f1f",x"3f39",x"3718",x"30c5",x"3be6",x"2ad9",x"3a28",x"3a68",x"1e72",x"3f3a",x"36eb",x"3b01",x"3745",x"3141",x"3a2c",x"3a6c",x"21d8",x"3f39",x"3719",x"3250",x"3bca",x"2f22",x"3a29",x"3a66"),
(x"a25f",x"3f33",x"36eb",x"bb99",x"345f",x"30d6",x"3a30",x"3a21",x"9bea",x"3f46",x"36eb",x"bb57",x"3625",x"2e99",x"3a2d",x"3a16",x"a16d",x"3f34",x"3711",x"bb70",x"3585",x"3014",x"3a2c",x"3a21"),
(x"1ecc",x"3f79",x"36eb",x"b74a",x"bb15",x"2de4",x"3b1f",x"3af6",x"9096",x"3f7b",x"36eb",x"3046",x"bbe8",x"2cb7",x"3b1f",x"3af2",x"1a19",x"3f7b",x"3712",x"b2e8",x"bbcb",x"2c10",x"3b1a",x"3af3"),
(x"9d97",x"3f90",x"36eb",x"38ae",x"3a73",x"2d47",x"3b3d",x"390a",x"9bdf",x"3f8f",x"36eb",x"b73f",x"3b1a",x"2d3c",x"3b3e",x"3909",x"9d28",x"3f8f",x"3712",x"3721",x"3b24",x"2bf9",x"3b39",x"3909"),
(x"231e",x"3f9c",x"36eb",x"3bbf",x"b113",x"322d",x"3b30",x"38c2",x"2078",x"3f8e",x"36eb",x"3aff",x"b73c",x"3197",x"3b2a",x"38bd",x"221f",x"3f9c",x"3713",x"3bc6",x"b1be",x"30de",x"3b2c",x"38c6"),
(x"a397",x"3f24",x"36eb",x"bbe6",x"2c77",x"308c",x"3a32",x"3a28",x"a25f",x"3f33",x"36eb",x"bb99",x"345f",x"30d6",x"3a30",x"3a21",x"a2e9",x"3f24",x"3711",x"bbe4",x"2d1d",x"308c",x"3a2e",x"3a2a"),
(x"22bc",x"3f73",x"3717",x"bb6f",x"b5e5",x"261e",x"3b19",x"3afa",x"2284",x"3f73",x"36eb",x"baaf",x"b860",x"2a70",x"3b1f",x"3afa",x"1f35",x"3f7a",x"3711",x"b934",x"ba0d",x"2c16",x"3b1a",x"3af5"),
(x"9f8c",x"3f92",x"36eb",x"2e29",x"3be6",x"3005",x"3b3d",x"390b",x"9d97",x"3f90",x"36eb",x"38ae",x"3a73",x"2d47",x"3b3d",x"390a",x"9ff6",x"3f91",x"3711",x"35dd",x"3b65",x"2eae",x"3b39",x"390b"),
(x"2273",x"3faa",x"3717",x"3bf0",x"af10",x"2aec",x"3b31",x"38cb",x"22be",x"3fa9",x"36eb",x"3bea",x"ae0a",x"2f10",x"3b35",x"38c7",x"221f",x"3f9c",x"3713",x"3bc6",x"b1be",x"30de",x"3b2c",x"38c6"),
(x"1e72",x"3f3a",x"36eb",x"3b01",x"3745",x"3141",x"3b34",x"3b18",x"1f1f",x"3f39",x"3718",x"30c5",x"3be6",x"2ad9",x"3b2e",x"3b19",x"1e5a",x"3f3a",x"3718",x"3af6",x"b7e0",x"2460",x"3b2f",x"3b1a"),
(x"a2ee",x"3f13",x"3714",x"bbec",x"ad02",x"2f4a",x"3a2f",x"3a32",x"a382",x"3f13",x"36eb",x"bbe8",x"ad68",x"3010",x"3a34",x"3a31",x"a2e9",x"3f24",x"3711",x"bbe4",x"2d1d",x"308c",x"3a2e",x"3a2a"),
(x"2365",x"3f6b",x"3715",x"bbfe",x"2412",x"2867",x"3b19",x"3aff",x"234c",x"3f6b",x"36eb",x"bbfa",x"ac62",x"2617",x"3b1f",x"3afe",x"22bc",x"3f73",x"3717",x"bb6f",x"b5e5",x"261e",x"3b19",x"3afa"),
(x"a2ba",x"3f92",x"36eb",x"b913",x"3a0d",x"310f",x"3b3d",x"390e",x"9f8c",x"3f92",x"36eb",x"2e29",x"3be6",x"3005",x"3b3d",x"390b",x"a20d",x"3f91",x"3712",x"b5a5",x"3b63",x"30cc",x"3b38",x"390d"),
(x"2414",x"3fb4",x"36eb",x"3be4",x"aadf",x"30ee",x"3b39",x"38ca",x"22be",x"3fa9",x"36eb",x"3bea",x"ae0a",x"2f10",x"3b35",x"38c7",x"2386",x"3fb5",x"370f",x"3bdd",x"b0de",x"2e6c",x"3b36",x"38ce"),
(x"2349",x"3f43",x"36eb",x"3bbf",x"b333",x"2ed0",x"3b35",x"3b1f",x"21d1",x"3f3e",x"36eb",x"3a0e",x"b929",x"2e76",x"3b35",x"3b1c",x"2288",x"3f43",x"3718",x"3b13",x"b732",x"2fec",x"3b2f",x"3b1f"),
(x"a269",x"3f0a",x"36eb",x"bab2",x"b834",x"30cb",x"3a35",x"3a36",x"a382",x"3f13",x"36eb",x"bbe8",x"ad68",x"3010",x"3a34",x"3a31",x"a1ea",x"3f0b",x"3712",x"bb45",x"b640",x"30a6",x"3a30",x"3a36"),
(x"99ac",x"3f1c",x"3710",x"bbcc",x"b228",x"2f2f",x"3a64",x"3a37",x"9b9c",x"3f1c",x"36eb",x"bbf4",x"9edc",x"2ebb",x"3a69",x"3a36",x"983c",x"3f20",x"3710",x"bb2f",x"36d9",x"2e52",x"3a64",x"3a35"),
(x"2308",x"3f60",x"3714",x"bb81",x"3558",x"2da5",x"3b19",x"3b04",x"22be",x"3f61",x"36eb",x"bbcf",x"32aa",x"2bc5",x"3b1e",x"3b04",x"2365",x"3f6b",x"3715",x"bbfe",x"2412",x"2867",x"3b19",x"3aff"),
(x"a3f7",x"3f8d",x"36eb",x"bbe5",x"adbc",x"3036",x"3b3c",x"3911",x"a2ba",x"3f92",x"36eb",x"b913",x"3a0d",x"310f",x"3b3d",x"390e",x"a34c",x"3f8d",x"3711",x"bbb2",x"332f",x"30f4",x"3b38",x"390f"),
(x"23bf",x"3fba",x"36eb",x"3af6",x"3714",x"32f0",x"3b3b",x"38cd",x"2414",x"3fb4",x"36eb",x"3be4",x"aadf",x"30ee",x"3b39",x"38ca",x"2312",x"3fb8",x"370d",x"3b0d",x"370c",x"3169",x"3b37",x"38cf"),
(x"2324",x"3f48",x"36eb",x"3bbf",x"3371",x"2dad",x"3b35",x"3b21",x"2349",x"3f43",x"36eb",x"3bbf",x"b333",x"2ed0",x"3b35",x"3b1f",x"22dc",x"3f47",x"3712",x"3bf0",x"2c20",x"2e95",x"3b30",x"3b22"),
(x"9dfd",x"3f02",x"36eb",x"b7cb",x"bae6",x"3068",x"3a36",x"3a3b",x"a269",x"3f0a",x"36eb",x"bab2",x"b834",x"30cb",x"3a35",x"3a36",x"9d7f",x"3f04",x"3715",x"b93c",x"b9e9",x"3110",x"3a31",x"3a3c"),
(x"20ef",x"3f58",x"3715",x"ba65",x"38c1",x"2d9c",x"3b19",x"3b09",x"207d",x"3f59",x"36eb",x"bac2",x"3833",x"2e8a",x"3b1f",x"3b09",x"2308",x"3f60",x"3714",x"bb81",x"3558",x"2da5",x"3b19",x"3b04"),
(x"a2c3",x"3f85",x"36eb",x"b902",x"ba23",x"306a",x"3b3a",x"3915",x"a3f7",x"3f8d",x"36eb",x"bbe5",x"adbc",x"3036",x"3b3c",x"3911",x"a273",x"3f87",x"3712",x"bae4",x"b7c3",x"30c9",x"3b36",x"3912"),
(x"2243",x"3fba",x"3713",x"3451",x"3bac",x"2d81",x"3b37",x"38d1",x"226e",x"3fbb",x"36eb",x"3571",x"3b6d",x"30cc",x"3b3b",x"38ce",x"2312",x"3fb8",x"370d",x"3b0d",x"370c",x"3169",x"3b37",x"38cf"),
(x"22c6",x"3f49",x"36eb",x"2eda",x"3bea",x"2e47",x"3b35",x"3b22",x"2324",x"3f48",x"36eb",x"3bbf",x"3371",x"2dad",x"3b35",x"3b21",x"2257",x"3f49",x"3712",x"3297",x"3bcc",x"2d84",x"3b30",x"3b23"),
(x"17aa",x"3f00",x"36eb",x"96f6",x"bbf5",x"2e97",x"3a36",x"3a3f",x"9dfd",x"3f02",x"36eb",x"b7cb",x"bae6",x"3068",x"3a36",x"3a3b",x"17a2",x"3f01",x"3715",x"9ef6",x"bbee",x"302a",x"3a31",x"3a40"),
(x"1d4c",x"3f53",x"3717",x"b939",x"3a0b",x"29e0",x"3b19",x"3b0c",x"1ce6",x"3f54",x"36eb",x"b9cd",x"3979",x"2caa",x"3b1f",x"3b0c",x"20ef",x"3f58",x"3715",x"ba65",x"38c1",x"2d9c",x"3b19",x"3b09"),
(x"9ff8",x"3f85",x"36eb",x"b3f1",x"bbbc",x"2b5c",x"3b39",x"3917",x"a2c3",x"3f85",x"36eb",x"b902",x"ba23",x"306a",x"3b3a",x"3915",x"a040",x"3f85",x"3713",x"b607",x"bb5e",x"2e4f",x"3b35",x"3914"),
(x"20f8",x"3fba",x"3716",x"38de",x"3a57",x"297d",x"3b38",x"38d2",x"210e",x"3fbb",x"36eb",x"3be3",x"2ce8",x"30c3",x"3b3c",x"38cf",x"2243",x"3fba",x"3713",x"3451",x"3bac",x"2d81",x"3b37",x"38d1"),
(x"2091",x"3f49",x"3717",x"2a07",x"3bfc",x"284d",x"3b2f",x"3b24",x"2058",x"3f49",x"36eb",x"2c56",x"3bf7",x"2bc1",x"3b35",x"3b25",x"2257",x"3f49",x"3712",x"3297",x"3bcc",x"2d84",x"3b30",x"3b23"),
(x"210b",x"3f04",x"3713",x"382e",x"baba",x"306c",x"3a31",x"3a44",x"20e4",x"3f02",x"36eb",x"366a",x"bb44",x"2f81",x"3a36",x"3a44",x"17a2",x"3f01",x"3715",x"9ef6",x"bbee",x"302a",x"3a31",x"3a40"),
(x"19fe",x"3f52",x"3717",x"2c95",x"3bf9",x"2918",x"3b19",x"3b0e",x"1a1b",x"3f52",x"36eb",x"35a6",x"3b74",x"2d53",x"3b1f",x"3b0d",x"1d4c",x"3f53",x"3717",x"b939",x"3a0b",x"29e0",x"3b19",x"3b0c"),
(x"9e8d",x"3f84",x"3716",x"bac7",x"383c",x"283f",x"3b34",x"3915",x"9efd",x"3f84",x"36eb",x"b94d",x"39f2",x"2dc5",x"3b38",x"3918",x"a040",x"3f85",x"3713",x"b607",x"bb5e",x"2e4f",x"3b35",x"3914"),
(x"1882",x"3fa8",x"370e",x"b004",x"a71d",x"3bef",x"3baa",x"3b2f",x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21",x"2273",x"3faa",x"3717",x"abf6",x"25ae",x"3bfb",x"3ba1",x"3b2f"),
(x"1f7b",x"3f4a",x"36eb",x"3b71",x"b58a",x"2fc3",x"3b35",x"3b26",x"2058",x"3f49",x"36eb",x"2c56",x"3bf7",x"2bc1",x"3b35",x"3b25",x"1f4b",x"3f49",x"3716",x"38f4",x"3a42",x"2c09",x"3b30",x"3b25"),
(x"2466",x"3f0a",x"3715",x"3ae0",x"b7cf",x"30d4",x"3a31",x"3a49",x"24bd",x"3f09",x"36eb",x"39f2",x"b938",x"30b5",x"3a36",x"3a4a",x"210b",x"3f04",x"3713",x"382e",x"baba",x"306c",x"3a31",x"3a44"),
(x"98cf",x"3f58",x"36eb",x"3976",x"39cc",x"2dcc",x"3b1f",x"3b12",x"1a1b",x"3f52",x"36eb",x"35a6",x"3b74",x"2d53",x"3b1f",x"3b0d",x"0e53",x"3f54",x"3714",x"39a7",x"399f",x"2d1e",x"3b1a",x"3b0f"),
(x"a282",x"3f82",x"36eb",x"b9ec",x"392b",x"31e4",x"3b37",x"391b",x"9efd",x"3f84",x"36eb",x"b94d",x"39f2",x"2dc5",x"3b38",x"3918",x"a17b",x"3f81",x"3711",x"b8c8",x"3a4e",x"30a8",x"3b33",x"3917"),
(x"1f7b",x"3f4a",x"36eb",x"3b71",x"b58a",x"2fc3",x"3b35",x"3b26",x"1f4b",x"3f49",x"3716",x"38f4",x"3a42",x"2c09",x"3b30",x"3b25",x"1e77",x"3f4b",x"3715",x"3ac2",x"b812",x"3146",x"3b30",x"3b26"),
(x"253f",x"3f13",x"3715",x"3bec",x"abe2",x"2fce",x"3a30",x"3a4e",x"2585",x"3f12",x"36eb",x"3bc4",x"b27a",x"3012",x"3a35",x"3a4f",x"2466",x"3f0a",x"3715",x"3ae0",x"b7cf",x"30d4",x"3a31",x"3a49"),
(x"9e13",x"3f5b",x"36eb",x"353f",x"3b87",x"2d28",x"3b20",x"3b14",x"98cf",x"3f58",x"36eb",x"3976",x"39cc",x"2dcc",x"3b1f",x"3b12",x"9e62",x"3f5a",x"3716",x"37d5",x"3af0",x"2d8e",x"3b1a",x"3b14"),
(x"a471",x"3f79",x"36eb",x"bbbc",x"3212",x"3175",x"3b34",x"391f",x"a282",x"3f82",x"36eb",x"b9ec",x"392b",x"31e4",x"3b37",x"391b",x"a407",x"3f79",x"370f",x"bb4b",x"35cc",x"3223",x"3b30",x"391b"),
(x"21ae",x"3fcd",x"36eb",x"3ade",x"37ab",x"31d3",x"3b41",x"38d7",x"229f",x"3fc1",x"36eb",x"3bdb",x"1c67",x"320a",x"3b3e",x"38d2",x"20f7",x"3fcc",x"370e",x"3b7b",x"34a9",x"3270",x"3b3d",x"38d9"),
(x"22bc",x"3f52",x"36eb",x"3adb",x"b7e7",x"30ac",x"3b35",x"3b2b",x"1e77",x"3f4b",x"3715",x"3ac2",x"b812",x"3146",x"3b30",x"3b26",x"2147",x"3f51",x"3718",x"3ac6",x"b7dc",x"3286",x"3b2f",x"3b2a"),
(x"24fc",x"3f1b",x"3717",x"3b55",x"35fd",x"307e",x"3a2f",x"3a53",x"255d",x"3f1c",x"36eb",x"3b6e",x"3575",x"309e",x"3a34",x"3a54",x"253f",x"3f13",x"3715",x"3bec",x"abe2",x"2fce",x"3a30",x"3a4e"),
(x"a16d",x"3f34",x"3711",x"b115",x"27d5",x"3be4",x"3bb6",x"3b90",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f",x"9c3a",x"3f30",x"3714",x"b05e",x"21a1",x"3bec",x"3bb1",x"3b94"),
(x"a172",x"3f5c",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"3b20",x"3b17",x"9e13",x"3f5b",x"36eb",x"353f",x"3b87",x"2d28",x"3b20",x"3b14",x"a13d",x"3f5b",x"3716",x"a345",x"3bf7",x"2dcc",x"3b1a",x"3b17"),
(x"a482",x"3f6f",x"36eb",x"bb61",x"b5a0",x"3119",x"3b30",x"3922",x"a471",x"3f79",x"36eb",x"bbbc",x"3212",x"3175",x"3b34",x"391f",x"a425",x"3f70",x"370f",x"bbd3",x"af46",x"3182",x"3b2d",x"391f"),
(x"2496",x"3f5d",x"36eb",x"3bba",x"b376",x"2f14",x"3b35",x"3b31",x"22bc",x"3f52",x"36eb",x"3adb",x"b7e7",x"30ac",x"3b35",x"3b2b",x"2442",x"3f5d",x"3714",x"3b6b",x"b587",x"3095",x"3b30",x"3b31"),
(x"2409",x"3f24",x"36eb",x"3884",x"3a69",x"324a",x"3a33",x"3a59",x"255d",x"3f1c",x"36eb",x"3b6e",x"3575",x"309e",x"3a34",x"3a54",x"2375",x"3f22",x"3711",x"38a4",x"3a69",x"309a",x"3a2f",x"3a57"),
(x"a38b",x"3f5a",x"36eb",x"bacc",x"3812",x"3065",x"3b20",x"3b19",x"a172",x"3f5c",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"3b20",x"3b17",x"a2d9",x"3f59",x"3714",x"b976",x"39c0",x"3024",x"3b1b",x"3b19"),
(x"a2ad",x"3f6a",x"36eb",x"b86e",x"ba87",x"313e",x"3b2e",x"3925",x"a482",x"3f6f",x"36eb",x"bb61",x"b5a0",x"3119",x"3b30",x"3922",x"a289",x"3f6b",x"370f",x"b891",x"ba72",x"30f5",x"3b2b",x"3921"),
(x"1a0c",x"3fd7",x"36eb",x"38a6",x"3a54",x"3207",x"3b44",x"38de",x"21ae",x"3fcd",x"36eb",x"3ade",x"37ab",x"31d3",x"3b41",x"38d7",x"1aac",x"3fd4",x"3712",x"38b5",x"3a3e",x"32bd",x"3b3f",x"38df"),
(x"250f",x"3f6a",x"36eb",x"3bef",x"2d0b",x"2e69",x"3b35",x"3b38",x"2496",x"3f5d",x"36eb",x"3bba",x"b376",x"2f14",x"3b35",x"3b31",x"24cc",x"3f69",x"3712",x"3bf0",x"aa00",x"2f46",x"3b31",x"3b38"),
(x"1f0f",x"3f25",x"3718",x"38ae",x"3a78",x"2b7c",x"3a2c",x"3a5b",x"1fad",x"3f26",x"36eb",x"360d",x"3b5a",x"2ef4",x"3a31",x"3a5d",x"2375",x"3f22",x"3711",x"38a4",x"3a69",x"309a",x"3a2f",x"3a57"),
(x"a422",x"3f54",x"36eb",x"bbcf",x"b174",x"303e",x"3b1f",x"3b1c",x"a38b",x"3f5a",x"36eb",x"bacc",x"3812",x"3065",x"3b20",x"3b19",x"a38f",x"3f55",x"3712",x"bbe0",x"2e5e",x"30a3",x"3b1b",x"3b1b"),
(x"a035",x"3f6a",x"3713",x"3583",x"bb63",x"3153",x"3b29",x"3922",x"9f83",x"3f68",x"36eb",x"35e4",x"bb4d",x"31a2",x"3b2b",x"3927",x"a289",x"3f6b",x"370f",x"b891",x"ba72",x"30f5",x"3b2b",x"3921"),
(x"91f4",x"3fd4",x"3716",x"badd",x"375a",x"334d",x"3b3f",x"38e1",x"980d",x"3fd7",x"36eb",x"b996",x"395e",x"33ec",x"3b44",x"38e0",x"1aac",x"3fd4",x"3712",x"38b5",x"3a3e",x"32bd",x"3b3f",x"38df"),
(x"2469",x"3f76",x"36eb",x"3b75",x"35a2",x"2d46",x"3b35",x"3b3e",x"250f",x"3f6a",x"36eb",x"3bef",x"2d0b",x"2e69",x"3b35",x"3b38",x"243c",x"3f75",x"3710",x"3b6a",x"35bb",x"2efe",x"3b31",x"3b3e"),
(x"1d9c",x"3f28",x"3718",x"3be6",x"309e",x"2baa",x"3a2c",x"3a5c",x"1e52",x"3f28",x"36eb",x"3be6",x"308f",x"2c41",x"3a31",x"3a5e",x"1f0f",x"3f25",x"3718",x"38ae",x"3a78",x"2b7c",x"3a2c",x"3a5b"),
(x"a30f",x"3f4f",x"36eb",x"b6fe",x"bb25",x"2ea4",x"3b1f",x"3b1f",x"a422",x"3f54",x"36eb",x"bbcf",x"b174",x"303e",x"3b1f",x"3b1c",x"a2cb",x"3f51",x"3714",x"b972",x"b9bb",x"30de",x"3b1a",x"3b1d"),
(x"a175",x"3f1a",x"3710",x"2828",x"260a",x"3bfe",x"3bb7",x"3ba6",x"a140",x"3f12",x"3714",x"2946",x"1ffc",x"3bfe",x"3bb7",x"3bac",x"a2ee",x"3f13",x"3714",x"2eb0",x"28fa",x"3bf3",x"3bb9",x"3bab"),
(x"a099",x"3f0e",x"3712",x"2953",x"27ae",x"3bfd",x"3bb6",x"3bb0",x"9ecc",x"3f0b",x"3714",x"a8bf",x"2c22",x"3bfa",x"3bb4",x"3bb3",x"a1ea",x"3f0b",x"3712",x"a587",x"208e",x"3bff",x"3bb8",x"3bb2"),
(x"9aa8",x"3f08",x"3714",x"231d",x"2b5f",x"3bfc",x"3bb2",x"3bb5",x"9d7f",x"3f04",x"3715",x"a0ea",x"2b00",x"3bfc",x"3bb3",x"3bb9",x"9ecc",x"3f0b",x"3714",x"a8bf",x"2c22",x"3bfa",x"3bb4",x"3bb3"),
(x"1a1e",x"3f06",x"3715",x"270a",x"a779",x"3bfe",x"3bad",x"3bb7",x"17a2",x"3f01",x"3715",x"27e2",x"29b5",x"3bfc",x"3bae",x"3bbb",x"9aa8",x"3f08",x"3714",x"231d",x"2b5f",x"3bfc",x"3bb2",x"3bb5"),
(x"20b2",x"3f08",x"3716",x"24bc",x"aceb",x"3bf9",x"3ba8",x"3bb6",x"210b",x"3f04",x"3713",x"2b1d",x"aee4",x"3bf0",x"3ba7",x"3bb9",x"1a1e",x"3f06",x"3715",x"270a",x"a779",x"3bfe",x"3bad",x"3bb7"),
(x"2335",x"3f0e",x"3714",x"a8e0",x"299e",x"3bfc",x"3ba4",x"3bb1",x"2466",x"3f0a",x"3715",x"a266",x"9d87",x"3bff",x"3ba1",x"3bb4",x"20b2",x"3f08",x"3716",x"24bc",x"aceb",x"3bf9",x"3ba8",x"3bb6"),
(x"23d3",x"3f13",x"3714",x"a538",x"a9ab",x"3bfd",x"3ba3",x"3bad",x"253f",x"3f13",x"3715",x"a891",x"a7ce",x"3bfd",x"3b9e",x"3bad",x"2335",x"3f0e",x"3714",x"a8e0",x"299e",x"3bfc",x"3ba4",x"3bb1"),
(x"23d3",x"3f13",x"3714",x"a538",x"a9ab",x"3bfd",x"3ba3",x"3bad",x"22d3",x"3f18",x"3715",x"ac67",x"28a5",x"3bf9",x"3ba4",x"3ba9",x"253f",x"3f13",x"3715",x"a891",x"a7ce",x"3bfd",x"3b9e",x"3bad"),
(x"20d5",x"3f18",x"3714",x"aa45",x"2b10",x"3bfa",x"3ba7",x"3ba8",x"2375",x"3f22",x"3711",x"a8d9",x"a52b",x"3bfe",x"3ba2",x"3ba0",x"22d3",x"3f18",x"3715",x"ac67",x"28a5",x"3bf9",x"3ba4",x"3ba9"),
(x"14bb",x"3f16",x"3710",x"a352",x"ae80",x"3bf5",x"3bae",x"3baa",x"951c",x"3f19",x"3711",x"abef",x"a8a8",x"3bfa",x"3baf",x"3ba7",x"1e4f",x"3f16",x"3711",x"aa66",x"b31a",x"3bca",x"3baa",x"3baa"),
(x"1d9c",x"3f28",x"3718",x"b420",x"1418",x"3bba",x"3ba9",x"3b9b",x"1f0f",x"3f25",x"3718",x"ab65",x"b528",x"3b8f",x"3ba8",x"3b9d",x"15a0",x"3f25",x"3713",x"b41f",x"ac3a",x"3bb6",x"3bad",x"3b9d"),
(x"16c6",x"3f29",x"3714",x"ade0",x"a4c2",x"3bf6",x"3bad",x"3b99",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f",x"1d4f",x"3f31",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3baa",x"3b93"),
(x"951c",x"3f19",x"3711",x"abef",x"a8a8",x"3bfa",x"3baf",x"3ba7",x"983c",x"3f20",x"3710",x"a856",x"a9ab",x"3bfc",x"3bb0",x"3ba1",x"20d5",x"3f18",x"3714",x"aa45",x"2b10",x"3bfa",x"3ba7",x"3ba8"),
(x"a3f1",x"3ec4",x"3718",x"a6a1",x"97c8",x"3bff",x"3981",x"31ad",x"a1bd",x"3ee0",x"3715",x"a1a1",x"23fc",x"3bff",x"3983",x"31eb",x"a069",x"3ec3",x"3718",x"a24c",x"a379",x"3bff",x"3985",x"31ab"),
(x"1e3f",x"3f34",x"3715",x"28bf",x"afdb",x"3bef",x"3ba9",x"3b91",x"1d4f",x"3f31",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3baa",x"3b93",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f"),
(x"13e1",x"3f25",x"36eb",x"bbf6",x"2a70",x"2d61",x"3a69",x"3a31",x"8dee",x"3f36",x"36eb",x"b469",x"bb91",x"316a",x"3a68",x"3a28",x"16c6",x"3f29",x"3714",x"bbf3",x"ae23",x"2b27",x"3a63",x"3a30"),
(x"20de",x"3dea",x"3715",x"ad56",x"a0d0",x"3bf8",x"3b6f",x"3b0e",x"1c89",x"3ddc",x"3716",x"b0f9",x"28af",x"3be5",x"3b6a",x"3b03",x"9e24",x"3de5",x"370e",x"afd2",x"a717",x"3bef",x"3b62",x"3b0b"),
(x"20de",x"3dea",x"3715",x"3bc5",x"ab9a",x"3358",x"3b8c",x"3a3c",x"2222",x"3de9",x"36eb",x"3b99",x"b315",x"330d",x"3b91",x"3a3c",x"1c89",x"3ddc",x"3716",x"3add",x"b75a",x"334d",x"3b8c",x"3a34"),
(x"1f0d",x"3e22",x"3713",x"2da3",x"af14",x"3beb",x"3b70",x"3b3f",x"1ba5",x"3e29",x"3714",x"2c39",x"a9a5",x"3bf9",x"3b6e",x"3b46",x"2079",x"3e21",x"3712",x"2a69",x"a87e",x"3bfc",x"3b72",x"3b3e"),
(x"242c",x"3e29",x"3712",x"2a73",x"aa97",x"3bfa",x"3b78",x"3b45",x"2498",x"3e24",x"3711",x"2481",x"a546",x"3bff",x"3b7a",x"3b40",x"21e0",x"3e1f",x"3711",x"2994",x"a977",x"3bfc",x"3b74",x"3b3d"),
(x"21e0",x"3e1f",x"3711",x"2994",x"a977",x"3bfc",x"3b74",x"3b3d",x"2079",x"3e21",x"3712",x"2a69",x"a87e",x"3bfc",x"3b72",x"3b3e",x"242c",x"3e29",x"3712",x"2a73",x"aa97",x"3bfa",x"3b78",x"3b45"),
(x"212c",x"3e2d",x"3716",x"2f15",x"b29c",x"3bc6",x"3b73",x"3b48",x"2000",x"3e2e",x"3718",x"2e36",x"2160",x"3bf6",x"3b72",x"3b49",x"2360",x"3e2f",x"3711",x"2fec",x"2c2c",x"3beb",x"3b77",x"3b4a"),
(x"1fdf",x"3e42",x"370f",x"ab8a",x"b0ae",x"3be6",x"3b73",x"3b5b",x"221a",x"3e47",x"3713",x"2e9c",x"b366",x"3bbd",x"3b76",x"3b5f",x"2010",x"3e3f",x"370e",x"a6d5",x"a5c2",x"3bfe",x"3b73",x"3b59"),
(x"2517",x"3e40",x"370f",x"2cd8",x"271d",x"3bf9",x"3b7d",x"3b59",x"219e",x"3e3b",x"3713",x"2538",x"2c79",x"3bfa",x"3b75",x"3b54",x"2437",x"3e45",x"370f",x"1df0",x"2631",x"3bff",x"3b7a",x"3b5d"),
(x"2517",x"3e40",x"370f",x"2cd8",x"271d",x"3bf9",x"3b7d",x"3b59",x"24fa",x"3e37",x"370f",x"2ec5",x"9a24",x"3bf4",x"3b7c",x"3b51",x"219e",x"3e3b",x"3713",x"2538",x"2c79",x"3bfa",x"3b75",x"3b54"),
(x"2360",x"3e2f",x"3711",x"2fec",x"2c2c",x"3beb",x"3b77",x"3b4a",x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d",x"2072",x"3e36",x"3710",x"2c5b",x"30a5",x"3be5",x"3b73",x"3b51"),
(x"9607",x"3e5d",x"3717",x"17c8",x"1f79",x"3c00",x"3b6a",x"3b72",x"9959",x"3e66",x"3715",x"26c2",x"2c63",x"3bfa",x"3b6a",x"3b7a",x"125b",x"3e5e",x"3717",x"2ff2",x"2a7d",x"3bed",x"3b6c",x"3b73"),
(x"2458",x"3e5f",x"3714",x"9553",x"2b62",x"3bfc",x"3b79",x"3b74",x"24ba",x"3e5b",x"3712",x"3163",x"2345",x"3be2",x"3b7b",x"3b71",x"2323",x"3e55",x"3716",x"2cd8",x"27e2",x"3bf9",x"3b77",x"3b6c"),
(x"2323",x"3e55",x"3716",x"2cd8",x"27e2",x"3bf9",x"3b77",x"3b6c",x"2116",x"3e56",x"3716",x"a818",x"2d04",x"3bf8",x"3b74",x"3b6c",x"2458",x"3e5f",x"3714",x"9553",x"2b62",x"3bfc",x"3b79",x"3b74"),
(x"1e07",x"3e59",x"3714",x"2504",x"2da9",x"3bf7",x"3b70",x"3b6f",x"2074",x"3e62",x"3711",x"a40b",x"2d5c",x"3bf8",x"3b73",x"3b77",x"2116",x"3e56",x"3716",x"a818",x"2d04",x"3bf8",x"3b74",x"3b6c"),
(x"1acb",x"3e5c",x"3714",x"3036",x"273e",x"3bed",x"3b6e",x"3b72",x"125b",x"3e5e",x"3717",x"2ff2",x"2a7d",x"3bed",x"3b6c",x"3b73",x"1f03",x"3e64",x"3711",x"327d",x"975f",x"3bd5",x"3b71",x"3b78"),
(x"2353",x"3e7c",x"3711",x"3115",x"a7d5",x"3be4",x"3b78",x"3b8d",x"1f3f",x"3e6b",x"3712",x"3146",x"ac91",x"3bde",x"3b71",x"3b7e",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c"),
(x"98e9",x"3e7d",x"3715",x"a8bf",x"2fdb",x"3bef",x"3b6a",x"3b8d",x"9aa8",x"3e77",x"3718",x"a138",x"2e95",x"3bf4",x"3b69",x"3b89",x"9ff6",x"3e78",x"3719",x"290e",x"2f00",x"3bf2",x"3b66",x"3b89"),
(x"98e9",x"3e7d",x"3715",x"a8bf",x"2fdb",x"3bef",x"3b6a",x"3b8d",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c",x"9aa8",x"3e77",x"3718",x"a138",x"2e95",x"3bf4",x"3b69",x"3b89"),
(x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"9920",x"3e76",x"3718",x"ab4f",x"a525",x"3bfc",x"3b6a",x"3b88",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c"),
(x"9dca",x"3e73",x"3715",x"ad65",x"2c5a",x"3bf3",x"3b67",x"3b85",x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"a0a3",x"3e6e",x"3718",x"acf2",x"991e",x"3bf9",x"3b64",x"3b81"),
(x"a072",x"3e68",x"3712",x"b542",x"b0b9",x"3b76",x"3b64",x"3b7b",x"a0f6",x"3e69",x"3712",x"b59c",x"b36a",x"3b42",x"3b64",x"3b7d",x"9d58",x"3e68",x"3717",x"ad2d",x"aecb",x"3bed",x"3b67",x"3b7c"),
(x"9d58",x"3e68",x"3717",x"ad2d",x"aecb",x"3bed",x"3b67",x"3b7c",x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"9b02",x"3e67",x"3716",x"3009",x"ada6",x"3be7",x"3b69",x"3b7b"),
(x"9959",x"3e66",x"3715",x"26c2",x"2c63",x"3bfa",x"3b6a",x"3b7a",x"9b02",x"3e67",x"3716",x"3009",x"ada6",x"3be7",x"3b69",x"3b7b",x"1e50",x"3e66",x"3712",x"2f67",x"2981",x"3bf0",x"3b71",x"3b7a"),
(x"9abe",x"3e63",x"3714",x"257a",x"2e8a",x"3bf4",x"3b69",x"3b78",x"9959",x"3e66",x"3715",x"26c2",x"2c63",x"3bfa",x"3b6a",x"3b7a",x"9607",x"3e5d",x"3717",x"17c8",x"1f79",x"3c00",x"3b6a",x"3b72"),
(x"9ec5",x"3e5f",x"3718",x"2c00",x"a90e",x"3bfa",x"3b66",x"3b75",x"9e13",x"3e58",x"3715",x"251e",x"ad06",x"3bf9",x"3b67",x"3b6e",x"a29f",x"3e53",x"3714",x"975f",x"ac2c",x"3bfb",x"3b61",x"3b6a"),
(x"a29f",x"3e53",x"3714",x"975f",x"ac2c",x"3bfb",x"3b61",x"3b6a",x"a123",x"3e50",x"3714",x"adba",x"a266",x"3bf7",x"3b63",x"3b68",x"a3b3",x"3e47",x"3712",x"b106",x"a73e",x"3be5",x"3b5f",x"3b60"),
(x"a3b3",x"3e47",x"3712",x"b106",x"a73e",x"3be5",x"3b5f",x"3b60",x"a180",x"3e45",x"3715",x"b468",x"a47a",x"3bb0",x"3b63",x"3b5e",x"a294",x"3e3b",x"3710",x"b550",x"ae33",x"3b81",x"3b61",x"3b55"),
(x"a294",x"3e3b",x"3710",x"b550",x"ae33",x"3b81",x"3b61",x"3b55",x"a0d7",x"3e3d",x"3717",x"b273",x"af43",x"3bc8",x"3b64",x"3b57",x"9faa",x"3e33",x"3712",x"ab5c",x"a345",x"3bfc",x"3b65",x"3b4f"),
(x"9faa",x"3e33",x"3712",x"ab5c",x"a345",x"3bfc",x"3b65",x"3b4f",x"9ad5",x"3e36",x"3711",x"2e24",x"aa2b",x"3bf4",x"3b69",x"3b51",x"11f0",x"3e35",x"3712",x"add2",x"304b",x"3be4",x"3b6c",x"3b50"),
(x"1d2c",x"3e2c",x"3716",x"2553",x"b2c7",x"3bd1",x"3b6f",x"3b48",x"1b46",x"3e2e",x"3716",x"af4b",x"2a5f",x"3bf0",x"3b6e",x"3b49",x"2000",x"3e2e",x"3718",x"2e36",x"2160",x"3bf6",x"3b72",x"3b49"),
(x"1d2c",x"3e2c",x"3716",x"2553",x"b2c7",x"3bd1",x"3b6f",x"3b48",x"2000",x"3e2e",x"3718",x"2e36",x"2160",x"3bf6",x"3b72",x"3b49",x"212c",x"3e2d",x"3716",x"2f15",x"b29c",x"3bc6",x"3b73",x"3b48"),
(x"1ba5",x"3e29",x"3714",x"2c39",x"a9a5",x"3bf9",x"3b6e",x"3b46",x"1f0d",x"3e22",x"3713",x"2da3",x"af14",x"3beb",x"3b70",x"3b3f",x"9aec",x"3e22",x"3717",x"30e7",x"b057",x"3bd4",x"3b68",x"3b3f"),
(x"9aec",x"3e22",x"3717",x"30e7",x"b057",x"3bd4",x"3b68",x"3b3f",x"16e7",x"3e1d",x"370f",x"2edc",x"acd0",x"3bee",x"3b6c",x"3b3b",x"a039",x"3e14",x"3713",x"29b8",x"26e9",x"3bfd",x"3b64",x"3b34"),
(x"a039",x"3e14",x"3713",x"29b8",x"26e9",x"3bfd",x"3b64",x"3b34",x"9631",x"3e13",x"3716",x"2adf",x"26b5",x"3bfc",x"3b69",x"3b32",x"a08e",x"3e07",x"3717",x"2bf6",x"a5ae",x"3bfb",x"3b62",x"3b29"),
(x"a08e",x"3e07",x"3717",x"2bf6",x"a5ae",x"3bfb",x"3b62",x"3b29",x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a",x"a1a0",x"3dfc",x"370f",x"b6ca",x"afac",x"3b2e",x"3b5f",x"3b1f"),
(x"a05e",x"3df6",x"3713",x"af9f",x"3907",x"3a25",x"3b61",x"3b1a",x"a12d",x"3df8",x"370d",x"b809",x"ae09",x"3add",x"3b5f",x"3b1c",x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a"),
(x"9e24",x"3de5",x"370e",x"afd2",x"a717",x"3bef",x"3b62",x"3b0b",x"9f80",x"3def",x"3712",x"a9f0",x"ab1d",x"3bfa",x"3b61",x"3b14",x"20de",x"3dea",x"3715",x"ad56",x"a0d0",x"3bf8",x"3b6f",x"3b0e"),
(x"2043",x"3df7",x"3715",x"3b81",x"3440",x"330f",x"3b8b",x"3a42",x"1624",x"3e08",x"370e",x"3b5f",x"35f1",x"2f4d",x"3b89",x"3a4c",x"2166",x"3df7",x"36eb",x"3b89",x"3473",x"31fc",x"3b90",x"3a43"),
(x"2307",x"3e8d",x"36eb",x"bba1",x"34cc",x"1f45",x"3b3d",x"3b5a",x"234d",x"3e9c",x"36eb",x"bbf5",x"ae59",x"2467",x"3b3d",x"3b53",x"235a",x"3e97",x"3710",x"bbfd",x"2997",x"a0a8",x"3b38",x"3b56"),
(x"1c29",x"3e7b",x"36eb",x"346a",x"3b91",x"316a",x"3b3c",x"3b66",x"2307",x"3e8d",x"36eb",x"bba1",x"34cc",x"1f45",x"3b3d",x"3b5a",x"2002",x"3e80",x"3714",x"bb1c",x"3754",x"223f",x"3b37",x"3b62"),
(x"234d",x"3e9c",x"36eb",x"bbf5",x"ae59",x"2467",x"3b3d",x"3b53",x"2237",x"3ea4",x"36eb",x"bab1",x"b862",x"21f0",x"3b3d",x"3b4f",x"227e",x"3ea3",x"3712",x"bb76",x"b5c5",x"204d",x"3b38",x"3b4f"),
(x"2237",x"3ea4",x"36eb",x"bab1",x"b862",x"21f0",x"3b3d",x"3b4f",x"1f6a",x"3ea8",x"36eb",x"b7e1",x"baf5",x"269a",x"3b3d",x"3b4b",x"214b",x"3ea6",x"3714",x"b95a",x"b9f1",x"2025",x"3b38",x"3b4d"),
(x"1f6a",x"3ea8",x"36eb",x"b7e1",x"baf5",x"269a",x"3b3d",x"3b4b",x"142d",x"3eaa",x"36eb",x"b03c",x"bbeb",x"299b",x"3b3d",x"3b48",x"1f1f",x"3ea8",x"3714",x"b5bf",x"bb76",x"27db",x"3b38",x"3b4b"),
(x"142d",x"3eaa",x"36eb",x"b03c",x"bbeb",x"299b",x"3b3d",x"3b48",x"9d76",x"3ea9",x"36eb",x"3868",x"baab",x"296a",x"3b3d",x"3b44",x"11db",x"3eaa",x"3715",x"2836",x"bbfd",x"294f",x"3b38",x"3b47"),
(x"9d99",x"3ea9",x"3716",x"386f",x"baa7",x"2604",x"3b38",x"3b44",x"9d76",x"3ea9",x"36eb",x"3868",x"baab",x"296a",x"3b3d",x"3b44",x"a14f",x"3ea3",x"3714",x"3b01",x"b7b5",x"2839",x"3b39",x"3b40"),
(x"a11a",x"3ea2",x"36eb",x"3af3",x"b7df",x"2b38",x"3b3e",x"3b40",x"a1ea",x"3e9d",x"36eb",x"3bf9",x"ad11",x"2511",x"3b3e",x"3b3d",x"a14f",x"3ea3",x"3714",x"3b01",x"b7b5",x"2839",x"3b39",x"3b40"),
(x"a1ea",x"3e9d",x"36eb",x"3bf9",x"ad11",x"2511",x"3b3e",x"3b3d",x"a11a",x"3e99",x"36eb",x"390c",x"3a34",x"2532",x"3b3e",x"3b3b",x"a1ee",x"3e9d",x"3714",x"3be6",x"310f",x"9bfc",x"3b39",x"3b3d"),
(x"a0ed",x"3e98",x"3715",x"3928",x"3a1d",x"1553",x"3b39",x"3b3a",x"a11a",x"3e99",x"36eb",x"390c",x"3a34",x"2532",x"3b3e",x"3b3b",x"9ddf",x"3e98",x"3714",x"afe4",x"3bee",x"28fd",x"3b39",x"3b38"),
(x"9ddf",x"3e98",x"3714",x"afe4",x"3bee",x"28fd",x"3b39",x"3b38",x"9d99",x"3e98",x"36eb",x"b5dd",x"3b6d",x"2be9",x"3b3e",x"3b38",x"9908",x"3e9a",x"3711",x"b64f",x"3b52",x"2d1b",x"3b3a",x"3b36"),
(x"1bc8",x"3e8d",x"36eb",x"39db",x"b96c",x"2c1a",x"3b3e",x"3b2b",x"199d",x"3e8c",x"36eb",x"3bf6",x"aa70",x"2d61",x"3b3e",x"3b29",x"1b8a",x"3e8e",x"3711",x"3a7a",x"b8af",x"2839",x"3b39",x"3b2c"),
(x"9908",x"3e9a",x"3711",x"b64f",x"3b52",x"2d1b",x"3b3a",x"3b36",x"99c6",x"3e9b",x"36eb",x"b2b1",x"3bc8",x"2e54",x"3b3f",x"3b37",x"1937",x"3e9a",x"3710",x"3416",x"3bad",x"2f8d",x"3b3a",x"3b33"),
(x"1e92",x"3e42",x"36eb",x"bb7d",x"3521",x"3096",x"3b1d",x"3b54",x"21a6",x"3e48",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b1f",x"3b51",x"1fdf",x"3e42",x"370f",x"ba9b",x"3854",x"30fa",x"3b19",x"3b52"),
(x"2043",x"3df7",x"3715",x"3b81",x"3440",x"330f",x"3b8b",x"3a42",x"2166",x"3df7",x"36eb",x"3b89",x"3473",x"31fc",x"3b90",x"3a43",x"20de",x"3dea",x"3715",x"3bc5",x"ab9a",x"3358",x"3b8c",x"3a3c"),
(x"a18f",x"3e8e",x"3711",x"28d9",x"252b",x"3bfe",x"3b63",x"3b9d",x"1de8",x"3e90",x"3710",x"2856",x"29ab",x"3bfc",x"3b71",x"3b9e",x"9a89",x"3e8b",x"3718",x"2b65",x"3528",x"3b8f",x"3b69",x"3b9a"),
(x"9e52",x"3df5",x"36eb",x"bbe3",x"ace8",x"30c3",x"3b8a",x"3a22",x"9e25",x"3df6",x"3716",x"b8de",x"ba57",x"297d",x"3b86",x"3a25",x"9de0",x"3df4",x"3715",x"bbd7",x"31f9",x"2c2a",x"3b86",x"3a26"),
(x"9faa",x"3e33",x"3712",x"b84e",x"bab0",x"2ec8",x"3a3a",x"3a41",x"a081",x"3e33",x"36eb",x"b958",x"b9de",x"2fdf",x"3a3f",x"3a41",x"a294",x"3e3b",x"3710",x"bb6a",x"b5bb",x"2efe",x"3a3b",x"3a3c"),
(x"1ab2",x"3e9b",x"36eb",x"337e",x"3bba",x"2ef6",x"3b3f",x"3b33",x"1e0f",x"3e99",x"36eb",x"3aa4",x"3859",x"2fe4",x"3b3f",x"3b31",x"1937",x"3e9a",x"3710",x"3416",x"3bad",x"2f8d",x"3b3a",x"3b33"),
(x"989a",x"3e7f",x"36eb",x"bbfa",x"20b5",x"2cb4",x"3b37",x"38b1",x"990f",x"3e89",x"36eb",x"bbe6",x"b08f",x"2c41",x"3b3a",x"38ac",x"9613",x"3e7f",x"3715",x"bbfa",x"2710",x"2c48",x"3b33",x"38ae"),
(x"1d11",x"3e98",x"3711",x"3a7e",x"3887",x"3089",x"3b3a",x"3b31",x"1e0f",x"3e99",x"36eb",x"3aa4",x"3859",x"2fe4",x"3b3f",x"3b31",x"1ea1",x"3e94",x"3710",x"3bcc",x"3228",x"2f2f",x"3b3a",x"3b30"),
(x"1f2f",x"3e3f",x"36eb",x"bb19",x"b744",x"2cf7",x"3b1c",x"3b55",x"1e92",x"3e42",x"36eb",x"bb7d",x"3521",x"3096",x"3b1d",x"3b54",x"2010",x"3e3f",x"370e",x"bb25",x"b70d",x"2d6a",x"3b19",x"3b53"),
(x"201d",x"3e63",x"36eb",x"37d8",x"3af6",x"2a35",x"3b42",x"3861",x"247a",x"3e61",x"36eb",x"36fe",x"3b25",x"2ea4",x"3b42",x"385c",x"2074",x"3e62",x"3711",x"34dc",x"3b97",x"2d61",x"3b3e",x"3861"),
(x"1edf",x"3e90",x"36eb",x"3b02",x"b776",x"2fc8",x"3b3e",x"3b2c",x"1bc8",x"3e8d",x"36eb",x"39db",x"b96c",x"2c1a",x"3b3e",x"3b2b",x"1de8",x"3e90",x"3710",x"3b2f",x"b6d9",x"2e52",x"3b3a",x"3b2d"),
(x"1b46",x"3e2e",x"3716",x"b7e9",x"baf1",x"2aa7",x"3a3a",x"3a48",x"1c1b",x"3e2d",x"36eb",x"b776",x"bb0b",x"2d41",x"3a3f",x"3a49",x"9faa",x"3e33",x"3712",x"b84e",x"bab0",x"2ec8",x"3a3a",x"3a41"),
(x"98e9",x"3e7d",x"3715",x"b95d",x"39e3",x"2de3",x"3b32",x"38af",x"9943",x"3e7e",x"36eb",x"b9df",x"3964",x"2d28",x"3b37",x"38b2",x"9613",x"3e7f",x"3715",x"bbfa",x"2710",x"2c48",x"3b33",x"38ae"),
(x"219e",x"3e3b",x"3713",x"bb5b",x"b634",x"2c03",x"3b17",x"3b55",x"2166",x"3e3a",x"36eb",x"bad3",x"b822",x"2c4d",x"3b1b",x"3b58",x"2010",x"3e3f",x"370e",x"bb25",x"b70d",x"2d6a",x"3b19",x"3b53"),
(x"9631",x"3e13",x"3716",x"3bff",x"a0c2",x"2138",x"3b87",x"3a51",x"95be",x"3e13",x"36eb",x"3bfe",x"9ea7",x"2828",x"3b8c",x"3a53",x"1624",x"3e08",x"370e",x"3b5f",x"35f1",x"2f4d",x"3b89",x"3a4c"),
(x"1cd4",x"3e2c",x"36eb",x"bb24",x"371c",x"2cde",x"3a3f",x"3a49",x"1c1b",x"3e2d",x"36eb",x"b776",x"bb0b",x"2d41",x"3a3f",x"3a49",x"1d2c",x"3e2c",x"3716",x"bbde",x"b1b6",x"2825",x"3a3a",x"3a49"),
(x"9ff6",x"3e78",x"3719",x"b9a6",x"3994",x"2fc6",x"3b30",x"38b3",x"a0ef",x"3e78",x"36eb",x"b9ed",x"394b",x"2f45",x"3b35",x"38b6",x"98e9",x"3e7d",x"3715",x"b95d",x"39e3",x"2de3",x"3b32",x"38af"),
(x"1f30",x"3e66",x"36eb",x"3bf8",x"2379",x"2d44",x"3b43",x"3863",x"201d",x"3e63",x"36eb",x"37d8",x"3af6",x"2a35",x"3b42",x"3861",x"1f03",x"3e64",x"3711",x"3b12",x"3763",x"2ca3",x"3b3e",x"3862"),
(x"21a8",x"3e39",x"3713",x"bb09",x"3791",x"2ab8",x"3b2f",x"382f",x"216e",x"3e39",x"36eb",x"b9e9",x"3955",x"2e31",x"3b34",x"382e",x"219e",x"3e3b",x"3713",x"bb5b",x"b634",x"2c03",x"3b2f",x"382e"),
(x"17ea",x"3e1d",x"36eb",x"3ab4",x"b859",x"2a66",x"3b8b",x"3a58",x"95be",x"3e13",x"36eb",x"3bfe",x"9ea7",x"2828",x"3b8c",x"3a53",x"16e7",x"3e1d",x"370f",x"3ad7",x"b821",x"29e6",x"3b87",x"3a57"),
(x"1986",x"3e2a",x"36eb",x"b97a",x"39b6",x"309a",x"3a3f",x"3a4b",x"1cd4",x"3e2c",x"36eb",x"bb24",x"371c",x"2cde",x"3a3f",x"3a49",x"1ba5",x"3e29",x"3714",x"b9e8",x"3951",x"2f27",x"3a3a",x"3a4a"),
(x"a09e",x"3e76",x"36eb",x"b2cb",x"bbc1",x"2fc5",x"3b35",x"38b7",x"a0ef",x"3e78",x"36eb",x"b9ed",x"394b",x"2f45",x"3b35",x"38b6",x"9fe7",x"3e77",x"3719",x"b250",x"bbca",x"2f22",x"3b30",x"38b3"),
(x"1fbf",x"3e6a",x"36eb",x"3b57",x"b625",x"2e99",x"3b43",x"3865",x"1f30",x"3e66",x"36eb",x"3bf8",x"2379",x"2d44",x"3b43",x"3863",x"1f3f",x"3e6b",x"3712",x"3b92",x"b509",x"2cb0",x"3b3e",x"3866"),
(x"1c5d",x"3e35",x"36eb",x"b046",x"3be8",x"2cb7",x"3b34",x"3832",x"216e",x"3e39",x"36eb",x"b9e9",x"3955",x"2e31",x"3b34",x"382e",x"2072",x"3e36",x"3710",x"b833",x"3ac7",x"2d1d",x"3b2f",x"3831"),
(x"1f0d",x"3e22",x"3713",x"37c3",x"baf3",x"2e28",x"3b86",x"3a5b",x"1fba",x"3e21",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b8a",x"3a5c",x"16e7",x"3e1d",x"370f",x"3ad7",x"b821",x"29e6",x"3b87",x"3a57"),
(x"9d26",x"3e23",x"36eb",x"baff",x"373c",x"3197",x"3a3f",x"3a50",x"1986",x"3e2a",x"36eb",x"b97a",x"39b6",x"309a",x"3a3f",x"3a4b",x"9aec",x"3e22",x"3717",x"ba77",x"3889",x"310e",x"3a3a",x"3a50"),
(x"9aa8",x"3e77",x"3718",x"b0c5",x"bbe6",x"2ad9",x"3b2f",x"38b5",x"9950",x"3e76",x"36eb",x"bb01",x"b745",x"3141",x"3b32",x"38b9",x"9fe7",x"3e77",x"3719",x"b250",x"bbca",x"2f22",x"3b30",x"38b3"),
(x"2422",x"3e7d",x"36eb",x"3b99",x"b45f",x"30d6",x"3b44",x"3870",x"1fbf",x"3e6a",x"36eb",x"3b57",x"b625",x"2e99",x"3b43",x"3865",x"2353",x"3e7c",x"3711",x"3b70",x"b585",x"3014",x"3b3f",x"3870"),
(x"9a03",x"3e37",x"36eb",x"374a",x"3b15",x"2de4",x"3b35",x"3836",x"1c5d",x"3e35",x"36eb",x"b046",x"3be8",x"2cb7",x"3b34",x"3832",x"11f0",x"3e35",x"3712",x"32e8",x"3bcb",x"2c10",x"3b30",x"3835"),
(x"20b1",x"3e20",x"36eb",x"b8ae",x"ba73",x"2d47",x"3b1b",x"3b2e",x"1fba",x"3e21",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b1b",x"3b2d",x"2079",x"3e21",x"3712",x"b721",x"bb24",x"2bf9",x"3b17",x"3b30"),
(x"a139",x"3e14",x"36eb",x"bbbf",x"3113",x"322d",x"3a3f",x"3a58",x"9d26",x"3e23",x"36eb",x"baff",x"373c",x"3197",x"3a3f",x"3a50",x"a039",x"3e14",x"3713",x"bbc6",x"31be",x"30de",x"3a3a",x"3a57"),
(x"24be",x"3e8c",x"36eb",x"3be6",x"ac77",x"308c",x"3b44",x"3878",x"2422",x"3e7d",x"36eb",x"3b99",x"b45f",x"30d6",x"3b44",x"3870",x"2467",x"3e8c",x"3711",x"3be4",x"ad1e",x"308c",x"3b40",x"3878"),
(x"a0d7",x"3e3d",x"3717",x"3b6f",x"35e5",x"261e",x"3b32",x"383c",x"a09f",x"3e3d",x"36eb",x"3aaf",x"3860",x"2a70",x"3b37",x"383a",x"9ad5",x"3e36",x"3711",x"3934",x"3a0d",x"2c18",x"3b31",x"3837"),
(x"21ab",x"3e1e",x"36eb",x"ae29",x"bbe6",x"3005",x"3b1c",x"3b2f",x"20b1",x"3e20",x"36eb",x"b8ae",x"ba73",x"2d47",x"3b1b",x"3b2e",x"21e0",x"3e1f",x"3711",x"b5dd",x"bb65",x"2eae",x"3b18",x"3b32"),
(x"a08e",x"3e07",x"3717",x"bbf0",x"2f10",x"2aec",x"3a39",x"3a5e",x"a0d9",x"3e07",x"36eb",x"bbea",x"2e09",x"2f12",x"3a3e",x"3a5f",x"a039",x"3e14",x"3713",x"bbc6",x"31be",x"30de",x"3a3a",x"3a57"),
(x"9950",x"3e76",x"36eb",x"bb01",x"b745",x"3141",x"3b82",x"396a",x"9aa8",x"3e77",x"3718",x"b0c5",x"bbe6",x"2ad9",x"3b82",x"3970",x"9920",x"3e76",x"3718",x"baf6",x"37e1",x"2460",x"3b82",x"3970"),
(x"2469",x"3e9d",x"3714",x"3bec",x"2d02",x"2f48",x"3b40",x"3881",x"24b3",x"3e9d",x"36eb",x"3be8",x"2d66",x"3010",x"3b45",x"3881",x"2467",x"3e8c",x"3711",x"3be4",x"ad1e",x"308c",x"3b40",x"3878"),
(x"a180",x"3e45",x"3715",x"3bfe",x"a412",x"2867",x"3b33",x"3840",x"a166",x"3e45",x"36eb",x"3bfa",x"2c62",x"2617",x"3b38",x"383e",x"a0d7",x"3e3d",x"3717",x"3b6f",x"35e5",x"261e",x"3b32",x"383c"),
(x"244f",x"3e1f",x"36eb",x"3913",x"ba0d",x"310f",x"3b1e",x"3b32",x"21ab",x"3e1e",x"36eb",x"ae29",x"bbe6",x"3005",x"3b1c",x"3b2f",x"23f2",x"3e20",x"3712",x"35a5",x"bb63",x"30cc",x"3b19",x"3b34"),
(x"a243",x"3dfc",x"36eb",x"bbe4",x"2adf",x"30ee",x"3a3d",x"3a65",x"a0d9",x"3e07",x"36eb",x"bbea",x"2e09",x"2f12",x"3a3e",x"3a5f",x"a1a0",x"3dfc",x"370f",x"bbdd",x"30de",x"2e6c",x"3a39",x"3a64"),
(x"a164",x"3e6e",x"36eb",x"bbbf",x"3333",x"2ed0",x"3b87",x"3969",x"9fd8",x"3e72",x"36eb",x"ba0e",x"3929",x"2e76",x"3b85",x"396a",x"a0a3",x"3e6e",x"3718",x"bb13",x"3732",x"2fec",x"3b87",x"396f"),
(x"2427",x"3ea6",x"36eb",x"3ab2",x"3834",x"30cb",x"3b45",x"3886",x"24b3",x"3e9d",x"36eb",x"3be8",x"2d66",x"3010",x"3b45",x"3881",x"23cf",x"3ea5",x"3712",x"3b45",x"3640",x"30a6",x"3b40",x"3885"),
(x"1ea1",x"3e94",x"3710",x"3bcc",x"3228",x"2f2f",x"3b3a",x"3b30",x"1f98",x"3e94",x"36eb",x"3bf4",x"1edc",x"2ebb",x"3b3f",x"3b2f",x"1de8",x"3e90",x"3710",x"3b2f",x"b6d9",x"2e52",x"3b3a",x"3b2d"),
(x"a123",x"3e50",x"3714",x"3b81",x"b558",x"2da5",x"3b35",x"3845",x"a0d8",x"3e4f",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"3b3a",x"3843",x"a180",x"3e45",x"3715",x"3bfe",x"a412",x"2867",x"3b33",x"3840"),
(x"24ee",x"3e23",x"36eb",x"3be5",x"2dbc",x"3036",x"3b1f",x"3b34",x"244f",x"3e1f",x"36eb",x"3913",x"ba0d",x"310f",x"3b1e",x"3b32",x"2498",x"3e24",x"3711",x"3bb2",x"b32f",x"30f4",x"3b1a",x"3b36"),
(x"a1da",x"3df6",x"36eb",x"baf6",x"b714",x"32f0",x"3a3d",x"3a68",x"a243",x"3dfc",x"36eb",x"bbe4",x"2adf",x"30ee",x"3a3d",x"3a65",x"a12d",x"3df8",x"370d",x"bb0d",x"b70c",x"3169",x"3a39",x"3a66"),
(x"a13e",x"3e68",x"36eb",x"bbbf",x"b370",x"2dad",x"3b8a",x"3969",x"a164",x"3e6e",x"36eb",x"bbbf",x"3333",x"2ed0",x"3b87",x"3969",x"a0f6",x"3e69",x"3712",x"bbf0",x"ac20",x"2e95",x"3b8a",x"396e"),
(x"20e4",x"3eae",x"36eb",x"37cb",x"3ae6",x"3068",x"3b45",x"388b",x"2427",x"3ea6",x"36eb",x"3ab2",x"3834",x"30cb",x"3b45",x"3886",x"20a5",x"3eac",x"3715",x"393c",x"39e9",x"3110",x"3b40",x"388b"),
(x"9e13",x"3e58",x"3715",x"3a65",x"b8c1",x"2d9c",x"3b36",x"384a",x"9d2f",x"3e57",x"36eb",x"3ac2",x"b833",x"2e8a",x"3b3b",x"3848",x"a123",x"3e50",x"3714",x"3b81",x"b558",x"2da5",x"3b35",x"3845"),
(x"2454",x"3e2b",x"36eb",x"3902",x"3a23",x"306a",x"3b20",x"3b38",x"24ee",x"3e23",x"36eb",x"3be5",x"2dbc",x"3036",x"3b1f",x"3b34",x"242c",x"3e29",x"3712",x"3ae4",x"37c3",x"30c9",x"3b1b",x"3b39"),
(x"a05e",x"3df6",x"3713",x"b451",x"bbac",x"2d81",x"3a38",x"3a67",x"a088",x"3df5",x"36eb",x"b571",x"bb6d",x"30cc",x"3a3d",x"3a69",x"a12d",x"3df8",x"370d",x"bb0d",x"b70c",x"3169",x"3a39",x"3a66"),
(x"a0e1",x"3e67",x"36eb",x"aeda",x"bbea",x"2e47",x"3b8b",x"3969",x"a13e",x"3e68",x"36eb",x"bbbf",x"b370",x"2dad",x"3b8a",x"3969",x"a072",x"3e68",x"3712",x"b297",x"bbcc",x"2d84",x"3b8b",x"396f"),
(x"177f",x"3eb0",x"36eb",x"175f",x"3bf5",x"2e99",x"3b44",x"3890",x"20e4",x"3eae",x"36eb",x"37cb",x"3ae6",x"3068",x"3b45",x"388b",x"1788",x"3eaf",x"3715",x"1ef6",x"3bee",x"302a",x"3b3f",x"388f"),
(x"9607",x"3e5d",x"3717",x"3939",x"ba0b",x"29e0",x"3b38",x"384d",x"9470",x"3e5c",x"36eb",x"39cd",x"b979",x"2caa",x"3b3c",x"384b",x"9e13",x"3e58",x"3715",x"3a65",x"b8c1",x"2d9c",x"3b36",x"384a"),
(x"21e1",x"3e2c",x"36eb",x"33f1",x"3bbc",x"2b5c",x"3b20",x"3b3b",x"2454",x"3e2b",x"36eb",x"3902",x"3a23",x"306a",x"3b20",x"3b38",x"2226",x"3e2b",x"3713",x"3607",x"3b5e",x"2e4f",x"3b1b",x"3b3b"),
(x"9e25",x"3df6",x"3716",x"b8de",x"ba57",x"297d",x"3a37",x"3a68",x"9e52",x"3df5",x"36eb",x"bbe3",x"ace8",x"30c3",x"3a3c",x"3a6b",x"a05e",x"3df6",x"3713",x"b451",x"bbac",x"2d81",x"3a38",x"3a67"),
(x"9d58",x"3e68",x"3717",x"aa07",x"bbfc",x"284d",x"3b8c",x"3970",x"9ce6",x"3e67",x"36eb",x"ac58",x"bbf7",x"2bc5",x"3b8d",x"396a",x"a072",x"3e68",x"3712",x"b297",x"bbcc",x"2d84",x"3b8b",x"396f"),
(x"9e4d",x"3ead",x"3713",x"b82e",x"3aba",x"306c",x"3b3f",x"3893",x"9dfd",x"3eae",x"36eb",x"b66a",x"3b44",x"2f81",x"3b43",x"3894",x"1788",x"3eaf",x"3715",x"1ef6",x"3bee",x"302a",x"3b3f",x"388f"),
(x"125b",x"3e5e",x"3717",x"ac95",x"bbf9",x"2918",x"3b38",x"384e",x"11e3",x"3e5e",x"36eb",x"b5a6",x"bb74",x"2d53",x"3b3d",x"384c",x"9607",x"3e5d",x"3717",x"3939",x"ba0b",x"29e0",x"3b38",x"384d"),
(x"212c",x"3e2d",x"3716",x"3ac7",x"b83c",x"283f",x"3b1b",x"3b3d",x"2164",x"3e2d",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b20",x"3b3c",x"2226",x"3e2b",x"3713",x"3607",x"3b5e",x"2e4f",x"3b1b",x"3b3b"),
(x"1624",x"3e08",x"370e",x"3004",x"271d",x"3bef",x"3b6b",x"3b29",x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a",x"a08e",x"3e07",x"3717",x"2bf6",x"a5ae",x"3bfb",x"3b62",x"3b29"),
(x"9b62",x"3e66",x"36eb",x"ba75",x"b8ad",x"2ccc",x"3b8e",x"396a",x"9ce6",x"3e67",x"36eb",x"ac58",x"bbf7",x"2bc5",x"3b8d",x"396a",x"9b02",x"3e67",x"3716",x"b8f4",x"ba42",x"2c09",x"3b8d",x"3970"),
(x"a2e7",x"3ea6",x"3715",x"bae0",x"37cf",x"30d4",x"3b3d",x"3898",x"a395",x"3ea8",x"36eb",x"b9f2",x"3938",x"30b5",x"3b42",x"389a",x"9e4d",x"3ead",x"3713",x"b82e",x"3aba",x"306c",x"3b3f",x"3893"),
(x"1e32",x"3e58",x"36eb",x"b976",x"b9cc",x"2dcc",x"3b3f",x"3850",x"11e3",x"3e5e",x"36eb",x"b5a6",x"bb74",x"2d53",x"3b3d",x"384c",x"1acb",x"3e5c",x"3714",x"b9a7",x"b99e",x"2d1e",x"3b39",x"3850"),
(x"2433",x"3e2e",x"36eb",x"39ec",x"b92b",x"31e4",x"3b20",x"3b3f",x"2164",x"3e2d",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b20",x"3b3c",x"2360",x"3e2f",x"3711",x"38c8",x"ba4e",x"30a8",x"3b1c",x"3b3f"),
(x"9b62",x"3e66",x"36eb",x"ba75",x"b8ad",x"2ccc",x"3b8e",x"396a",x"9b02",x"3e67",x"3716",x"b8f4",x"ba42",x"2c09",x"3b8d",x"3970",x"9959",x"3e66",x"3715",x"bb3f",x"b6b6",x"2b9d",x"3b8e",x"3970"),
(x"a44d",x"3e9d",x"3715",x"bbec",x"2be2",x"2fce",x"3b3c",x"389d",x"a493",x"3e9e",x"36eb",x"bbc4",x"327a",x"3012",x"3b40",x"389e",x"a2e7",x"3ea6",x"3715",x"bae0",x"37cf",x"30d4",x"3b3d",x"3898"),
(x"20ef",x"3e55",x"36eb",x"b53f",x"bb87",x"2d28",x"3b40",x"3852",x"1e32",x"3e58",x"36eb",x"b976",x"b9cc",x"2dcc",x"3b3f",x"3850",x"2116",x"3e56",x"3716",x"b7d5",x"baf0",x"2d8e",x"3b3b",x"3854"),
(x"2563",x"3e37",x"36eb",x"3bbc",x"b212",x"3175",x"3b20",x"3b44",x"2433",x"3e2e",x"36eb",x"39ec",x"b92b",x"31e4",x"3b20",x"3b3f",x"24fa",x"3e37",x"370f",x"3b4b",x"b5cc",x"3223",x"3b1c",x"3b44"),
(x"9f92",x"3de3",x"36eb",x"bade",x"b7ab",x"31d3",x"3b8f",x"3a2a",x"a0ba",x"3def",x"36eb",x"bbdb",x"9c67",x"320a",x"3b8c",x"3a25",x"9e24",x"3de5",x"370e",x"bb7b",x"b4a9",x"3270",x"3b8b",x"3a2c"),
(x"a0d7",x"3e5f",x"36eb",x"bafe",x"375c",x"30f4",x"3a3d",x"3a29",x"9959",x"3e66",x"3715",x"ba5f",x"3874",x"3388",x"3a37",x"3a24",x"9ec5",x"3e5f",x"3718",x"bac6",x"37dc",x"3286",x"3a38",x"3a28"),
(x"a409",x"3e95",x"3717",x"bb55",x"b5fd",x"307e",x"3b3a",x"38a1",x"a46a",x"3e94",x"36eb",x"bb6e",x"b575",x"309e",x"3b3f",x"38a3",x"a44d",x"3e9d",x"3715",x"bbec",x"2be2",x"2fce",x"3b3c",x"389d"),
(x"2353",x"3e7c",x"3711",x"3115",x"a7d5",x"3be4",x"3b78",x"3b8d",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c",x"2002",x"3e80",x"3714",x"305e",x"a194",x"3bec",x"3b72",x"3b90"),
(x"2357",x"3e54",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3b41",x"3854",x"20ef",x"3e55",x"36eb",x"b53f",x"bb87",x"2d28",x"3b40",x"3852",x"2323",x"3e55",x"3716",x"2345",x"bbf7",x"2dcc",x"3b3c",x"3856"),
(x"2574",x"3e41",x"36eb",x"3b61",x"35a0",x"3119",x"3b20",x"3b4a",x"2563",x"3e37",x"36eb",x"3bbc",x"b212",x"3175",x"3b20",x"3b44",x"2517",x"3e40",x"370f",x"3bd3",x"2f46",x"3182",x"3b1c",x"3b49"),
(x"a348",x"3e53",x"36eb",x"bbba",x"3376",x"2f14",x"3a3e",x"3a2f",x"a0d7",x"3e5f",x"36eb",x"bafe",x"375c",x"30f4",x"3a3d",x"3a29",x"a29f",x"3e53",x"3714",x"bb6b",x"3587",x"3096",x"3a39",x"3a2f"),
(x"a22e",x"3e8d",x"36eb",x"b884",x"ba69",x"324a",x"3b3d",x"38a8",x"a46a",x"3e94",x"36eb",x"bb6e",x"b575",x"309e",x"3b3f",x"38a3",x"a18f",x"3e8e",x"3711",x"b8a4",x"ba69",x"309a",x"3b39",x"38a5"),
(x"24b8",x"3e56",x"36eb",x"3acc",x"b812",x"3064",x"3b41",x"3856",x"2357",x"3e54",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3b41",x"3854",x"245f",x"3e57",x"3714",x"3976",x"b9c0",x"3023",x"3b3c",x"3858"),
(x"2449",x"3e47",x"36eb",x"386e",x"3a87",x"313e",x"3b20",x"3b4e",x"2574",x"3e41",x"36eb",x"3b61",x"35a0",x"3119",x"3b20",x"3b4a",x"2437",x"3e45",x"370f",x"3891",x"3a72",x"30f5",x"3b1b",x"3b4c"),
(x"1222",x"3dd9",x"36eb",x"b8a6",x"ba54",x"3207",x"3b91",x"3a31",x"9f92",x"3de3",x"36eb",x"bade",x"b7ab",x"31d3",x"3b8f",x"3a2a",x"0f4a",x"3ddc",x"3712",x"b8b5",x"ba3e",x"32bd",x"3b8d",x"3a32"),
(x"a41c",x"3e46",x"36eb",x"bbef",x"ad09",x"2e69",x"3a3f",x"3a36",x"a348",x"3e53",x"36eb",x"bbba",x"3376",x"2f14",x"3a3e",x"3a2f",x"a3b3",x"3e47",x"3712",x"bbf0",x"2a00",x"2f46",x"3a3a",x"3a36"),
(x"9a89",x"3e8b",x"3718",x"b8ae",x"ba78",x"2b7c",x"3b36",x"38a8",x"9bc5",x"3e8b",x"36eb",x"b60d",x"bb5a",x"2ef3",x"3b3a",x"38ab",x"a18f",x"3e8e",x"3711",x"b8a4",x"ba69",x"309a",x"3b39",x"38a5"),
(x"2515",x"3e5c",x"36eb",x"3bcf",x"3174",x"303e",x"3b42",x"3859",x"24b8",x"3e56",x"36eb",x"3acc",x"b812",x"3064",x"3b41",x"3856",x"24ba",x"3e5b",x"3712",x"3be0",x"ae5e",x"30a3",x"3b3d",x"385a"),
(x"221a",x"3e47",x"3713",x"b583",x"3b63",x"3153",x"3b1a",x"3b4f",x"21a6",x"3e48",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b1f",x"3b51",x"2437",x"3e45",x"370f",x"3891",x"3a72",x"30f5",x"3b1b",x"3b4c"),
(x"1c89",x"3ddc",x"3716",x"3add",x"b75a",x"334d",x"3b8c",x"3a34",x"1dd1",x"3dd9",x"36eb",x"3996",x"b95e",x"33ec",x"3b92",x"3a33",x"0f4a",x"3ddc",x"3712",x"b8b5",x"ba3e",x"32bd",x"3b8d",x"3a32"),
(x"a2ed",x"3e3a",x"36eb",x"bb75",x"b5a2",x"2d46",x"3a3f",x"3a3c",x"a41c",x"3e46",x"36eb",x"bbef",x"ad09",x"2e69",x"3a3f",x"3a36",x"a294",x"3e3b",x"3710",x"bb6a",x"b5bb",x"2efe",x"3a3b",x"3a3c"),
(x"9747",x"3e88",x"3718",x"bbe6",x"b09f",x"2baa",x"3b35",x"38aa",x"990f",x"3e89",x"36eb",x"bbe6",x"b08f",x"2c41",x"3b3a",x"38ac",x"9a89",x"3e8b",x"3718",x"b8ae",x"ba78",x"2b7c",x"3b36",x"38a8"),
(x"247a",x"3e61",x"36eb",x"36fe",x"3b25",x"2ea4",x"3b42",x"385c",x"2515",x"3e5c",x"36eb",x"3bcf",x"3174",x"303e",x"3b42",x"3859",x"2458",x"3e5f",x"3714",x"3972",x"39bb",x"30de",x"3b3d",x"385c"),
(x"235a",x"3e97",x"3710",x"a828",x"a60a",x"3bfe",x"3b78",x"3ba3",x"2325",x"3e9e",x"3714",x"a946",x"9ffc",x"3bfe",x"3b78",x"3baa",x"2469",x"3e9d",x"3714",x"aeb0",x"a8fa",x"3bf3",x"3b7b",x"3ba9"),
(x"227e",x"3ea3",x"3712",x"a953",x"a7b4",x"3bfd",x"3b77",x"3bad",x"214b",x"3ea6",x"3714",x"28bf",x"ac22",x"3bfa",x"3b76",x"3bb0",x"23cf",x"3ea5",x"3712",x"2587",x"a09b",x"3bff",x"3b79",x"3baf"),
(x"1f1f",x"3ea8",x"3714",x"a31d",x"ab5f",x"3bfc",x"3b73",x"3bb3",x"20a5",x"3eac",x"3715",x"20ea",x"aafd",x"3bfc",x"3b75",x"3bb6",x"214b",x"3ea6",x"3714",x"28bf",x"ac22",x"3bfa",x"3b76",x"3bb0"),
(x"11db",x"3eaa",x"3715",x"a70a",x"2773",x"3bfe",x"3b6e",x"3bb4",x"1788",x"3eaf",x"3715",x"a7e2",x"a9b5",x"3bfc",x"3b6f",x"3bb9",x"1f1f",x"3ea8",x"3714",x"a31d",x"ab5f",x"3bfc",x"3b73",x"3bb3"),
(x"9d99",x"3ea9",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3b69",x"3bb4",x"9e4d",x"3ead",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3b69",x"3bb7",x"11db",x"3eaa",x"3715",x"a70a",x"2773",x"3bfe",x"3b6e",x"3bb4"),
(x"a14f",x"3ea3",x"3714",x"28e0",x"a99e",x"3bfc",x"3b65",x"3baf",x"a2e7",x"3ea6",x"3715",x"2266",x"1d87",x"3bff",x"3b62",x"3bb2",x"9d99",x"3ea9",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3b69",x"3bb4"),
(x"a1ee",x"3e9d",x"3714",x"2538",x"29ab",x"3bfd",x"3b63",x"3baa",x"a44d",x"3e9d",x"3715",x"2891",x"27ce",x"3bfd",x"3b5f",x"3baa",x"a14f",x"3ea3",x"3714",x"28e0",x"a99e",x"3bfc",x"3b65",x"3baf"),
(x"a1ee",x"3e9d",x"3714",x"2538",x"29ab",x"3bfd",x"3b63",x"3baa",x"a0ed",x"3e98",x"3715",x"2c67",x"a8a5",x"3bf9",x"3b65",x"3ba6",x"a44d",x"3e9d",x"3715",x"2891",x"27ce",x"3bfd",x"3b5f",x"3baa"),
(x"9ddf",x"3e98",x"3714",x"2a45",x"ab10",x"3bfa",x"3b68",x"3ba5",x"a18f",x"3e8e",x"3711",x"28d9",x"252b",x"3bfe",x"3b63",x"3b9d",x"a0ed",x"3e98",x"3715",x"2c67",x"a8a5",x"3bf9",x"3b65",x"3ba6"),
(x"1937",x"3e9a",x"3710",x"2352",x"2e7e",x"3bf5",x"3b6f",x"3ba7",x"1d11",x"3e98",x"3711",x"2bef",x"28a8",x"3bfa",x"3b71",x"3ba4",x"9908",x"3e9a",x"3711",x"2a66",x"331a",x"3bca",x"3b6b",x"3ba7"),
(x"9747",x"3e88",x"3718",x"3420",x"9418",x"3bba",x"3b6a",x"3b97",x"9a89",x"3e8b",x"3718",x"2b65",x"3528",x"3b8f",x"3b69",x"3b9a",x"18c5",x"3e8c",x"3713",x"341f",x"2c3a",x"3bb6",x"3b6e",x"3b9a"),
(x"1832",x"3e87",x"3714",x"2de0",x"24c2",x"3bf6",x"3b6e",x"3b96",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c",x"9613",x"3e7f",x"3715",x"27ae",x"24ea",x"3bfe",x"3b6b",x"3b8f"),
(x"1d11",x"3e98",x"3711",x"2bef",x"28a8",x"3bfa",x"3b71",x"3ba4",x"1de8",x"3e90",x"3710",x"2856",x"29ab",x"3bfc",x"3b71",x"3b9e",x"9ddf",x"3e98",x"3714",x"2a45",x"ab10",x"3bfa",x"3b68",x"3ba5"),
(x"98e9",x"3e7d",x"3715",x"a8bf",x"2fdb",x"3bef",x"3b6a",x"3b8d",x"9613",x"3e7f",x"3715",x"27ae",x"24ea",x"3bfe",x"3b6b",x"3b8f",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c"),
(x"199d",x"3e8c",x"36eb",x"3bf6",x"aa70",x"2d61",x"3b3e",x"3b29",x"1c29",x"3e7b",x"36eb",x"346a",x"3b91",x"316a",x"3b3c",x"3b21",x"1832",x"3e87",x"3714",x"3bf3",x"2e23",x"2b27",x"3b38",x"3b28"),
(x"22bc",x"3f52",x"36eb",x"3adb",x"b7e7",x"30ac",x"3b35",x"3b2b",x"1f7b",x"3f4a",x"36eb",x"3b71",x"b58a",x"2fc3",x"3b35",x"3b26",x"1e77",x"3f4b",x"3715",x"3ac2",x"b812",x"3146",x"3b30",x"3b26"),
(x"b931",x"3d45",x"3710",x"bbe9",x"26a1",x"309e",x"3a36",x"33ca",x"b930",x"3d5c",x"3710",x"bbeb",x"2604",x"3075",x"3a49",x"33c0",x"b92b",x"3d45",x"3732",x"bb64",x"243f",x"361b",x"3a35",x"33aa"),
(x"b92b",x"3d45",x"3732",x"bb64",x"243f",x"361b",x"3a35",x"33aa",x"b92a",x"3d5c",x"3733",x"bb1e",x"251e",x"3748",x"3a49",x"339f",x"b924",x"3d45",x"3749",x"ba3b",x"267a",x"3902",x"3a35",x"3392"),
(x"b924",x"3d45",x"3749",x"ba3b",x"267a",x"3902",x"3a35",x"3392",x"b922",x"3d5c",x"3748",x"b86c",x"29d9",x"3aa7",x"3a48",x"3388",x"b91f",x"3d45",x"374e",x"ac96",x"29b2",x"3bf8",x"3a34",x"3387"),
(x"b91f",x"3d45",x"374e",x"ac96",x"29b2",x"3bf8",x"3a34",x"3387",x"b91b",x"3d5c",x"3749",x"3594",x"2b76",x"3b7b",x"3a48",x"337b",x"b918",x"3d45",x"374b",x"38f0",x"29d6",x"3a48",x"3a34",x"337b"),
(x"b907",x"3d5d",x"3713",x"2f5d",x"3bdb",x"30c1",x"3bc3",x"39d6",x"b913",x"3d5c",x"373b",x"381d",x"3a67",x"34eb",x"3bbd",x"39cf",x"b90e",x"3d5d",x"370e",x"3754",x"3ae5",x"32eb",x"3bc0",x"39d7"),
(x"b91b",x"3d5e",x"374a",x"3544",x"b37e",x"3b51",x"3bb9",x"39cc",x"b913",x"3d5e",x"373a",x"3ae3",x"2b4f",x"380a",x"3bbc",x"39cf",x"b91b",x"3d5c",x"3749",x"382b",x"a439",x"3ad3",x"3bbb",x"39cb"),
(x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e",x"b906",x"3d45",x"3710",x"2e12",x"a66c",x"3bf6",x"3a34",x"333e",x"b90c",x"3d45",x"3724",x"3af5",x"1a59",x"37e2",x"3a34",x"3352"),
(x"b90f",x"3d73",x"3727",x"3bc1",x"a904",x"33bf",x"3bfb",x"3974",x"b90d",x"3d73",x"3711",x"3be1",x"a6cf",x"3179",x"3bfb",x"396f",x"b90e",x"3d5d",x"370e",x"3bcb",x"a946",x"330f",x"3bea",x"3970"),
(x"b91a",x"3d72",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"397c",x"b913",x"3d73",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"3978",x"b91b",x"3d5e",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"397d"),
(x"b922",x"3d72",x"3751",x"a11e",x"aa52",x"3bfd",x"3bfb",x"397f",x"b91a",x"3d72",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"397c",x"b924",x"3d5e",x"374d",x"af62",x"aa90",x"3bef",x"3beb",x"3980"),
(x"b92b",x"3d5e",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"3984",x"b928",x"3d72",x"374d",x"b867",x"a907",x"3aab",x"3bfb",x"3982",x"b924",x"3d5e",x"374d",x"af62",x"aa90",x"3bef",x"3beb",x"3980"),
(x"b930",x"3d5e",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"3986",x"b92f",x"3d72",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"3986",x"b92b",x"3d5e",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"3984"),
(x"b938",x"3d5e",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"398f",x"b935",x"3d73",x"3725",x"bb50",x"a638",x"3678",x"3bfb",x"398b",x"b930",x"3d5e",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"3986"),
(x"b935",x"3d73",x"3725",x"bb50",x"a638",x"3678",x"3bfb",x"398b",x"b938",x"3d5e",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"398f",x"b93a",x"3d73",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3bfb",x"398f"),
(x"b938",x"3d5e",x"3710",x"b678",x"bb4d",x"2af3",x"3bba",x"39ba",x"b930",x"3d5e",x"3738",x"b75b",x"bae5",x"32d3",x"3bb7",x"39c3",x"b930",x"3d5c",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bbd",x"39bd"),
(x"b912",x"3d45",x"373c",x"3aea",x"2832",x"3802",x"3a34",x"336a",x"b918",x"3d45",x"374b",x"38f0",x"29d6",x"3a48",x"3a34",x"337b",x"b913",x"3d5c",x"373b",x"3aa1",x"2559",x"3879",x"3a48",x"3369"),
(x"b924",x"3d5e",x"374d",x"b1cf",x"b808",x"3ac1",x"3bb8",x"39c9",x"b91b",x"3d5e",x"374a",x"3544",x"b37e",x"3b51",x"3bb9",x"39cc",x"b922",x"3d5c",x"3748",x"b511",x"b92e",x"398b",x"3bba",x"39c9"),
(x"b924",x"3d5e",x"374d",x"b1cf",x"b808",x"3ac1",x"3bb8",x"39c9",x"b922",x"3d5c",x"3748",x"b511",x"b92e",x"398b",x"3bba",x"39c9",x"b92b",x"3d5e",x"3744",x"b778",x"ba1b",x"3724",x"3bb7",x"39c5"),
(x"b92a",x"3d5c",x"3733",x"b800",x"ba99",x"3437",x"3bba",x"39c3",x"b930",x"3d5e",x"3738",x"b75b",x"bae5",x"32d3",x"3bb7",x"39c3",x"b92b",x"3d5e",x"3744",x"b778",x"ba1b",x"3724",x"3bb7",x"39c5"),
(x"b92a",x"3d74",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3849",x"b935",x"3d73",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3843",x"b931",x"3d74",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3842"),
(x"b925",x"3d74",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"384d",x"b92f",x"3d72",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3848",x"b92a",x"3d74",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3849"),
(x"b920",x"3d74",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"384f",x"b928",x"3d72",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"384c",x"b925",x"3d74",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"384d"),
(x"b920",x"3d74",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"384f",x"b922",x"3d72",x"3751",x"9a8d",x"39ac",x"39a3",x"3b24",x"384f",x"b928",x"3d72",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"384c"),
(x"b919",x"3d74",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3851",x"b91a",x"3d72",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3851",x"b920",x"3d74",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"384f"),
(x"b913",x"3d74",x"373e",x"3b0f",x"a04d",x"3786",x"3b1e",x"3853",x"b913",x"3d73",x"373e",x"3a5b",x"3409",x"386a",x"3b1f",x"3854",x"b919",x"3d74",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3851"),
(x"b90b",x"3d74",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3857",x"b90f",x"3d73",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3857",x"b913",x"3d74",x"373e",x"3b0f",x"a04d",x"3786",x"3b1e",x"3853"),
(x"b90b",x"3d74",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3857",x"b90d",x"3d73",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"385a",x"b90f",x"3d73",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3857"),
(x"b906",x"3d73",x"3713",x"2edc",x"bb7b",x"3565",x"3b16",x"3858",x"b90d",x"3d73",x"3711",x"368c",x"bb0e",x"3375",x"3b18",x"385a",x"b90b",x"3d74",x"371c",x"391c",x"b988",x"3561",x"3b19",x"3857"),
(x"b90e",x"3d5d",x"370e",x"b4eb",x"a6e9",x"3b9c",x"3a49",x"334b",x"b90d",x"3d73",x"3711",x"b36e",x"a40b",x"3bc7",x"3a5b",x"3349",x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e"),
(x"b931",x"3d8b",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a6f",x"33c9",x"b92f",x"3d8b",x"372b",x"bbac",x"a891",x"347c",x"3a6f",x"33b1",x"b931",x"3d74",x"3710",x"bbea",x"a7ae",x"307d",x"3a5b",x"33c4"),
(x"b92a",x"3d74",x"3739",x"bb13",x"a8dd",x"3771",x"3a5c",x"339e",x"b92f",x"3d8b",x"372b",x"bbac",x"a891",x"347c",x"3a6f",x"33b1",x"b92c",x"3d8b",x"373a",x"baa5",x"a5fd",x"3872",x"3a6f",x"33a3"),
(x"b925",x"3d74",x"3746",x"b918",x"a84d",x"3a28",x"3a5c",x"338e",x"b92a",x"3d74",x"3739",x"bb13",x"a8dd",x"3771",x"3a5c",x"339e",x"b925",x"3d8a",x"3749",x"b926",x"a7c8",x"3a1d",x"3a6f",x"3391"),
(x"b91f",x"3d8a",x"374f",x"a812",x"a959",x"3bfd",x"3a6f",x"3385",x"b920",x"3d74",x"374b",x"b451",x"a960",x"3bb2",x"3a5c",x"3385",x"b925",x"3d8a",x"3749",x"b926",x"a7c8",x"3a1d",x"3a6f",x"3391"),
(x"b918",x"3d8a",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a6f",x"3378",x"b919",x"3d74",x"3749",x"3647",x"a97a",x"3b59",x"3a5c",x"3379",x"b91f",x"3d8a",x"374f",x"a812",x"a959",x"3bfd",x"3a6f",x"3385"),
(x"b911",x"3d8a",x"373c",x"3ac9",x"a6b5",x"383a",x"3a6f",x"3366",x"b913",x"3d74",x"373e",x"3ac8",x"a7bb",x"383c",x"3a5c",x"336a",x"b918",x"3d8a",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a6f",x"3378"),
(x"b90b",x"3d74",x"371c",x"3aa9",x"a818",x"386b",x"3a5c",x"334a",x"b913",x"3d74",x"373e",x"3ac8",x"a7bb",x"383c",x"3a5c",x"336a",x"b90b",x"3d8a",x"3722",x"3b0f",x"a82c",x"3781",x"3a6f",x"334c"),
(x"b906",x"3d73",x"3713",x"29ab",x"208e",x"3bfd",x"3a5b",x"333d",x"b90b",x"3d74",x"371c",x"3aa9",x"a818",x"386b",x"3a5c",x"334a",x"b907",x"3d8a",x"3718",x"38f7",x"a86d",x"3a44",x"3a6f",x"3340"),
(x"b135",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"24c1",x"b116",x"3d6c",x"3710",x"0000",x"8000",x"3c00",x"3a55",x"2451",x"b135",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"24c1"),
(x"b161",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"255f",x"b135",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"24c1",x"b161",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"255f"),
(x"b161",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"255f",x"b161",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"255f",x"b1a1",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2643"),
(x"b1c1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"26b3",x"b1a1",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2643",x"b1c1",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"26b3"),
(x"b1fd",x"3d79",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"278b",x"b1c1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"26b3",x"b1fd",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"278b"),
(x"b1fd",x"3d79",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"278b",x"b1fd",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"278b",x"b22d",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"281a"),
(x"b261",x"3d79",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2878",x"b22d",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"281a",x"b261",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2878"),
(x"b261",x"3d79",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2878",x"b261",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2878",x"b2aa",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"28fb"),
(x"b2d6",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2949",x"b2aa",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"28fb",x"b2d6",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2949"),
(x"b326",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a58",x"29d7",x"b2d6",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2949",x"b326",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4b",x"29d7"),
(x"b326",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a58",x"29d7",x"b326",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4b",x"29d7",x"b34f",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2a20"),
(x"b451",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2c3f",x"b451",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2c3f",x"b50c",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2d8d"),
(x"b441",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2c23",x"b451",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2c3f",x"b441",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2c23"),
(x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b",x"b441",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2c23",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b"),
(x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b",x"b34f",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2a20"),
(x"b413",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2ba0",x"b40b",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2b84",x"b413",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"2ba0"),
(x"b413",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"2ba0",x"b3f4",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2b48",x"b409",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2b7d"),
(x"b409",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2b7d",x"b3d2",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2b0a",x"b407",x"3d7d",x"3710",x"0000",x"8cea",x"3c00",x"3a63",x"2b76"),
(x"b3f4",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2b48",x"b40b",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2b84",x"b413",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2ba0"),
(x"b3d2",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2b0a",x"b3f4",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2b48",x"b409",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2b7d"),
(x"b3a5",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2aba",x"b3d2",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2b0a",x"b407",x"3d53",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2b76"),
(x"b368",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2a4d",x"b3a5",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2aba",x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b"),
(x"b407",x"3d7d",x"3710",x"0000",x"8cea",x"3c00",x"3a63",x"2b76",x"b3a5",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2aba",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b"),
(x"b368",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a68",x"2a4d",x"b340",x"3d7c",x"3710",x"0000",x"8000",x"3c00",x"3a63",x"2a04",x"b351",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2a22"),
(x"b526",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2dbb",x"b50c",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2d8d",x"b526",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2dbb"),
(x"b5ce",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2ee7",x"b62a",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2f8b",x"b5ce",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2ee7"),
(x"b5bd",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2ec9",x"b5ce",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2ee7",x"b5bd",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ec9"),
(x"b5a1",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2e97",x"b5bd",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2ec9",x"b5a1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2e97"),
(x"b581",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2e5e",x"b5a1",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2e97",x"b581",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2e5e"),
(x"b581",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2e5e",x"b581",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2e5e",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b52b",x"3d8d",x"3710",x"0000",x"8000",x"3c00",x"3a72",x"2dc4",x"b50d",x"3d8e",x"3710",x"0000",x"8000",x"3c00",x"3a72",x"2d8e",x"b4f5",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"2d63"),
(x"b544",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"2df0",x"b52b",x"3d8d",x"3710",x"0000",x"8000",x"3c00",x"3a72",x"2dc4",x"b4f2",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2d5e"),
(x"b52b",x"3d42",x"3710",x"0000",x"8000",x"3c00",x"3a31",x"2dc4",x"b4f5",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"2d63",x"b50d",x"3d41",x"3710",x"0000",x"8000",x"3c00",x"3a30",x"2d8e"),
(x"b544",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2df0",x"b4f2",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2d5e",x"b52b",x"3d42",x"3710",x"0000",x"8000",x"3c00",x"3a31",x"2dc4"),
(x"b558",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2e14",x"b568",x"3d46",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"2e32",x"b575",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2e47"),
(x"b544",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2df0",x"b558",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2e14",x"b569",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"2e33"),
(x"b575",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2e49",x"b568",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"2e32",x"b575",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2e47"),
(x"b575",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2e47",x"b558",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"2e14",x"b569",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"2e33"),
(x"b4d8",x"3d7c",x"3710",x"0000",x"8000",x"3c00",x"3a63",x"2d2f",x"b4e1",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2d40",x"b4da",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2d33"),
(x"b51a",x"3d58",x"3710",x"0000",x"8000",x"3c00",x"3a44",x"2da6",x"b4e1",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2d40",x"b4da",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2d33"),
(x"b528",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2dbf",x"b51a",x"3d58",x"3710",x"0000",x"8000",x"3c00",x"3a44",x"2da6",x"b4f2",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2d5e"),
(x"b4da",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2d33",x"b51a",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5f",x"2da6",x"b4f2",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2d5e"),
(x"b4f2",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2d5e",x"b528",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2dbf",x"b544",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"2df0"),
(x"b4f2",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2d5e",x"b544",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2df0",x"b528",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2dbf"),
(x"b569",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"2e33",x"b528",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2dbf",x"b568",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2e30"),
(x"b52c",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2dc5",x"b528",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2dbf",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b526",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2dbb",x"b526",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2dbb",x"b52c",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2dc5"),
(x"b568",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2e30",x"b52c",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2dc5",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b63d",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2fac",x"b62a",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2f8b",x"b63d",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2fac"),
(x"b669",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2ffc",x"b669",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ffc",x"b63d",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2fac"),
(x"b721",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"30a2",x"b669",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ffc",x"b721",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"30a2"),
(x"b72d",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"30ad",x"b72d",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"30ad",x"b721",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"30a2"),
(x"b794",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"3109",x"b7c0",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"3130",x"b794",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"3109"),
(x"b794",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"3109",x"b794",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"3109",x"b77a",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30f1"),
(x"b77a",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30f1",x"b77a",x"3d76",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"30f1",x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed"),
(x"b72d",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"30ad",x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed",x"b72d",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"30ad"),
(x"b705",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"3088",x"b6fb",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"3080",x"b6f1",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"3076"),
(x"b73e",x"3d44",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30bc",x"b721",x"3d59",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30a2",x"b705",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"3088"),
(x"b705",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"3088",x"b6f1",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"3076",x"b6fb",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"3080"),
(x"b73e",x"3d8c",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"30bc",x"b705",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"3088",x"b721",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5e",x"30a2"),
(x"b783",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"30f9",x"b73e",x"3d8c",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"30bc",x"b72e",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"30ae"),
(x"b783",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30f9",x"b72e",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"30ae",x"b73e",x"3d44",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30bc"),
(x"b7a4",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3117",x"b7c7",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"3135",x"b7bd",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3d",x"312d"),
(x"b7c7",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a68",x"3136",x"b7c7",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"3135",x"b7bd",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"312d"),
(x"b7bd",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"312d",x"b7a4",x"3d87",x"3710",x"0000",x"8000",x"3c00",x"3a6c",x"3117",x"b7a8",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"311a"),
(x"b783",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30f9",x"b7a4",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3117",x"b7a8",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"311a"),
(x"b72d",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"30ad",x"b72e",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"30ae",x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed"),
(x"b77b",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"30f2",x"b72e",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"30ae",x"b776",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"30ed"),
(x"b783",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30f9",x"b77b",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"30f2",x"b72e",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"30ae"),
(x"b77b",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"30f2",x"b783",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"30f9",x"b72e",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"30ae"),
(x"b801",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"316b",x"b801",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"316b",x"b7c0",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"3130"),
(x"b820",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"31a2",x"b820",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"31a2",x"b801",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"316b"),
(x"b83a",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"31d0",x"b83a",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"31d0",x"b820",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"31a2"),
(x"b84a",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"31ed",x"b84a",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"31ed",x"b83a",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"31d0"),
(x"b85e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3211",x"b85e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3211",x"b84a",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"31ed"),
(x"b865",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"321d",x"b865",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"321d",x"b85e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3211"),
(x"b867",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"3222",x"b867",x"3d81",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"3222",x"b865",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"321d"),
(x"b86e",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"322d",x"b867",x"3d81",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"3222",x"b86e",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"322d"),
(x"b87d",x"3d50",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"3248",x"b87d",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"3248",x"b86e",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"322d"),
(x"b88f",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"3269",x"b88f",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"3269",x"b87d",x"3d50",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"3248"),
(x"b89e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3284",x"b89e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3284",x"b88f",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"3269"),
(x"b8a3",x"3d47",x"3710",x"2081",x"9ea7",x"3bff",x"3a35",x"328d",x"b8a3",x"3d89",x"3710",x"2160",x"1cd0",x"3bff",x"3a6e",x"328d",x"b89e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3284"),
(x"b906",x"3d73",x"3713",x"29ab",x"208e",x"3bfd",x"3a5b",x"333d",x"b8a3",x"3d89",x"3710",x"2160",x"1cd0",x"3bff",x"3a6e",x"328d",x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e"),
(x"b907",x"3d8a",x"3718",x"38f7",x"a86d",x"3a44",x"3a6f",x"3340",x"b8ff",x"3d8a",x"3710",x"2904",x"26d5",x"3bfd",x"3a6f",x"3331",x"b906",x"3d73",x"3713",x"29ab",x"208e",x"3bfd",x"3a5b",x"333d"),
(x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e",x"b8a3",x"3d47",x"3710",x"2081",x"9ea7",x"3bff",x"3a35",x"328d",x"b906",x"3d45",x"3710",x"2e12",x"a66c",x"3bf6",x"3a34",x"333e"),
(x"b911",x"3d8a",x"373c",x"2504",x"3bff",x"2111",x"3bc3",x"3a1b",x"b918",x"3d8a",x"374b",x"270a",x"3bfd",x"287a",x"3bc0",x"3a1e",x"b925",x"3d8a",x"3749",x"257a",x"3bfd",x"28f4",x"3bc0",x"3a23"),
(x"b90b",x"3d8a",x"3722",x"2773",x"3bfe",x"22dc",x"3bc8",x"3a19",x"b911",x"3d8a",x"373c",x"2504",x"3bff",x"2111",x"3bc3",x"3a1b",x"b92c",x"3d8b",x"373a",x"25e9",x"3bff",x"17c8",x"3bc3",x"3a25"),
(x"b907",x"3d8a",x"3718",x"25bc",x"3bfe",x"2680",x"3bc9",x"3a17",x"b90b",x"3d8a",x"3722",x"2773",x"3bfe",x"22dc",x"3bc8",x"3a19",x"b92f",x"3d8b",x"372b",x"26c2",x"3bfe",x"24a2",x"3bc6",x"3a27"),
(x"b8ff",x"3d8a",x"3710",x"257a",x"3bff",x"15bc",x"3bcb",x"3a14",x"b907",x"3d8a",x"3718",x"25bc",x"3bfe",x"2680",x"3bc9",x"3a17",x"b931",x"3d8b",x"3710",x"2418",x"3bff",x"1a24",x"3bcb",x"3a28"),
(x"b912",x"3d45",x"373c",x"184d",x"bbff",x"26c2",x"3a57",x"3a57",x"b924",x"3d45",x"3749",x"1ef6",x"bbff",x"23ef",x"3a5a",x"3a5e",x"b918",x"3d45",x"374b",x"2511",x"bbff",x"2259",x"3a5a",x"3a5a"),
(x"b90c",x"3d45",x"3724",x"9e3f",x"bbff",x"a00b",x"3a53",x"3a55",x"b92b",x"3d45",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a55",x"3a61",x"b912",x"3d45",x"373c",x"184d",x"bbff",x"26c2",x"3a57",x"3a57"),
(x"b906",x"3d45",x"3710",x"2546",x"bbff",x"9624",x"3a4f",x"3a53",x"b931",x"3d45",x"3710",x"9edc",x"bc00",x"9da1",x"3a4f",x"3a63",x"b90c",x"3d45",x"3724",x"9e3f",x"bbff",x"a00b",x"3a53",x"3a55"),
(x"b1fd",x"3d56",x"3710",x"375d",x"bb1a",x"0000",x"3a6a",x"3b8f",x"b1fd",x"3d56",x"36da",x"35da",x"bb72",x"8000",x"3a5f",x"3b8f",x"b22d",x"3d55",x"3710",x"2c28",x"bbfb",x"0000",x"3a6a",x"3b94"),
(x"b6fb",x"3d54",x"3710",x"37ed",x"3af2",x"0000",x"3a3e",x"39d2",x"b6fb",x"3d54",x"36da",x"38e1",x"3a57",x"0000",x"3a33",x"39d2",x"b6ef",x"3d51",x"3710",x"3b57",x"3658",x"868d",x"3a3e",x"39d5"),
(x"b63d",x"3d74",x"3710",x"affc",x"3bf0",x"0000",x"3a32",x"3b80",x"b63d",x"3d74",x"36da",x"ab45",x"3bfc",x"0000",x"3a3d",x"3b80",x"b62a",x"3d74",x"3710",x"2fbb",x"3bf1",x"0000",x"3a32",x"3b7d"),
(x"b1c1",x"3d5b",x"3710",x"3680",x"bb4f",x"8000",x"3a6a",x"3b88",x"b1c1",x"3d5b",x"36da",x"37bd",x"bb00",x"0000",x"3a5f",x"3b88",x"b1fd",x"3d56",x"3710",x"375d",x"bb1a",x"0000",x"3a6a",x"3b8f"),
(x"b906",x"3d45",x"3710",x"2546",x"bbff",x"9624",x"3a4f",x"3a53",x"b906",x"3d45",x"36da",x"224c",x"bbff",x"0000",x"3a44",x"3a53",x"b931",x"3d45",x"3710",x"9edc",x"bc00",x"9da1",x"3a4f",x"3a63"),
(x"b721",x"3d59",x"3710",x"37a6",x"3b06",x"8000",x"3a3e",x"39ca",x"b721",x"3d59",x"36da",x"3711",x"3b2d",x"0000",x"3a33",x"39ca",x"b6fb",x"3d54",x"3710",x"37ed",x"3af2",x"0000",x"3a3e",x"39d2"),
(x"b575",x"3d83",x"3710",x"ba67",x"b8cb",x"868d",x"3a32",x"3b4e",x"b575",x"3d83",x"36da",x"bb59",x"b650",x"8000",x"3a3d",x"3b4e",x"b575",x"3d86",x"3710",x"bb97",x"350d",x"8000",x"3a32",x"3b4c"),
(x"b1a1",x"3d5c",x"3710",x"2ede",x"bbf4",x"0000",x"3a6a",x"3b85",x"b1a1",x"3d5c",x"36da",x"314f",x"bbe3",x"0000",x"3a5f",x"3b85",x"b1c1",x"3d5b",x"3710",x"3680",x"bb4f",x"8000",x"3a6a",x"3b88"),
(x"b72e",x"3d5b",x"3710",x"3b4f",x"367e",x"0000",x"3a3e",x"39c7",x"b72e",x"3d5b",x"36da",x"39a7",x"39a9",x"0000",x"3a33",x"39c7",x"b721",x"3d59",x"3710",x"37a6",x"3b06",x"8000",x"3a3e",x"39ca"),
(x"b62a",x"3d74",x"3710",x"2fbb",x"3bf1",x"0000",x"3a32",x"3b7d",x"b62a",x"3d74",x"36da",x"303b",x"3bed",x"8000",x"3a3d",x"3b7d",x"b5ce",x"3d71",x"3710",x"2f26",x"3bf3",x"0000",x"3a32",x"3b6a"),
(x"b161",x"3d5d",x"3710",x"3407",x"bbbd",x"8000",x"3a6a",x"3b7f",x"b161",x"3d5d",x"36da",x"30d8",x"bbe8",x"8000",x"3a5f",x"3b7f",x"b1a1",x"3d5c",x"3710",x"2ede",x"bbf4",x"0000",x"3a6a",x"3b85"),
(x"b72d",x"3d5d",x"3710",x"3778",x"bb13",x"0000",x"3a3e",x"39c5",x"b72d",x"3d5d",x"36da",x"3a45",x"b8f8",x"0000",x"3a33",x"39c5",x"b72e",x"3d5b",x"3710",x"3b4f",x"367e",x"0000",x"3a3e",x"39c7"),
(x"b5ce",x"3d71",x"3710",x"2f26",x"3bf3",x"0000",x"3a32",x"3b6a",x"b5ce",x"3d71",x"36da",x"2ae9",x"3bfc",x"8000",x"3a3d",x"3b6a",x"b5bd",x"3d71",x"3710",x"b559",x"3b8a",x"0000",x"3a32",x"3b67"),
(x"b135",x"3d5f",x"3710",x"3934",x"ba13",x"0000",x"3a6a",x"3b7b",x"b135",x"3d5f",x"36da",x"3822",x"bad9",x"8000",x"3a5f",x"3b7b",x"b161",x"3d5d",x"3710",x"3407",x"bbbd",x"8000",x"3a6a",x"3b7f"),
(x"b721",x"3d5e",x"3710",x"0cea",x"bc00",x"0000",x"3a17",x"3b9a",x"b721",x"3d5e",x"36da",x"2560",x"bbff",x"8000",x"3a0c",x"3b9a",x"b72d",x"3d5d",x"3710",x"3778",x"bb13",x"0000",x"3a17",x"3b9c"),
(x"b5bd",x"3d71",x"3710",x"b559",x"3b8a",x"0000",x"3a32",x"3b67",x"b5bd",x"3d71",x"36da",x"b6e1",x"3b38",x"0000",x"3a3d",x"3b67",x"b5a1",x"3d75",x"3710",x"b72c",x"3b26",x"8000",x"3a32",x"3b60"),
(x"b93a",x"3d73",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"383f",x"b93a",x"3d73",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"3838",x"b931",x"3d74",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3842"),
(x"b116",x"3d64",x"3710",x"3bdf",x"b1b0",x"068d",x"3a6a",x"3b76",x"b116",x"3d64",x"36da",x"3b51",x"b675",x"8000",x"3a5f",x"3b76",x"b135",x"3d5f",x"3710",x"3934",x"ba13",x"0000",x"3a6a",x"3b7b"),
(x"b568",x"3d46",x"3710",x"b810",x"bae4",x"0000",x"3a17",x"3b39",x"b568",x"3d46",x"36da",x"b919",x"ba29",x"0000",x"3a0c",x"3b39",x"b575",x"3d4a",x"3710",x"bab5",x"b85c",x"0000",x"3a17",x"3b3c"),
(x"b5a1",x"3d75",x"3710",x"b72c",x"3b26",x"8000",x"3a32",x"3b60",x"b5a1",x"3d75",x"36da",x"b67b",x"3b50",x"0000",x"3a3d",x"3b60",x"b581",x"3d78",x"3710",x"b794",x"3b0b",x"0000",x"3a32",x"3b5a"),
(x"b669",x"3d5d",x"3710",x"abaa",x"bbfc",x"0000",x"3a17",x"3b77",x"b669",x"3d5d",x"36da",x"a65f",x"bbff",x"0000",x"3a0c",x"3b77",x"b721",x"3d5e",x"3710",x"0cea",x"bc00",x"0000",x"3a17",x"3b9a"),
(x"b581",x"3d78",x"3710",x"b794",x"3b0b",x"0000",x"3a32",x"3b5a",x"b581",x"3d78",x"36da",x"b89f",x"3a87",x"0000",x"3a3d",x"3b5a",x"b568",x"3d7e",x"3710",x"b9f3",x"3958",x"0000",x"3a32",x"3b53"),
(x"b8a3",x"3d47",x"3710",x"2a1e",x"bbfd",x"0000",x"3a4f",x"3a2e",x"b8a3",x"3d47",x"36da",x"2850",x"bbfe",x"8000",x"3a44",x"3a2e",x"b906",x"3d45",x"3710",x"2546",x"bbff",x"9624",x"3a4f",x"3a53"),
(x"b63d",x"3d5c",x"3710",x"ab45",x"bbfc",x"0000",x"3a17",x"3b6e",x"b63d",x"3d5c",x"36da",x"affc",x"bbf0",x"8000",x"3a0c",x"3b6e",x"b669",x"3d5d",x"3710",x"abaa",x"bbfc",x"0000",x"3a17",x"3b77"),
(x"b568",x"3d89",x"3710",x"b919",x"3a29",x"0000",x"3a32",x"3b48",x"b568",x"3d89",x"36da",x"b810",x"3ae4",x"8000",x"3a3d",x"3b48",x"b558",x"3d8b",x"3710",x"b3cc",x"3bc2",x"8000",x"3a32",x"3b44"),
(x"b62a",x"3d5c",x"3710",x"303b",x"bbed",x"0000",x"3a17",x"3b6b",x"b62a",x"3d5c",x"36da",x"2fb9",x"bbf1",x"0000",x"3a0c",x"3b6b",x"b63d",x"3d5c",x"3710",x"ab45",x"bbfc",x"0000",x"3a17",x"3b6e"),
(x"b558",x"3d8b",x"3710",x"b3cc",x"3bc2",x"8000",x"3a32",x"3b44",x"b558",x"3d8b",x"36da",x"b02d",x"3bee",x"0000",x"3a3d",x"3b44",x"b544",x"3d8b",x"3710",x"b138",x"3be4",x"0000",x"3a32",x"3b40"),
(x"b575",x"3d4a",x"3710",x"bab5",x"b85c",x"0000",x"3a17",x"3b3c",x"b575",x"3d4a",x"36da",x"bb97",x"b50d",x"8000",x"3a0c",x"3b3c",x"b575",x"3d4c",x"3710",x"bb59",x"3650",x"8000",x"3a17",x"3b3e"),
(x"b544",x"3d8b",x"3710",x"b138",x"3be4",x"0000",x"3a32",x"3b40",x"b544",x"3d8b",x"36da",x"b46b",x"3bb0",x"0000",x"3a3d",x"3b40",x"b52b",x"3d8d",x"3710",x"b472",x"3baf",x"0000",x"3a32",x"3b3b"),
(x"b5ce",x"3d5f",x"3710",x"2ae9",x"bbfc",x"0000",x"3a17",x"3b59",x"b5ce",x"3d5f",x"36da",x"2f26",x"bbf3",x"0000",x"3a0c",x"3b59",x"b62a",x"3d5c",x"3710",x"303b",x"bbed",x"0000",x"3a17",x"3b6b"),
(x"b52b",x"3d8d",x"3710",x"b472",x"3baf",x"0000",x"3a32",x"3b3b",x"b52b",x"3d8d",x"36da",x"b238",x"3bd8",x"8000",x"3a3d",x"3b3b",x"b50d",x"3d8e",x"3710",x"253f",x"3bff",x"0000",x"3a32",x"3b35"),
(x"b5bd",x"3d5e",x"3710",x"b6e1",x"bb38",x"0000",x"3a17",x"3b56",x"b5bd",x"3d5e",x"36da",x"b559",x"bb8a",x"0000",x"3a0c",x"3b56",x"b5ce",x"3d5f",x"3710",x"2ae9",x"bbfc",x"0000",x"3a17",x"3b59"),
(x"b50d",x"3d8e",x"3710",x"253f",x"3bff",x"0000",x"3a32",x"3b35",x"b50d",x"3d8e",x"36da",x"324a",x"3bd8",x"8000",x"3a3d",x"3b35",x"b4f9",x"3d8c",x"3710",x"38a5",x"3a82",x"0000",x"3a32",x"3b31"),
(x"b5a1",x"3d5a",x"3710",x"b67b",x"bb50",x"8000",x"3a17",x"3b50",x"b5a1",x"3d5a",x"36da",x"b72c",x"bb26",x"8000",x"3a0c",x"3b50",x"b5bd",x"3d5e",x"3710",x"b6e1",x"bb38",x"0000",x"3a17",x"3b56"),
(x"b4f9",x"3d8c",x"3710",x"38a5",x"3a82",x"0000",x"3a32",x"3b31",x"b4f9",x"3d8c",x"36da",x"3a57",x"38e0",x"8000",x"3a3d",x"3b31",x"b4f5",x"3d89",x"3710",x"3bbb",x"341b",x"8000",x"3a32",x"3b2e"),
(x"b581",x"3d57",x"3710",x"b89f",x"ba87",x"0000",x"3a17",x"3b4a",x"b581",x"3d57",x"36da",x"b794",x"bb0b",x"0000",x"3a0c",x"3b4a",x"b5a1",x"3d5a",x"3710",x"b67b",x"bb50",x"8000",x"3a17",x"3b50"),
(x"b4f5",x"3d89",x"3710",x"3bbb",x"341b",x"8000",x"3a32",x"3b2e",x"b4f5",x"3d89",x"36da",x"3bc4",x"33a2",x"0000",x"3a3d",x"3b2e",x"b4f2",x"3d86",x"3710",x"3aea",x"3805",x"8000",x"3a32",x"3b2c"),
(x"b931",x"3d74",x"3710",x"bbea",x"a7ae",x"307d",x"3a5b",x"33c4",x"b931",x"3d74",x"36da",x"bbff",x"a4d0",x"0000",x"3a5a",x"33f3",x"b931",x"3d8b",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a6f",x"33c9"),
(x"b8ff",x"3d8a",x"3710",x"257a",x"3bff",x"15bc",x"3bcb",x"3a14",x"b8ff",x"3d8a",x"36da",x"26a7",x"3bff",x"8000",x"3bd5",x"3a14",x"b8a3",x"3d89",x"3710",x"286a",x"3bfe",x"8000",x"3bcb",x"39f0"),
(x"b568",x"3d51",x"3710",x"bb03",x"b7b2",x"0000",x"3a17",x"3b43",x"b568",x"3d51",x"36da",x"b9f3",x"b958",x"0000",x"3a0c",x"3b43",x"b581",x"3d57",x"3710",x"b89f",x"ba87",x"0000",x"3a17",x"3b4a"),
(x"b4f2",x"3d86",x"3710",x"3aea",x"3805",x"8000",x"3a32",x"3b2c",x"b4f2",x"3d86",x"36da",x"3a46",x"38f6",x"0000",x"3a3d",x"3b2c",x"b4da",x"3d7f",x"3710",x"3a4b",x"38ef",x"068d",x"3a32",x"3b25"),
(x"b8a3",x"3d89",x"3710",x"286a",x"3bfe",x"8000",x"3bcb",x"39f0",x"b8a3",x"3d89",x"36da",x"2a59",x"3bfd",x"0000",x"3bd5",x"39f0",x"b89e",x"3d88",x"3710",x"36f0",x"3b35",x"0000",x"3bcb",x"39ee"),
(x"b558",x"3d45",x"3710",x"b02d",x"bbee",x"0000",x"3a17",x"3b35",x"b558",x"3d45",x"36da",x"b3cc",x"bbc2",x"8000",x"3a0c",x"3b35",x"b568",x"3d46",x"3710",x"b810",x"bae4",x"0000",x"3a17",x"3b39"),
(x"b4da",x"3d7f",x"3710",x"3a4b",x"38ef",x"068d",x"3a32",x"3b25",x"b4da",x"3d7f",x"36da",x"3afc",x"37cc",x"0000",x"3a3d",x"3b25",x"b4d8",x"3d7c",x"3710",x"3be5",x"b11d",x"068d",x"3a32",x"3b22"),
(x"b89e",x"3d88",x"3710",x"36f0",x"3b35",x"0000",x"3bcb",x"39ee",x"b89e",x"3d88",x"36da",x"380f",x"3ae4",x"0000",x"3bd5",x"39ee",x"b88f",x"3d84",x"3710",x"380a",x"3ae7",x"0000",x"3bcb",x"39e7"),
(x"b544",x"3d45",x"3710",x"b46b",x"bbb0",x"0000",x"3a17",x"3b31",x"b544",x"3d45",x"36da",x"b138",x"bbe4",x"0000",x"3a0c",x"3b31",x"b558",x"3d45",x"3710",x"b02d",x"bbee",x"0000",x"3a17",x"3b35"),
(x"b4d8",x"3d7c",x"3710",x"3be5",x"b11d",x"068d",x"3a32",x"3b22",x"b4d8",x"3d7c",x"36da",x"3af9",x"b7d7",x"068d",x"3a3d",x"3b22",x"b4e1",x"3d7a",x"3710",x"3599",x"bb7e",x"0000",x"3a32",x"3b20"),
(x"b88f",x"3d84",x"3710",x"380a",x"3ae7",x"0000",x"3bcb",x"39e7",x"b88f",x"3d84",x"36da",x"377a",x"3b12",x"0000",x"3bd5",x"39e7",x"b87d",x"3d7f",x"3710",x"3541",x"3b8e",x"0000",x"3bcb",x"39df"),
(x"b52b",x"3d42",x"3710",x"b238",x"bbd8",x"8000",x"3a17",x"3b2c",x"b52b",x"3d42",x"36da",x"b472",x"bbaf",x"0000",x"3a0c",x"3b2c",x"b544",x"3d45",x"3710",x"b46b",x"bbb0",x"0000",x"3a17",x"3b31"),
(x"b4e1",x"3d7a",x"3710",x"3599",x"bb7e",x"0000",x"3a32",x"3b20",x"b4e1",x"3d7a",x"36da",x"33d2",x"bbc1",x"8000",x"3a3d",x"3b20",x"b51a",x"3d77",x"3710",x"332b",x"bbcb",x"8000",x"3a32",x"3b14"),
(x"b87d",x"3d7f",x"3710",x"3541",x"3b8e",x"0000",x"3bcb",x"39df",x"b87d",x"3d7f",x"36da",x"3244",x"3bd8",x"0000",x"3bd5",x"39df",x"b86e",x"3d7f",x"3710",x"ad01",x"3bf9",x"0000",x"3bcb",x"39d8"),
(x"b50d",x"3d41",x"3710",x"324a",x"bbd8",x"8000",x"3a17",x"3b27",x"b50d",x"3d41",x"36da",x"253f",x"bbff",x"068d",x"3a0c",x"3b27",x"b52b",x"3d42",x"3710",x"b238",x"bbd8",x"8000",x"3a17",x"3b2c"),
(x"b51a",x"3d77",x"3710",x"332b",x"bbcb",x"8000",x"3a32",x"3b14",x"b51a",x"3d77",x"36da",x"347c",x"bbad",x"0000",x"3a3d",x"3b14",x"b528",x"3d75",x"3710",x"37fe",x"baed",x"0000",x"3a32",x"3b11"),
(x"b86e",x"3d7f",x"3710",x"ad01",x"3bf9",x"0000",x"3bcb",x"39d8",x"b86e",x"3d7f",x"36da",x"b406",x"3bbe",x"0000",x"3bd5",x"39d8",x"b867",x"3d81",x"3710",x"b975",x"39d9",x"0000",x"3bcb",x"39d5"),
(x"b4f9",x"3d43",x"3710",x"3a57",x"b8e0",x"0000",x"3a17",x"3b22",x"b4f9",x"3d43",x"36da",x"38a5",x"ba82",x"8000",x"3a0c",x"3b22",x"b50d",x"3d41",x"3710",x"324a",x"bbd8",x"8000",x"3a17",x"3b27"),
(x"b528",x"3d75",x"3710",x"37fe",x"baed",x"0000",x"3a32",x"3b11",x"b528",x"3d75",x"36da",x"38ed",x"ba4d",x"8000",x"3a3d",x"3b11",x"b52c",x"3d74",x"3710",x"3bfc",x"ab6c",x"0000",x"3a32",x"3b10"),
(x"b867",x"3d81",x"3710",x"b975",x"39d9",x"0000",x"3bcb",x"39d5",x"b867",x"3d81",x"36da",x"baa2",x"3877",x"0000",x"3bd5",x"39d5",x"b865",x"3d84",x"3710",x"bb0e",x"378a",x"8000",x"3bcb",x"39d3"),
(x"b4f5",x"3d47",x"3710",x"3bc4",x"b3a2",x"8000",x"3a17",x"3b20",x"b4f5",x"3d47",x"36da",x"3bbb",x"b41b",x"8000",x"3a0c",x"3b20",x"b4f9",x"3d43",x"3710",x"3a57",x"b8e0",x"0000",x"3a17",x"3b22"),
(x"b52c",x"3d74",x"3710",x"3bfc",x"ab6c",x"0000",x"3b11",x"39ae",x"b52c",x"3d74",x"36da",x"3b0d",x"378c",x"0000",x"3b06",x"39ae",x"b526",x"3d73",x"3710",x"35f8",x"3b6b",x"0000",x"3b11",x"39af"),
(x"b865",x"3d84",x"3710",x"bb0e",x"378a",x"8000",x"3bcb",x"39d3",x"b865",x"3d84",x"36da",x"baaf",x"3865",x"8000",x"3bd5",x"39d3",x"b85e",x"3d88",x"3710",x"b878",x"3aa2",x"0000",x"3bcb",x"39ce"),
(x"b4f2",x"3d4a",x"3710",x"3a46",x"b8f6",x"0000",x"3a17",x"3b1d",x"b4f2",x"3d4a",x"36da",x"3aea",x"b805",x"8000",x"3a0c",x"3b1d",x"b4f5",x"3d47",x"3710",x"3bc4",x"b3a2",x"8000",x"3a17",x"3b20"),
(x"b526",x"3d73",x"3710",x"35f8",x"3b6b",x"0000",x"3b11",x"39af",x"b526",x"3d73",x"36da",x"33bb",x"3bc3",x"0000",x"3b06",x"39af",x"b50c",x"3d72",x"3710",x"292b",x"3bfe",x"8000",x"3b11",x"39b4"),
(x"b116",x"3d6c",x"3710",x"3b51",x"3675",x"0000",x"3a6a",x"3b70",x"b116",x"3d6c",x"36da",x"3bdf",x"31b0",x"868d",x"3a5f",x"3b70",x"b116",x"3d64",x"3710",x"3bdf",x"b1b0",x"068d",x"3a6a",x"3b76"),
(x"b85e",x"3d88",x"3710",x"b878",x"3aa2",x"0000",x"3bcb",x"39ce",x"b85e",x"3d88",x"36da",x"b5f3",x"3b6d",x"068d",x"3bd5",x"39ce",x"b84a",x"3d8b",x"3710",x"ac15",x"3bfb",x"8000",x"3bcb",x"39c6"),
(x"b4da",x"3d51",x"3710",x"3afc",x"b7cc",x"8000",x"3a17",x"3b17",x"b4da",x"3d51",x"36da",x"3a4b",x"b8ef",x"8000",x"3a0c",x"3b17",x"b4f2",x"3d4a",x"3710",x"3a46",x"b8f6",x"0000",x"3a17",x"3b1d"),
(x"b451",x"3d72",x"3710",x"a0ea",x"3c00",x"0000",x"3b11",x"39d8",x"b451",x"3d72",x"36da",x"a987",x"3bfe",x"8000",x"3b06",x"39d8",x"b441",x"3d73",x"3710",x"b6f3",x"3b34",x"0000",x"3b11",x"39db"),
(x"b89e",x"3d47",x"3710",x"380f",x"bae4",x"0000",x"3a4f",x"3a2c",x"b89e",x"3d47",x"36da",x"36f0",x"bb35",x"0000",x"3a44",x"3a2c",x"b8a3",x"3d47",x"3710",x"2a1e",x"bbfd",x"0000",x"3a4f",x"3a2e"),
(x"b84a",x"3d8b",x"3710",x"ac15",x"3bfb",x"8000",x"3bcb",x"39c6",x"b84a",x"3d8b",x"36da",x"30e0",x"3be8",x"8000",x"3bd5",x"39c6",x"b83a",x"3d88",x"3710",x"3890",x"3a92",x"0000",x"3bcb",x"39bf"),
(x"b4d8",x"3d54",x"3710",x"3af9",x"37d7",x"868d",x"3a17",x"3b14",x"b4d8",x"3d54",x"36da",x"3be5",x"311d",x"068d",x"3a0c",x"3b14",x"b4da",x"3d51",x"3710",x"3afc",x"b7cc",x"8000",x"3a17",x"3b17"),
(x"b50c",x"3d72",x"3710",x"292b",x"3bfe",x"8000",x"3b11",x"39b4",x"b50c",x"3d72",x"36da",x"236c",x"3bff",x"0000",x"3b06",x"39b4",x"b451",x"3d72",x"3710",x"a0ea",x"3c00",x"0000",x"3b11",x"39d8"),
(x"b88f",x"3d4c",x"3710",x"377a",x"bb12",x"8000",x"3a4f",x"3a25",x"b88f",x"3d4c",x"36da",x"380a",x"bae7",x"0000",x"3a44",x"3a25",x"b89e",x"3d47",x"3710",x"380f",x"bae4",x"0000",x"3a4f",x"3a2c"),
(x"b568",x"3d7e",x"3710",x"b9f3",x"3958",x"0000",x"3a32",x"3b53",x"b568",x"3d7e",x"36da",x"bb03",x"37b2",x"868d",x"3a3d",x"3b53",x"b569",x"3d80",x"3710",x"bb2d",x"b70f",x"0000",x"3a32",x"3b51"),
(x"b4e1",x"3d56",x"3710",x"33d2",x"3bc1",x"868d",x"3a17",x"3b12",x"b4e1",x"3d56",x"36da",x"3599",x"3b7e",x"0000",x"3a0c",x"3b12",x"b4d8",x"3d54",x"3710",x"3af9",x"37d7",x"868d",x"3a17",x"3b14"),
(x"b441",x"3d73",x"3710",x"b6f3",x"3b34",x"0000",x"3b11",x"39db",x"b441",x"3d73",x"36da",x"b7a3",x"3b07",x"0000",x"3b06",x"39db",x"b40d",x"3d7a",x"3710",x"b83a",x"3aca",x"0000",x"3b11",x"39e6"),
(x"b87d",x"3d50",x"3710",x"3244",x"bbd8",x"0000",x"3a4f",x"3a1d",x"b87d",x"3d50",x"36da",x"3541",x"bb8e",x"0000",x"3a44",x"3a1d",x"b88f",x"3d4c",x"3710",x"377a",x"bb12",x"8000",x"3a4f",x"3a25"),
(x"b83a",x"3d88",x"3710",x"3890",x"3a92",x"0000",x"3bcb",x"39bf",x"b83a",x"3d88",x"36da",x"3953",x"39f7",x"8000",x"3bd5",x"39bf",x"b820",x"3d7a",x"3710",x"391f",x"3a25",x"0000",x"3bcb",x"39b0"),
(x"b51a",x"3d58",x"3710",x"347c",x"3bad",x"8000",x"3a17",x"3b07",x"b51a",x"3d58",x"36da",x"332b",x"3bcb",x"0000",x"3a0c",x"3b07",x"b4e1",x"3d56",x"3710",x"33d2",x"3bc1",x"868d",x"3a17",x"3b12"),
(x"b40d",x"3d7a",x"3710",x"b83a",x"3aca",x"0000",x"3b11",x"39e6",x"b40d",x"3d7a",x"36da",x"b8bf",x"3a70",x"068d",x"3b06",x"39e6",x"b407",x"3d7d",x"3710",x"bb61",x"3629",x"0000",x"3b11",x"39e8"),
(x"b86e",x"3d51",x"3710",x"b406",x"bbbe",x"0000",x"3a4f",x"3a17",x"b86e",x"3d51",x"36da",x"ad01",x"bbf9",x"0000",x"3a44",x"3a17",x"b87d",x"3d50",x"3710",x"3244",x"bbd8",x"0000",x"3a4f",x"3a1d"),
(x"b569",x"3d80",x"3710",x"bb2d",x"b70f",x"0000",x"3a32",x"3b51",x"b569",x"3d80",x"36da",x"ba4b",x"b8f0",x"0000",x"3a3d",x"3b51",x"b575",x"3d83",x"3710",x"ba67",x"b8cb",x"868d",x"3a32",x"3b4e"),
(x"b528",x"3d5a",x"3710",x"38ed",x"3a4d",x"0000",x"3a17",x"3b04",x"b528",x"3d5a",x"36da",x"37fe",x"3aed",x"0000",x"3a0c",x"3b04",x"b51a",x"3d58",x"3710",x"347c",x"3bad",x"8000",x"3a17",x"3b07"),
(x"b407",x"3d7d",x"3710",x"bb61",x"3629",x"0000",x"3b11",x"39e8",x"b407",x"3d7d",x"36da",x"bbf7",x"2ddb",x"0000",x"3b06",x"39e8",x"b409",x"3d7e",x"3710",x"bb1a",x"b75c",x"8000",x"3b11",x"39e9"),
(x"b867",x"3d4f",x"3710",x"baa2",x"b877",x"0000",x"3a4f",x"3a15",x"b867",x"3d4f",x"36da",x"b975",x"b9d8",x"0000",x"3a44",x"3a15",x"b86e",x"3d51",x"3710",x"b406",x"bbbe",x"0000",x"3a4f",x"3a17"),
(x"b820",x"3d7a",x"3710",x"391f",x"3a25",x"0000",x"3bcb",x"39b0",x"b820",x"3d7a",x"36da",x"385c",x"3ab4",x"0000",x"3bd5",x"39b0",x"b801",x"3d73",x"3710",x"3561",x"3b88",x"0000",x"3bcb",x"39a3"),
(x"b52c",x"3d5b",x"3710",x"3b0d",x"b78c",x"0000",x"3a17",x"3b03",x"b52c",x"3d5b",x"36da",x"3bfc",x"2b6c",x"0000",x"3a0c",x"3b03",x"b528",x"3d5a",x"3710",x"38ed",x"3a4d",x"0000",x"3a17",x"3b04"),
(x"b409",x"3d7e",x"3710",x"bb1a",x"b75c",x"8000",x"3b11",x"39e9",x"b409",x"3d7e",x"36da",x"bab5",x"b85b",x"0000",x"3b06",x"39e9",x"b413",x"3d82",x"3710",x"bb08",x"b7a0",x"0000",x"3b11",x"39ed"),
(x"b865",x"3d4c",x"3710",x"baaf",x"b865",x"8000",x"3a4f",x"3a12",x"b865",x"3d4c",x"36da",x"bb0e",x"b78a",x"8000",x"3a44",x"3a12",x"b867",x"3d4f",x"3710",x"baa2",x"b877",x"0000",x"3a4f",x"3a15"),
(x"b801",x"3d73",x"3710",x"3561",x"3b88",x"0000",x"3bcb",x"39a3",x"b801",x"3d73",x"36da",x"3346",x"3bca",x"0000",x"3bd5",x"39a3",x"b7c0",x"3d71",x"3710",x"29e3",x"3bfd",x"0000",x"3bcb",x"3996"),
(x"b526",x"3d5d",x"3710",x"33bc",x"bbc3",x"0000",x"3a23",x"3a1a",x"b526",x"3d5d",x"36da",x"35f9",x"bb6b",x"0000",x"3a18",x"3a1a",x"b52c",x"3d5b",x"3710",x"3b0d",x"b78c",x"0000",x"3a23",x"3a1b"),
(x"b413",x"3d82",x"3710",x"bb08",x"b7a0",x"0000",x"3b11",x"39ed",x"b413",x"3d82",x"36da",x"bba9",x"b499",x"0000",x"3b06",x"39ed",x"b413",x"3d84",x"3710",x"bb8c",x"354a",x"8000",x"3b11",x"39ee"),
(x"b85e",x"3d47",x"3710",x"b5f3",x"bb6d",x"8000",x"3a4f",x"3a0e",x"b85e",x"3d47",x"36da",x"b878",x"baa2",x"0000",x"3a44",x"3a0e",x"b865",x"3d4c",x"3710",x"baaf",x"b865",x"8000",x"3a4f",x"3a12"),
(x"b7c0",x"3d71",x"3710",x"29e3",x"3bfd",x"0000",x"3bcb",x"3996",x"b7c0",x"3d71",x"36da",x"a984",x"3bfe",x"8000",x"3bd5",x"3996",x"b794",x"3d73",x"3710",x"b358",x"3bc9",x"0000",x"3bcb",x"398d"),
(x"b50c",x"3d5e",x"3710",x"236c",x"bbff",x"0000",x"3a23",x"3a15",x"b50c",x"3d5e",x"36da",x"292b",x"bbfe",x"8000",x"3a18",x"3a15",x"b526",x"3d5d",x"3710",x"33bc",x"bbc3",x"0000",x"3a23",x"3a1a"),
(x"b413",x"3d84",x"3710",x"bb8c",x"354a",x"8000",x"3b11",x"39ee",x"b413",x"3d84",x"36da",x"ba12",x"3935",x"868d",x"3b06",x"39ee",x"b40b",x"3d85",x"3710",x"b3aa",x"3bc4",x"8000",x"3b11",x"39f0"),
(x"b84a",x"3d45",x"3710",x"30e0",x"bbe8",x"8000",x"3a4f",x"3a06",x"b84a",x"3d45",x"36da",x"ac15",x"bbfb",x"868d",x"3a44",x"3a06",x"b85e",x"3d47",x"3710",x"b5f3",x"bb6d",x"8000",x"3a4f",x"3a0e"),
(x"b794",x"3d73",x"3710",x"b358",x"3bc9",x"0000",x"3bcb",x"398d",x"b794",x"3d73",x"36da",x"b51c",x"3b94",x"0000",x"3bd5",x"398d",x"b77a",x"3d76",x"3710",x"b83f",x"3ac7",x"0000",x"3bcb",x"3987"),
(x"b441",x"3d5d",x"3710",x"b7a3",x"bb07",x"0000",x"3a23",x"39ee",x"b441",x"3d5d",x"36da",x"b6f3",x"bb34",x"0000",x"3a18",x"39ee",x"b451",x"3d5e",x"3710",x"a987",x"bbfe",x"8000",x"3a23",x"39f1"),
(x"b40b",x"3d85",x"3710",x"b3aa",x"3bc4",x"8000",x"3b11",x"39f0",x"b40b",x"3d85",x"36da",x"aabe",x"3bfd",x"868d",x"3b06",x"39f0",x"b3f4",x"3d85",x"3710",x"3149",x"3be3",x"0000",x"3b11",x"39f3"),
(x"b83a",x"3d48",x"3710",x"3953",x"b9f7",x"8000",x"3a4f",x"39ff",x"b83a",x"3d48",x"36da",x"3890",x"ba92",x"0000",x"3a44",x"39ff",x"b84a",x"3d45",x"3710",x"30e0",x"bbe8",x"8000",x"3a4f",x"3a06"),
(x"b77a",x"3d76",x"3710",x"b83f",x"3ac7",x"0000",x"3bcb",x"3987",x"b77a",x"3d76",x"36da",x"b97c",x"39d2",x"0000",x"3bd5",x"3987",x"b776",x"3d78",x"3710",x"bbee",x"3037",x"0000",x"3bcb",x"3985"),
(x"b451",x"3d5e",x"3710",x"a987",x"bbfe",x"8000",x"3a23",x"39f1",x"b451",x"3d5e",x"36da",x"a0ea",x"bc00",x"0000",x"3a18",x"39f1",x"b50c",x"3d5e",x"3710",x"236c",x"bbff",x"0000",x"3a23",x"3a15"),
(x"b3f4",x"3d85",x"3710",x"3149",x"3be3",x"0000",x"3b11",x"39f3",x"b3f4",x"3d85",x"36da",x"3408",x"3bbd",x"0000",x"3b06",x"39f3",x"b3d2",x"3d83",x"3710",x"2ffb",x"3bf0",x"0000",x"3b11",x"39f7"),
(x"b569",x"3d4f",x"3710",x"ba4b",x"38f0",x"0000",x"3a17",x"3b41",x"b569",x"3d4f",x"36da",x"bb2d",x"370f",x"0000",x"3a0c",x"3b41",x"b568",x"3d51",x"3710",x"bb03",x"b7b2",x"0000",x"3a17",x"3b43"),
(x"b776",x"3d78",x"3710",x"bbee",x"3037",x"0000",x"3bcb",x"3985",x"b776",x"3d78",x"36da",x"bbce",x"b2fb",x"0000",x"3bd5",x"3985",x"b77b",x"3d7a",x"3710",x"b937",x"ba10",x"0000",x"3bcb",x"3983"),
(x"b40d",x"3d55",x"3710",x"b8bf",x"ba70",x"8000",x"3a23",x"39e3",x"b40d",x"3d55",x"36da",x"b83a",x"baca",x"0000",x"3a18",x"39e3",x"b441",x"3d5d",x"3710",x"b7a3",x"bb07",x"0000",x"3a23",x"39ee"),
(x"b3d2",x"3d83",x"3710",x"2ffb",x"3bf0",x"0000",x"3b11",x"39f7",x"b3d2",x"3d83",x"36da",x"abf9",x"3bfc",x"0000",x"3b06",x"39f7",x"b3a5",x"3d85",x"3710",x"24fd",x"3bff",x"0000",x"3b11",x"39fb"),
(x"b820",x"3d55",x"3710",x"385c",x"bab4",x"8000",x"3a4f",x"39f1",x"b820",x"3d55",x"36da",x"391f",x"ba25",x"0000",x"3a44",x"39f1",x"b83a",x"3d48",x"3710",x"3953",x"b9f7",x"8000",x"3a4f",x"39ff"),
(x"b77b",x"3d7a",x"3710",x"b937",x"ba10",x"0000",x"3a9e",x"3ac5",x"b77b",x"3d7a",x"36da",x"b853",x"baba",x"0000",x"3a93",x"3ac5",x"b790",x"3d7d",x"3710",x"b606",x"bb69",x"0000",x"3a9e",x"3ac9"),
(x"b407",x"3d53",x"3710",x"bbf7",x"addb",x"0000",x"3a23",x"39e1",x"b407",x"3d53",x"36da",x"bb61",x"b629",x"0000",x"3a18",x"39e1",x"b40d",x"3d55",x"3710",x"b8bf",x"ba70",x"8000",x"3a23",x"39e3"),
(x"b3a5",x"3d85",x"3710",x"24fd",x"3bff",x"0000",x"3b11",x"39fb",x"b3a5",x"3d85",x"36da",x"32b6",x"3bd2",x"0000",x"3b06",x"39fb",x"b368",x"3d82",x"3710",x"37ea",x"3af3",x"8000",x"3b11",x"3a01"),
(x"b575",x"3d4c",x"3710",x"bb59",x"3650",x"8000",x"3a17",x"3b3e",x"b575",x"3d4c",x"36da",x"ba67",x"38cb",x"068d",x"3a0c",x"3b3e",x"b569",x"3d4f",x"3710",x"ba4b",x"38f0",x"0000",x"3a17",x"3b41"),
(x"b790",x"3d7d",x"3710",x"b606",x"bb69",x"0000",x"3a9e",x"3ac9",x"b790",x"3d7d",x"36da",x"b461",x"bbb1",x"0000",x"3a93",x"3ac9",x"b7a8",x"3d7e",x"3710",x"b360",x"bbc8",x"0000",x"3a9e",x"3ace"),
(x"b409",x"3d51",x"3710",x"bab5",x"385b",x"0000",x"3a23",x"39e0",x"b409",x"3d51",x"36da",x"bb1a",x"375d",x"0000",x"3a18",x"39e0",x"b407",x"3d53",x"3710",x"bbf7",x"addb",x"0000",x"3a23",x"39e1"),
(x"b368",x"3d82",x"3710",x"37ea",x"3af3",x"8000",x"3b11",x"3a01",x"b368",x"3d82",x"36da",x"3912",x"3a2f",x"8000",x"3b06",x"3a01",x"b340",x"3d7c",x"3710",x"3aba",x"3853",x"0000",x"3b11",x"3a07"),
(x"b801",x"3d5d",x"3710",x"3346",x"bbca",x"0000",x"3a4f",x"39e4",x"b801",x"3d5d",x"36da",x"3561",x"bb88",x"0000",x"3a44",x"39e4",x"b820",x"3d55",x"3710",x"385c",x"bab4",x"8000",x"3a4f",x"39f1"),
(x"b7a8",x"3d7e",x"3710",x"b360",x"bbc8",x"0000",x"3a9e",x"3ace",x"b7a8",x"3d7e",x"36da",x"b4b8",x"bba4",x"8000",x"3a93",x"3ace",x"b7bd",x"3d80",x"3710",x"b6d2",x"bb3c",x"0000",x"3a9e",x"3ad2"),
(x"b413",x"3d4e",x"3710",x"bba9",x"3498",x"0000",x"3a23",x"39dc",x"b413",x"3d4e",x"36da",x"bb08",x"37a1",x"068d",x"3a18",x"39dc",x"b409",x"3d51",x"3710",x"bab5",x"385b",x"0000",x"3a23",x"39e0"),
(x"b340",x"3d7c",x"3710",x"3aba",x"3853",x"0000",x"3b11",x"3a07",x"b340",x"3d7c",x"36da",x"3b6b",x"35fb",x"8000",x"3b06",x"3a07",x"b33a",x"3d77",x"3710",x"3bf6",x"ae02",x"868d",x"3b11",x"3a0b"),
(x"b7c0",x"3d5f",x"3710",x"a984",x"bbfe",x"0000",x"3a4f",x"39d8",x"b7c0",x"3d5f",x"36da",x"29e3",x"bbfd",x"0000",x"3a44",x"39d8",x"b801",x"3d5d",x"3710",x"3346",x"bbca",x"0000",x"3a4f",x"39e4"),
(x"b7bd",x"3d80",x"3710",x"b6d2",x"bb3c",x"0000",x"3a9e",x"3ad2",x"b7bd",x"3d80",x"36da",x"b821",x"bada",x"8000",x"3a93",x"3ad2",x"b7c7",x"3d82",x"3710",x"ba01",x"b948",x"8a8d",x"3a9e",x"3ad5"),
(x"b931",x"3d45",x"3710",x"bbe9",x"26a1",x"309e",x"3a36",x"33ca",x"b931",x"3d45",x"36da",x"bbff",x"26b5",x"0000",x"3a38",x"33fa",x"b930",x"3d5c",x"3710",x"bbeb",x"2604",x"3075",x"3a49",x"33c0"),
(x"b413",x"3d4c",x"3710",x"ba12",x"b935",x"868d",x"3a23",x"39db",x"b413",x"3d4c",x"36da",x"bb8c",x"b54a",x"8000",x"3a18",x"39db",x"b413",x"3d4e",x"3710",x"bba9",x"3498",x"0000",x"3a23",x"39dc"),
(x"b33a",x"3d77",x"3710",x"3bf6",x"ae02",x"868d",x"3b11",x"3a0b",x"b33a",x"3d77",x"36da",x"3b88",x"b564",x"8000",x"3b06",x"3a0b",x"b351",x"3d72",x"3710",x"3b23",x"b738",x"0000",x"3b11",x"3a0f"),
(x"b794",x"3d5d",x"3710",x"b51c",x"bb94",x"0000",x"3a4f",x"39cf",x"b794",x"3d5d",x"36da",x"b358",x"bbc9",x"0000",x"3a44",x"39cf",x"b7c0",x"3d5f",x"3710",x"a984",x"bbfe",x"0000",x"3a4f",x"39d8"),
(x"b7c7",x"3d82",x"3710",x"ba01",x"b948",x"8a8d",x"3a9e",x"3ad5",x"b7c7",x"3d82",x"36da",x"bb43",x"b6b4",x"0000",x"3a93",x"3ad5",x"b7c7",x"3d84",x"3710",x"b8b7",x"3a76",x"0000",x"3a9e",x"3ad6"),
(x"b40b",x"3d4b",x"3710",x"aabe",x"bbfd",x"068d",x"3a23",x"39d9",x"b40b",x"3d4b",x"36da",x"b3aa",x"bbc4",x"0000",x"3a18",x"39d9",x"b413",x"3d4c",x"3710",x"ba12",x"b935",x"868d",x"3a23",x"39db"),
(x"b351",x"3d72",x"3710",x"3b23",x"b738",x"0000",x"3b11",x"3a0f",x"b351",x"3d72",x"36da",x"3bb2",x"b458",x"0000",x"3b06",x"3a0f",x"b34f",x"3d70",x"3710",x"3913",x"3a2f",x"0000",x"3b11",x"3a11"),
(x"b77a",x"3d5a",x"3710",x"b97c",x"b9d2",x"0000",x"3a4f",x"39ca",x"b77a",x"3d5a",x"36da",x"b83f",x"bac7",x"0000",x"3a44",x"39ca",x"b794",x"3d5d",x"3710",x"b51c",x"bb94",x"0000",x"3a4f",x"39cf"),
(x"b7c7",x"3d84",x"3710",x"b8b7",x"3a76",x"0000",x"3a9e",x"3ad6",x"b7c7",x"3d84",x"36da",x"b744",x"3b20",x"8a8d",x"3a93",x"3ad6",x"b7a4",x"3d87",x"3710",x"b654",x"3b58",x"0000",x"3a9e",x"3add"),
(x"b3f4",x"3d4b",x"3710",x"3408",x"bbbd",x"0000",x"3a23",x"39d6",x"b3f4",x"3d4b",x"36da",x"3149",x"bbe3",x"0000",x"3a18",x"39d6",x"b40b",x"3d4b",x"3710",x"aabe",x"bbfd",x"068d",x"3a23",x"39d9"),
(x"b34f",x"3d70",x"3710",x"3913",x"3a2f",x"0000",x"3a6a",x"3b35",x"b34f",x"3d70",x"36da",x"3448",x"3bb5",x"0000",x"3a5f",x"3b35",x"b326",x"3d70",x"3710",x"a5e3",x"3bff",x"0000",x"3a6a",x"3b39"),
(x"b776",x"3d57",x"3710",x"bbce",x"32fb",x"0000",x"3a3e",x"3a17",x"b776",x"3d57",x"36da",x"bbee",x"b037",x"0000",x"3a33",x"3a17",x"b77a",x"3d5a",x"3710",x"b97c",x"b9d2",x"0000",x"3a3e",x"3a19"),
(x"b7a4",x"3d87",x"3710",x"b654",x"3b58",x"0000",x"3a9e",x"3add",x"b7a4",x"3d87",x"36da",x"b64a",x"3b5a",x"8000",x"3a93",x"3add",x"b783",x"3d8b",x"3710",x"b33d",x"3bca",x"0000",x"3a9e",x"3ae4"),
(x"b3d2",x"3d4c",x"3710",x"abf9",x"bbfc",x"8000",x"3a23",x"39d2",x"b3d2",x"3d4c",x"36da",x"2ffb",x"bbf0",x"0000",x"3a18",x"39d2",x"b3f4",x"3d4b",x"3710",x"3408",x"bbbd",x"0000",x"3a23",x"39d6"),
(x"b326",x"3d70",x"3710",x"a5e3",x"3bff",x"0000",x"3a6a",x"3b39",x"b326",x"3d70",x"36da",x"ad8e",x"3bf8",x"0000",x"3a5f",x"3b39",x"b2d6",x"3d71",x"3710",x"b287",x"3bd4",x"0000",x"3a6a",x"3b40"),
(x"b77b",x"3d55",x"3710",x"b853",x"3aba",x"0000",x"3a3e",x"3a15",x"b77b",x"3d55",x"36da",x"b937",x"3a10",x"8000",x"3a33",x"3a15",x"b776",x"3d57",x"3710",x"bbce",x"32fb",x"0000",x"3a3e",x"3a17"),
(x"b783",x"3d8b",x"3710",x"b33d",x"3bca",x"0000",x"3a9e",x"3ae4",x"b783",x"3d8b",x"36da",x"afa0",x"3bf1",x"0000",x"3a93",x"3ae4",x"b73e",x"3d8c",x"3710",x"27ae",x"3bfe",x"0000",x"3a9e",x"3af1"),
(x"b3a5",x"3d4b",x"3710",x"32b6",x"bbd2",x"868d",x"3a23",x"39ce",x"b3a5",x"3d4b",x"36da",x"2504",x"bbff",x"0000",x"3a18",x"39ce",x"b3d2",x"3d4c",x"3710",x"abf9",x"bbfc",x"8000",x"3a23",x"39d2"),
(x"b2d6",x"3d71",x"3710",x"b287",x"3bd4",x"0000",x"3a6a",x"3b40",x"b2d6",x"3d71",x"36da",x"b4dc",x"3b9f",x"0000",x"3a5f",x"3b40",x"b2aa",x"3d74",x"3710",x"b78b",x"3b0e",x"0000",x"3a6a",x"3b45"),
(x"b790",x"3d52",x"3710",x"b461",x"3bb1",x"0000",x"3a3e",x"3a11",x"b790",x"3d52",x"36da",x"b606",x"3b69",x"0000",x"3a33",x"3a11",x"b77b",x"3d55",x"3710",x"b853",x"3aba",x"0000",x"3a3e",x"3a15"),
(x"b73e",x"3d8c",x"3710",x"27ae",x"3bfe",x"0000",x"3a9e",x"3af1",x"b73e",x"3d8c",x"36da",x"2f57",x"3bf2",x"8000",x"3a93",x"3af1",x"b705",x"3d89",x"3710",x"34b8",x"3ba4",x"0000",x"3a9e",x"3afc"),
(x"b368",x"3d4e",x"3710",x"3912",x"ba2f",x"8000",x"3a23",x"39c8",x"b368",x"3d4e",x"36da",x"37ea",x"baf3",x"8000",x"3a18",x"39c8",x"b3a5",x"3d4b",x"3710",x"32b6",x"bbd2",x"868d",x"3a23",x"39ce"),
(x"b2aa",x"3d74",x"3710",x"b78b",x"3b0e",x"0000",x"3a6a",x"3b45",x"b2aa",x"3d74",x"36da",x"b7e2",x"3af5",x"0000",x"3a5f",x"3b45",x"b261",x"3d79",x"3710",x"b72e",x"3b26",x"8000",x"3a6a",x"3b4d"),
(x"b7a8",x"3d51",x"3710",x"b4b8",x"3ba4",x"8000",x"3a3e",x"3a0c",x"b7a8",x"3d51",x"36da",x"b360",x"3bc8",x"8000",x"3a33",x"3a0c",x"b790",x"3d52",x"3710",x"b461",x"3bb1",x"0000",x"3a3e",x"3a11"),
(x"b705",x"3d89",x"3710",x"34b8",x"3ba4",x"0000",x"3a9e",x"3afc",x"b705",x"3d89",x"36da",x"36ee",x"3b35",x"0000",x"3a93",x"3afc",x"b6f1",x"3d84",x"3710",x"3a69",x"38c9",x"068d",x"3a9e",x"3b01"),
(x"b340",x"3d54",x"3710",x"3b6b",x"b5fb",x"0000",x"3a23",x"39c2",x"b340",x"3d54",x"36da",x"3aba",x"b853",x"8000",x"3a18",x"39c2",x"b368",x"3d4e",x"3710",x"3912",x"ba2f",x"8000",x"3a23",x"39c8"),
(x"b261",x"3d79",x"3710",x"b72e",x"3b26",x"8000",x"3a6a",x"3b4d",x"b261",x"3d79",x"36da",x"b5e0",x"3b70",x"8000",x"3a5f",x"3b4d",x"b22d",x"3d7b",x"3710",x"ae88",x"3bf5",x"0000",x"3a6a",x"3b52"),
(x"b7bd",x"3d4f",x"3710",x"b821",x"3ad9",x"0000",x"3a3e",x"3a08",x"b7bd",x"3d4f",x"36da",x"b6d2",x"3b3c",x"0000",x"3a33",x"3a08",x"b7a8",x"3d51",x"3710",x"b4b8",x"3ba4",x"8000",x"3a3e",x"3a0c"),
(x"b6f1",x"3d84",x"3710",x"3a69",x"38c9",x"068d",x"3a9e",x"3b01",x"b6f1",x"3d84",x"36da",x"3b73",x"35d3",x"8000",x"3a93",x"3b01",x"b6ef",x"3d7f",x"3710",x"3be9",x"b0b7",x"0000",x"3a9e",x"3b05"),
(x"b33a",x"3d59",x"3710",x"3b88",x"3564",x"868d",x"3a23",x"39be",x"b33a",x"3d59",x"36da",x"3bf6",x"2e02",x"8000",x"3a18",x"39be",x"b340",x"3d54",x"3710",x"3b6b",x"b5fb",x"0000",x"3a23",x"39c2"),
(x"b22d",x"3d7b",x"3710",x"ae88",x"3bf5",x"0000",x"3a6a",x"3b52",x"b22d",x"3d7b",x"36da",x"2c28",x"3bfb",x"0000",x"3a5f",x"3b52",x"b1fd",x"3d79",x"3710",x"35da",x"3b72",x"0000",x"3a6a",x"3b57"),
(x"b7c7",x"3d4d",x"3710",x"bb43",x"36b4",x"0000",x"3a3e",x"3a06",x"b7c7",x"3d4d",x"36da",x"ba01",x"3948",x"8000",x"3a33",x"3a06",x"b7bd",x"3d4f",x"3710",x"b821",x"3ad9",x"0000",x"3a3e",x"3a08"),
(x"b6ef",x"3d7f",x"3710",x"3be9",x"b0b7",x"0000",x"3a9e",x"3b05",x"b6ef",x"3d7f",x"36da",x"3b57",x"b658",x"8000",x"3a93",x"3b05",x"b6fb",x"3d7b",x"3710",x"38e1",x"ba57",x"0000",x"3a9e",x"3b08"),
(x"b351",x"3d5d",x"3710",x"3bb2",x"3458",x"8000",x"3a23",x"39ba",x"b351",x"3d5d",x"36da",x"3b23",x"3738",x"0000",x"3a18",x"39ba",x"b33a",x"3d59",x"3710",x"3b88",x"3564",x"868d",x"3a23",x"39be"),
(x"b1fd",x"3d79",x"3710",x"35da",x"3b72",x"0000",x"3a6a",x"3b57",x"b1fd",x"3d79",x"36da",x"375d",x"3b1a",x"8000",x"3a5f",x"3b57",x"b1c1",x"3d75",x"3710",x"37bc",x"3b00",x"0000",x"3a6a",x"3b5d"),
(x"b7c7",x"3d4c",x"3710",x"b744",x"bb20",x"0000",x"3a3e",x"3a05",x"b7c7",x"3d4c",x"36da",x"b8b7",x"ba76",x"0000",x"3a33",x"3a05",x"b7c7",x"3d4d",x"3710",x"bb43",x"36b4",x"0000",x"3a3e",x"3a06"),
(x"b6fb",x"3d7b",x"3710",x"38e1",x"ba57",x"0000",x"3a9e",x"3b08",x"b6fb",x"3d7b",x"36da",x"37ed",x"baf2",x"868d",x"3a93",x"3b08",x"b721",x"3d77",x"3710",x"3711",x"bb2d",x"0000",x"3a9e",x"3b10"),
(x"b34f",x"3d60",x"3710",x"3448",x"bbb5",x"0000",x"3a23",x"39b8",x"b34f",x"3d60",x"36da",x"3913",x"ba2f",x"0000",x"3a18",x"39b8",x"b351",x"3d5d",x"3710",x"3bb2",x"3458",x"8000",x"3a23",x"39ba"),
(x"b1c1",x"3d75",x"3710",x"37bc",x"3b00",x"0000",x"3a6a",x"3b5d",x"b1c1",x"3d75",x"36da",x"367f",x"3b4f",x"8000",x"3a5f",x"3b5d",x"b1a1",x"3d73",x"3710",x"314f",x"3be3",x"8000",x"3a6a",x"3b60"),
(x"b7a4",x"3d48",x"3710",x"b64a",x"bb5a",x"0000",x"3a3e",x"39fd",x"b7a4",x"3d48",x"36da",x"b654",x"bb58",x"8000",x"3a33",x"39fd",x"b7c7",x"3d4c",x"3710",x"b744",x"bb20",x"0000",x"3a3e",x"3a05"),
(x"b721",x"3d77",x"3710",x"3711",x"bb2d",x"0000",x"3a9e",x"3b10",x"b721",x"3d77",x"36da",x"37a6",x"bb06",x"0000",x"3a93",x"3b10",x"b72e",x"3d75",x"3710",x"39a7",x"b9a8",x"0000",x"3a9e",x"3b13"),
(x"b326",x"3d60",x"3710",x"ad8e",x"bbf8",x"0000",x"3a6a",x"3bad",x"b326",x"3d60",x"36da",x"a5e3",x"bbff",x"0000",x"3a5f",x"3bad",x"b34f",x"3d60",x"3710",x"3448",x"bbb5",x"0000",x"3a6a",x"3bb1"),
(x"b1a1",x"3d73",x"3710",x"314f",x"3be3",x"8000",x"3a6a",x"3b60",x"b1a1",x"3d73",x"36da",x"2ede",x"3bf4",x"0000",x"3a5f",x"3b60",x"b161",x"3d73",x"3710",x"30d8",x"3be8",x"8000",x"3a6a",x"3b66"),
(x"b783",x"3d45",x"3710",x"afa0",x"bbf1",x"0000",x"3a3e",x"39f7",x"b783",x"3d45",x"36da",x"b33d",x"bbca",x"8000",x"3a33",x"39f7",x"b7a4",x"3d48",x"3710",x"b64a",x"bb5a",x"0000",x"3a3e",x"39fd"),
(x"b72e",x"3d75",x"3710",x"39a7",x"b9a8",x"0000",x"3a32",x"3bb1",x"b72e",x"3d75",x"36da",x"3b4f",x"b67e",x"8000",x"3a3d",x"3bb1",x"b72d",x"3d73",x"3710",x"3a45",x"38f8",x"0000",x"3a32",x"3bb0"),
(x"b2d6",x"3d5f",x"3710",x"b4dc",x"bb9f",x"0000",x"3a6a",x"3ba5",x"b2d6",x"3d5f",x"36da",x"b287",x"bbd4",x"0000",x"3a5f",x"3ba5",x"b326",x"3d60",x"3710",x"ad8e",x"bbf8",x"0000",x"3a6a",x"3bad"),
(x"b161",x"3d73",x"3710",x"30d8",x"3be8",x"8000",x"3a6a",x"3b66",x"b161",x"3d73",x"36da",x"3408",x"3bbd",x"0000",x"3a5f",x"3b66",x"b135",x"3d71",x"3710",x"3822",x"3ad9",x"0000",x"3a6a",x"3b6b"),
(x"b73e",x"3d44",x"3710",x"2f57",x"bbf2",x"0000",x"3a3e",x"39ea",x"b73e",x"3d44",x"36da",x"27ae",x"bbff",x"0000",x"3a33",x"39ea",x"b783",x"3d45",x"3710",x"afa0",x"bbf1",x"0000",x"3a3e",x"39f7"),
(x"b72d",x"3d73",x"3710",x"3a45",x"38f8",x"0000",x"3a32",x"3bb0",x"b72d",x"3d73",x"36da",x"3778",x"3b13",x"0000",x"3a3d",x"3bb0",x"b721",x"3d72",x"3710",x"2560",x"3bff",x"0000",x"3a32",x"3bad"),
(x"b2aa",x"3d5c",x"3710",x"b7e2",x"baf5",x"0000",x"3a6a",x"3ba1",x"b2aa",x"3d5c",x"36da",x"b78b",x"bb0e",x"0000",x"3a5f",x"3ba1",x"b2d6",x"3d5f",x"3710",x"b4dc",x"bb9f",x"0000",x"3a6a",x"3ba5"),
(x"b135",x"3d71",x"3710",x"3822",x"3ad9",x"0000",x"3a6a",x"3b6b",x"b135",x"3d71",x"36da",x"3934",x"3a13",x"8000",x"3a5f",x"3b6b",x"b116",x"3d6c",x"3710",x"3b51",x"3675",x"0000",x"3a6a",x"3b70"),
(x"b705",x"3d47",x"3710",x"36ee",x"bb35",x"0000",x"3a3e",x"39de",x"b705",x"3d47",x"36da",x"34b8",x"bba4",x"868d",x"3a33",x"39de",x"b73e",x"3d44",x"3710",x"2f57",x"bbf2",x"0000",x"3a3e",x"39ea"),
(x"b575",x"3d86",x"3710",x"bb97",x"350d",x"8000",x"3a32",x"3b4c",x"b575",x"3d86",x"36da",x"bab5",x"385c",x"068d",x"3a3d",x"3b4c",x"b568",x"3d89",x"3710",x"b919",x"3a29",x"0000",x"3a32",x"3b48"),
(x"b938",x"3d5e",x"3710",x"bbc9",x"a82f",x"3347",x"3beb",x"398f",x"b938",x"3d5e",x"36da",x"bbfe",x"a8f0",x"0000",x"3bea",x"3999",x"b93a",x"3d73",x"3710",x"bbf8",x"a8ed",x"2cf9",x"3bfb",x"398f"),
(x"b261",x"3d57",x"3710",x"b5e0",x"bb70",x"8000",x"3a6a",x"3b99",x"b261",x"3d57",x"36da",x"b72e",x"bb26",x"0000",x"3a5f",x"3b99",x"b2aa",x"3d5c",x"3710",x"b7e2",x"baf5",x"0000",x"3a6a",x"3ba1"),
(x"b931",x"3d8b",x"3710",x"2418",x"3bff",x"1a24",x"3bcb",x"3a28",x"b931",x"3d8b",x"36da",x"23ae",x"3bff",x"0000",x"3bd5",x"3a28",x"b8ff",x"3d8a",x"3710",x"257a",x"3bff",x"15bc",x"3bcb",x"3a14"),
(x"b6f1",x"3d4b",x"3710",x"3b73",x"b5d3",x"0000",x"3a3e",x"39d9",x"b6f1",x"3d4b",x"36da",x"3a69",x"b8c9",x"8000",x"3a33",x"39d9",x"b705",x"3d47",x"3710",x"36ee",x"bb35",x"0000",x"3a3e",x"39de"),
(x"b721",x"3d72",x"3710",x"2560",x"3bff",x"0000",x"3a32",x"3bad",x"b721",x"3d72",x"36da",x"0cea",x"3c00",x"0000",x"3a3d",x"3bad",x"b669",x"3d72",x"3710",x"a666",x"3bff",x"0000",x"3a32",x"3b89"),
(x"b22d",x"3d55",x"3710",x"2c28",x"bbfb",x"0000",x"3a6a",x"3b94",x"b22d",x"3d55",x"36da",x"ae8a",x"bbf5",x"8000",x"3a5f",x"3b94",x"b261",x"3d57",x"3710",x"b5e0",x"bb70",x"8000",x"3a6a",x"3b99"),
(x"b6ef",x"3d51",x"3710",x"3b57",x"3658",x"868d",x"3a3e",x"39d5",x"b6ef",x"3d51",x"36da",x"3be9",x"30b7",x"068d",x"3a33",x"39d5",x"b6f1",x"3d4b",x"3710",x"3b73",x"b5d3",x"0000",x"3a3e",x"39d9"),
(x"b669",x"3d72",x"3710",x"a666",x"3bff",x"0000",x"3a32",x"3b89",x"b669",x"3d72",x"36da",x"abae",x"3bfc",x"8000",x"3a3d",x"3b89",x"b63d",x"3d74",x"3710",x"affc",x"3bf0",x"0000",x"3a32",x"3b80"),
(x"b930",x"3d5c",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bbd",x"39bd",x"b930",x"3d5c",x"36da",x"b67a",x"bb50",x"0000",x"3bc3",x"39b4",x"b938",x"3d5e",x"3710",x"b678",x"bb4d",x"2af3",x"3bba",x"39ba"),
(x"b930",x"4041",x"3710",x"bbeb",x"2604",x"3075",x"39c5",x"33c0",x"b92a",x"4041",x"3733",x"bb1e",x"2518",x"3748",x"39c4",x"339f",x"b92b",x"4036",x"3732",x"bb64",x"243f",x"361b",x"39b1",x"33aa"),
(x"b92a",x"4041",x"3733",x"bb1e",x"2518",x"3748",x"39c4",x"339f",x"b922",x"4041",x"3748",x"b86c",x"29d9",x"3aa7",x"39c4",x"3388",x"b924",x"4036",x"3749",x"ba3b",x"2680",x"3902",x"39b0",x"3392"),
(x"b922",x"4041",x"3748",x"b86c",x"29d9",x"3aa7",x"39c4",x"3388",x"b91b",x"4041",x"3749",x"3594",x"2b76",x"3b7b",x"39c3",x"337b",x"b91f",x"4036",x"374e",x"ac96",x"29b2",x"3bf8",x"39b0",x"3387"),
(x"b91b",x"4041",x"3749",x"3594",x"2b76",x"3b7b",x"39c3",x"337b",x"b913",x"4041",x"373b",x"3aa1",x"2559",x"3879",x"39c3",x"3369",x"b918",x"4036",x"374b",x"38f0",x"29d6",x"3a48",x"39b0",x"337b"),
(x"b913",x"4041",x"373b",x"381d",x"3a67",x"34eb",x"3b1c",x"3899",x"b913",x"4042",x"373a",x"3ae3",x"2b4b",x"380a",x"3b1b",x"3899",x"b90e",x"4042",x"370e",x"3754",x"3ae5",x"32eb",x"3b1f",x"38a1"),
(x"b913",x"4042",x"373a",x"3ae3",x"2b4b",x"380a",x"3b1b",x"3899",x"b913",x"4041",x"373b",x"381d",x"3a67",x"34eb",x"3b1c",x"3899",x"b91b",x"4041",x"3749",x"382b",x"a439",x"3ad3",x"3b1a",x"3895"),
(x"b913",x"4042",x"373a",x"3b64",x"a9cc",x"3612",x"3beb",x"39a8",x"b913",x"404d",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"39a7",x"b90f",x"404d",x"3727",x"3bc1",x"a907",x"33c0",x"3bfb",x"39a3"),
(x"b90f",x"404d",x"3727",x"3bc1",x"a907",x"33c0",x"3bfb",x"39a3",x"b90e",x"4042",x"370e",x"3bcb",x"a949",x"330f",x"3bea",x"399f",x"b913",x"4042",x"373a",x"3b64",x"a9cc",x"3612",x"3beb",x"39a8"),
(x"b913",x"404d",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"39a7",x"b913",x"4042",x"373a",x"3b64",x"a9cc",x"3612",x"3beb",x"39a8",x"b91b",x"4042",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"39ac"),
(x"b91a",x"404d",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"39ab",x"b91b",x"4042",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"39ac",x"b924",x"4043",x"374d",x"af62",x"aa90",x"3bef",x"3bec",x"39af"),
(x"b928",x"404d",x"374d",x"b867",x"a907",x"3aab",x"3bfc",x"39b1",x"b922",x"404d",x"3751",x"a111",x"aa52",x"3bfd",x"3bfc",x"39af",x"b924",x"4043",x"374d",x"af62",x"aa90",x"3bef",x"3bec",x"39af"),
(x"b92f",x"404d",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"39b5",x"b928",x"404d",x"374d",x"b867",x"a907",x"3aab",x"3bfc",x"39b1",x"b92b",x"4043",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"39b3"),
(x"b935",x"404d",x"3725",x"bb50",x"a63f",x"3678",x"3bfb",x"39ba",x"b92f",x"404d",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"39b5",x"b930",x"4043",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"39b6"),
(x"b930",x"4043",x"3738",x"b75b",x"bae5",x"32d3",x"3b16",x"388d",x"b92a",x"4041",x"3733",x"b800",x"ba99",x"3435",x"3b19",x"388d",x"b930",x"4041",x"3710",x"b700",x"bb23",x"2f0f",x"3b1b",x"3887"),
(x"b913",x"4041",x"373b",x"3aa1",x"2559",x"3879",x"39c3",x"3369",x"b90c",x"4036",x"3724",x"3af5",x"1a59",x"37e2",x"39b0",x"3352",x"b912",x"4036",x"373c",x"3aea",x"2832",x"3802",x"39b0",x"336a"),
(x"b913",x"4041",x"373b",x"3aa1",x"2559",x"3879",x"39c3",x"3369",x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e",x"b90c",x"4036",x"3724",x"3af5",x"1a59",x"37e2",x"39b0",x"3352"),
(x"b91b",x"4042",x"374a",x"3544",x"b37e",x"3b51",x"3b18",x"3896",x"b91b",x"4041",x"3749",x"382b",x"a439",x"3ad3",x"3b1a",x"3895",x"b922",x"4041",x"3748",x"b511",x"b92e",x"398b",x"3b18",x"3893"),
(x"b922",x"4041",x"3748",x"b511",x"b92e",x"398b",x"3b18",x"3893",x"b92a",x"4041",x"3733",x"b800",x"ba99",x"3435",x"3b19",x"388d",x"b92b",x"4043",x"3744",x"b779",x"ba1b",x"3724",x"3b16",x"388f"),
(x"b935",x"404d",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3821",x"b93a",x"404d",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"381d",x"b931",x"404d",x"3710",x"b3e2",x"3bbf",x"28bf",x"3b1e",x"3820"),
(x"b92f",x"404d",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3826",x"b935",x"404d",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3821",x"b92a",x"404d",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3827"),
(x"b928",x"404d",x"374d",x"b4d8",x"3aa1",x"3784",x"3b25",x"382a",x"b92f",x"404d",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3826",x"b925",x"404d",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"382b"),
(x"b91a",x"404d",x"374d",x"35fb",x"37c0",x"3a53",x"3b22",x"3830",x"b922",x"404d",x"3751",x"9ac2",x"39ac",x"39a3",x"3b24",x"382d",x"b920",x"404d",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"382d"),
(x"b913",x"404d",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3832",x"b91a",x"404d",x"374d",x"35fb",x"37c0",x"3a53",x"3b22",x"3830",x"b919",x"404e",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"382f"),
(x"b90f",x"404d",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3835",x"b913",x"404d",x"373e",x"3a5b",x"3408",x"386a",x"3b1f",x"3832",x"b913",x"404e",x"373e",x"3b0f",x"a05a",x"3786",x"3b1e",x"3831"),
(x"b90d",x"404d",x"3711",x"b36d",x"a40b",x"3bc7",x"39d6",x"3349",x"b906",x"404d",x"3713",x"29ab",x"208e",x"3bfd",x"39d7",x"333d",x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e"),
(x"b92f",x"4059",x"372b",x"bbac",x"a891",x"347c",x"39eb",x"33b1",x"b92a",x"404d",x"3739",x"bb13",x"a8dd",x"3771",x"39d7",x"339e",x"b931",x"404d",x"3710",x"bbea",x"a7ae",x"307d",x"39d7",x"33c4"),
(x"b92a",x"404d",x"3739",x"bb13",x"a8dd",x"3771",x"39d7",x"339e",x"b92c",x"4059",x"373a",x"baa5",x"a5fd",x"3872",x"39eb",x"33a3",x"b925",x"4059",x"3749",x"b926",x"a7c8",x"3a1d",x"39eb",x"3391"),
(x"b920",x"404d",x"374b",x"b451",x"a960",x"3bb2",x"39d8",x"3385",x"b925",x"404d",x"3746",x"b918",x"a84d",x"3a28",x"39d8",x"338e",x"b925",x"4059",x"3749",x"b926",x"a7c8",x"3a1d",x"39eb",x"3391"),
(x"b919",x"404e",x"3749",x"3647",x"a97a",x"3b59",x"39d8",x"3379",x"b920",x"404d",x"374b",x"b451",x"a960",x"3bb2",x"39d8",x"3385",x"b91f",x"4059",x"374f",x"a812",x"a959",x"3bfd",x"39eb",x"3384"),
(x"b913",x"404e",x"373e",x"3ac8",x"a7bb",x"383c",x"39d8",x"336a",x"b919",x"404e",x"3749",x"3647",x"a97a",x"3b59",x"39d8",x"3379",x"b918",x"4059",x"374b",x"38ec",x"a7f6",x"3a4c",x"39eb",x"3378"),
(x"b913",x"404e",x"373e",x"3ac8",x"a7bb",x"383c",x"39d8",x"336a",x"b911",x"4059",x"373c",x"3ac9",x"a6b5",x"383a",x"39eb",x"3366",x"b90b",x"4059",x"3722",x"3b0f",x"a82c",x"3781",x"39ea",x"334c"),
(x"b90b",x"404d",x"371c",x"3aa9",x"a818",x"386b",x"39d7",x"334a",x"b90b",x"4059",x"3722",x"3b0f",x"a82c",x"3781",x"39ea",x"334c",x"b907",x"4059",x"3718",x"38f7",x"a86d",x"3a44",x"39eb",x"3340"),
(x"b116",x"404a",x"3710",x"0000",x"8000",x"3c00",x"39d1",x"2450",x"b116",x"4045",x"3710",x"0000",x"8000",x"3c00",x"39c9",x"2450",x"b135",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"24c1"),
(x"b135",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"24c1",x"b161",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"255f",x"b161",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"255f"),
(x"b161",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"255f",x"b1a1",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2642",x"b1a1",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2642"),
(x"b1a1",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2642",x"b1a1",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2642",x"b1c1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"26b3"),
(x"b1c1",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"26b3",x"b1fd",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39be",x"278b",x"b1fd",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"278b"),
(x"b1fd",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"278b",x"b1fd",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39be",x"278b",x"b22d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"281a"),
(x"b22d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"281a",x"b22d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"281a",x"b261",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39be",x"2878"),
(x"b261",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dc",x"2878",x"b261",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39be",x"2878",x"b2aa",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"28fa"),
(x"b2aa",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"28fa",x"b2d6",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2949",x"b2d6",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2949"),
(x"b2d6",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2949",x"b2d6",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2949",x"b326",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"29d7"),
(x"b326",x"404b",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"29d7",x"b326",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"29d7",x"b34f",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2a20"),
(x"b50c",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2d8d",x"b50c",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2d8d",x"b451",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2c3f"),
(x"b451",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2c3f",x"b441",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2c23",x"b441",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2c23"),
(x"b441",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2c23",x"b441",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2c23",x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b"),
(x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b",x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b",x"b34f",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d4",x"2a20"),
(x"b40b",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2b83",x"b3f4",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2b47",x"b413",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2ba0"),
(x"b3f4",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2b47",x"b3d2",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"2b0a",x"b409",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2b7d"),
(x"b3d2",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"2b0a",x"b3a5",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2ab9",x"b407",x"4052",x"3710",x"0000",x"8000",x"3c00",x"39df",x"2b76"),
(x"b40b",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2b83",x"b413",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"2ba0",x"b413",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2ba0"),
(x"b3f4",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2b47",x"b413",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2ba0",x"b409",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2b7d"),
(x"b3d2",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2b0a",x"b409",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2b7d",x"b407",x"403d",x"3710",x"8000",x"0cea",x"3c00",x"39bb",x"2b76"),
(x"b3a5",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"2ab9",x"b407",x"403d",x"3710",x"8000",x"0cea",x"3c00",x"39bb",x"2b76",x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b"),
(x"b3a5",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2ab9",x"b368",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2a4d",x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b"),
(x"b368",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2a4d",x"b340",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"2a05",x"b351",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2a24"),
(x"b50c",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2d8d",x"b526",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2dbb",x"b526",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2dbb"),
(x"b62a",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2f8b",x"b62a",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2f8b",x"b5ce",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ee7"),
(x"b5ce",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ee7",x"b5bd",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ec9",x"b5bd",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2ec9"),
(x"b5bd",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"2ec9",x"b5bd",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"2ec9",x"b5a1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2e97"),
(x"b5a1",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2e97",x"b581",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"2e5e",x"b581",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"2e5e"),
(x"b581",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"2e5e",x"b581",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"2e5e",x"b568",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2e30"),
(x"b50d",x"405b",x"3710",x"0000",x"8000",x"3c00",x"39ee",x"2d8e",x"b4f9",x"405a",x"3710",x"0000",x"8000",x"3c00",x"39ec",x"2d6a",x"b4f5",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"2d63"),
(x"b52b",x"405a",x"3710",x"0000",x"8000",x"3c00",x"39ed",x"2dc4",x"b4f5",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"2d63",x"b4f2",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2d5e"),
(x"b4f5",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"2d63",x"b4f9",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ae",x"2d6a",x"b50d",x"4034",x"3710",x"0000",x"8000",x"3c00",x"39ac",x"2d8e"),
(x"b4f2",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2d5e",x"b4f5",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"2d63",x"b52b",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ad",x"2dc4"),
(x"b568",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b0",x"2e32",x"b575",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2e49",x"b575",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2e47"),
(x"b558",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2e14",x"b575",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"2e47",x"b569",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"2e33"),
(x"b568",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39ea",x"2e32",x"b558",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2e14",x"b575",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e4",x"2e47"),
(x"b558",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2e14",x"b544",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2df0",x"b569",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"2e33"),
(x"b4e1",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2d3f",x"b51a",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"2da6",x"b4da",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"2d33"),
(x"b4e1",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39be",x"2d3f",x"b4d8",x"403d",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"2d2f",x"b4da",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"2d33"),
(x"b51a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"2da6",x"b4da",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"2d33",x"b4f2",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b4",x"2d5e"),
(x"b51a",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"2da6",x"b528",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2dbf",x"b4f2",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e6",x"2d5e"),
(x"b528",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2dbf",x"b569",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"2e33",x"b544",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"2df0"),
(x"b544",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"2df0",x"b569",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"2e33",x"b528",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"2dbf"),
(x"b528",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"2dbf",x"b52c",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2dc5",x"b568",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"2e30"),
(x"b528",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"2dbf",x"b569",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"2e33",x"b568",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2e30"),
(x"b526",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2dbb",x"b52c",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2dc5",x"b52c",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2dc5"),
(x"b52c",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2dc5",x"b52c",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2dc5",x"b568",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"2e30"),
(x"b63d",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2fac",x"b62a",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d7",x"2f8b",x"b62a",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2f8b"),
(x"b669",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2ffc",x"b63d",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"2fac",x"b63d",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c3",x"2fac"),
(x"b721",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30a2",x"b669",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2ffc",x"b669",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"2ffc"),
(x"b721",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30a2",x"b721",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30a2",x"b72d",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30ad"),
(x"b794",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"3109",x"b7c0",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"3130",x"b7c0",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"3130"),
(x"b794",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"3109",x"b794",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"3109",x"b77a",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"30f1"),
(x"b77a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c1",x"30f1",x"b77a",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d9",x"30f1",x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed"),
(x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed",x"b72d",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30ad",x"b72d",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"30ad"),
(x"b6fb",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"3080",x"b6ef",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"3075",x"b6f1",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3076"),
(x"b721",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"30a2",x"b6fb",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"3080",x"b705",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3088"),
(x"b6f1",x"4056",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3076",x"b6ef",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"3075",x"b6fb",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"3080"),
(x"b705",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3088",x"b6fb",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"3080",x"b721",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"30a2"),
(x"b73e",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39ec",x"30bc",x"b721",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"30a2",x"b72e",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"30ae"),
(x"b72e",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"30ae",x"b721",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39c0",x"30a2",x"b73e",x"4035",x"3710",x"0000",x"8000",x"3c00",x"39ae",x"30bc"),
(x"b7c7",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3135",x"b7c7",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b6",x"3136",x"b7bd",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"312d"),
(x"b7c7",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3135",x"b7a4",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"3117",x"b7bd",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"312d"),
(x"b7a4",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"3117",x"b783",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"30f9",x"b7a8",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e0",x"311a"),
(x"b7a4",x"4038",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"3117",x"b7bd",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"312d",x"b7a8",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"311a"),
(x"b72e",x"4041",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"30ae",x"b77b",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"30f2",x"b776",x"403f",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"30ed"),
(x"b72e",x"404e",x"3710",x"0000",x"8000",x"3c00",x"39d8",x"30ae",x"b72d",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"30ad",x"b776",x"4050",x"3710",x"0000",x"8000",x"3c00",x"39db",x"30ed"),
(x"b801",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"316b",x"b7c0",x"404c",x"3710",x"0000",x"8000",x"3c00",x"39d5",x"3130",x"b7c0",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c5",x"3130"),
(x"b801",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"316b",x"b801",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c4",x"316b",x"b820",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"31a2"),
(x"b83a",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"31d0",x"b820",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"31a2",x"b820",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"31a2"),
(x"b84a",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"31ed",x"b83a",x"4057",x"3710",x"0000",x"8000",x"3c00",x"39e8",x"31d0",x"b83a",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b2",x"31d0"),
(x"b85e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3211",x"b84a",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"31ed",x"b84a",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"31ed"),
(x"b85e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3211",x"b85e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3211",x"b865",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"321d"),
(x"b867",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"3222",x"b865",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"321d",x"b865",x"4039",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"321d"),
(x"b867",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e2",x"3222",x"b867",x"403b",x"3710",x"0000",x"8000",x"3c00",x"39b8",x"3222",x"b86e",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"322d"),
(x"b87d",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"3248",x"b86e",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"322d",x"b86e",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"322d"),
(x"b88f",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3269",x"b87d",x"4053",x"3710",x"0000",x"8000",x"3c00",x"39e1",x"3248",x"b87d",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39b9",x"3248"),
(x"b88f",x"4055",x"3710",x"0000",x"8000",x"3c00",x"39e5",x"3269",x"b88f",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b5",x"3269",x"b89e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3284"),
(x"b8a3",x"4058",x"3710",x"2160",x"1cd0",x"3bff",x"39e9",x"328d",x"b89e",x"4058",x"3710",x"0000",x"8000",x"3c00",x"39e9",x"3284",x"b89e",x"4037",x"3710",x"0000",x"8000",x"3c00",x"39b1",x"3284"),
(x"b8a3",x"4058",x"3710",x"2160",x"1cd0",x"3bff",x"39e9",x"328d",x"b8a3",x"4037",x"3710",x"2081",x"9ea7",x"3bff",x"39b1",x"328d",x"b907",x"4042",x"3713",x"2c13",x"9f5f",x"3bfb",x"39c4",x"333e"),
(x"b8ff",x"4059",x"3710",x"2904",x"26d5",x"3bfd",x"39eb",x"3331",x"b8a3",x"4058",x"3710",x"2160",x"1cd0",x"3bff",x"39e9",x"328d",x"b906",x"404d",x"3713",x"29ab",x"208e",x"3bfd",x"39d7",x"333d"),
(x"b918",x"4059",x"374b",x"270a",x"3bfd",x"287a",x"3a18",x"3ba9",x"b91f",x"4059",x"374f",x"28f4",x"3bfa",x"ac2c",x"3a17",x"3bac",x"b925",x"4059",x"3749",x"257a",x"3bfd",x"28f7",x"3a18",x"3bae"),
(x"b911",x"4059",x"373c",x"2504",x"3bff",x"2111",x"3a1b",x"3ba6",x"b925",x"4059",x"3749",x"257a",x"3bfd",x"28f7",x"3a18",x"3bae",x"b92c",x"4059",x"373a",x"25e9",x"3bff",x"17c8",x"3a1b",x"3bb1"),
(x"b90b",x"4059",x"3722",x"2773",x"3bfe",x"22dc",x"3a1f",x"3ba4",x"b92c",x"4059",x"373a",x"25e9",x"3bff",x"17c8",x"3a1b",x"3bb1",x"b92f",x"4059",x"372b",x"26c2",x"3bfe",x"24a2",x"3a1e",x"3bb2"),
(x"b907",x"4059",x"3718",x"25bc",x"3bfe",x"2673",x"3a21",x"3ba2",x"b92f",x"4059",x"372b",x"26c2",x"3bfe",x"24a2",x"3a1e",x"3bb2",x"b931",x"4059",x"3710",x"2418",x"3bff",x"1a24",x"3a23",x"3bb3"),
(x"b924",x"4036",x"3749",x"1ef6",x"bbff",x"23ef",x"3a12",x"3bab",x"b91f",x"4036",x"374e",x"281b",x"bbe6",x"b0f0",x"3a13",x"3ba9",x"b918",x"4036",x"374b",x"2511",x"bbff",x"224c",x"3a12",x"3ba6"),
(x"b92b",x"4036",x"3732",x"9cd0",x"bc00",x"1bc8",x"3a0d",x"3bae",x"b924",x"4036",x"3749",x"1ef6",x"bbff",x"23ef",x"3a12",x"3bab",x"b912",x"4036",x"373c",x"184d",x"bbff",x"26c8",x"3a0f",x"3ba4"),
(x"b931",x"4036",x"3710",x"9ec2",x"bc00",x"9da1",x"3a07",x"3bb0",x"b92b",x"4036",x"3732",x"9cd0",x"bc00",x"1bc8",x"3a0d",x"3bae",x"b90c",x"4036",x"3724",x"9e3f",x"bbff",x"a025",x"3a0b",x"3ba2"),
(x"b1fd",x"403f",x"36da",x"35da",x"bb72",x"0000",x"3a50",x"3b8e",x"b22d",x"403e",x"36da",x"ae8a",x"bbf5",x"8000",x"3a50",x"3b93",x"b22d",x"403e",x"3710",x"2c28",x"bbfb",x"0000",x"3a5a",x"3b93"),
(x"b6fb",x"403e",x"36da",x"38e1",x"3a57",x"0000",x"3a72",x"3ad4",x"b6ef",x"403c",x"36da",x"3be9",x"30b7",x"868d",x"3a72",x"3ad8",x"b6ef",x"403c",x"3710",x"3b57",x"3658",x"8000",x"3a7c",x"3ad8"),
(x"b63d",x"404e",x"36da",x"ab45",x"3bfc",x"0000",x"3a8b",x"3b47",x"b62a",x"404d",x"36da",x"303b",x"3bed",x"8000",x"3a8b",x"3b4a",x"b62a",x"404d",x"3710",x"2fbb",x"3bf1",x"0000",x"3a96",x"3b4a"),
(x"b1c1",x"4041",x"36da",x"37bc",x"bb00",x"0000",x"3a50",x"3b87",x"b1fd",x"403f",x"36da",x"35da",x"bb72",x"0000",x"3a50",x"3b8e",x"b1fd",x"403f",x"3710",x"375d",x"bb1a",x"0000",x"3a5a",x"3b8e"),
(x"b906",x"4036",x"36da",x"2273",x"bbff",x"0000",x"39fd",x"3b9f",x"b931",x"4036",x"36da",x"9e3f",x"bc00",x"0000",x"39fd",x"3bb0",x"b931",x"4036",x"3710",x"9ec2",x"bc00",x"9da1",x"3a07",x"3bb0"),
(x"b721",x"4040",x"36da",x"3711",x"3b2d",x"0000",x"3a72",x"3acc",x"b6fb",x"403e",x"36da",x"38e1",x"3a57",x"0000",x"3a72",x"3ad4",x"b6fb",x"403e",x"3710",x"37ed",x"3af2",x"0000",x"3a7c",x"3ad4"),
(x"b575",x"4055",x"36da",x"bb59",x"b650",x"8000",x"3a8b",x"3b77",x"b575",x"4056",x"36da",x"bab5",x"385c",x"8000",x"3a8b",x"3b79",x"b575",x"4056",x"3710",x"bb97",x"350c",x"8000",x"3a96",x"3b79"),
(x"b1a1",x"4042",x"36da",x"314f",x"bbe3",x"0000",x"3a50",x"3b84",x"b1c1",x"4041",x"36da",x"37bc",x"bb00",x"0000",x"3a50",x"3b87",x"b1c1",x"4041",x"3710",x"367f",x"bb4f",x"0000",x"3a5a",x"3b87"),
(x"b72e",x"4041",x"36da",x"39a7",x"39a9",x"0000",x"3a72",x"3ac9",x"b721",x"4040",x"36da",x"3711",x"3b2d",x"0000",x"3a72",x"3acc",x"b721",x"4040",x"3710",x"37a6",x"3b06",x"8000",x"3a7c",x"3acc"),
(x"b62a",x"404d",x"36da",x"303b",x"3bed",x"8000",x"3a8b",x"3b4a",x"b5ce",x"404c",x"36da",x"2ae9",x"3bfc",x"8000",x"3a8b",x"3b5c",x"b5ce",x"404c",x"3710",x"2f26",x"3bf3",x"0000",x"3a96",x"3b5c"),
(x"b161",x"4042",x"36da",x"30d8",x"bbe8",x"8000",x"3a50",x"3b7e",x"b1a1",x"4042",x"36da",x"314f",x"bbe3",x"0000",x"3a50",x"3b84",x"b1a1",x"4042",x"3710",x"2ede",x"bbf4",x"0000",x"3a5a",x"3b84"),
(x"b72d",x"4042",x"36da",x"3a45",x"b8f8",x"0000",x"3a72",x"3ac8",x"b72e",x"4041",x"36da",x"39a7",x"39a9",x"0000",x"3a72",x"3ac9",x"b72e",x"4041",x"3710",x"3b4f",x"367e",x"8000",x"3a7c",x"3ac9"),
(x"b5ce",x"404c",x"36da",x"2ae9",x"3bfc",x"8000",x"3a8b",x"3b5c",x"b5bd",x"404c",x"36da",x"b6e1",x"3b38",x"0000",x"3a8b",x"3b5f",x"b5bd",x"404c",x"3710",x"b559",x"3b8a",x"0000",x"3a96",x"3b5f"),
(x"b135",x"4043",x"36da",x"3822",x"bad9",x"8000",x"3a50",x"3b7a",x"b161",x"4042",x"36da",x"30d8",x"bbe8",x"8000",x"3a50",x"3b7e",x"b161",x"4042",x"3710",x"3407",x"bbbd",x"8000",x"3a5a",x"3b7e"),
(x"b721",x"4042",x"36da",x"2560",x"bbff",x"8000",x"3a42",x"3bad",x"b72d",x"4042",x"36da",x"3a45",x"b8f8",x"0000",x"3a42",x"3bb0",x"b72d",x"4042",x"3710",x"3778",x"bb13",x"0000",x"3a4c",x"3bb0"),
(x"b5bd",x"404c",x"36da",x"b6e1",x"3b38",x"0000",x"3a8b",x"3b5f",x"b5a1",x"404e",x"36da",x"b67b",x"3b50",x"0000",x"3a8b",x"3b65",x"b5a1",x"404e",x"3710",x"b72d",x"3b26",x"8000",x"3a96",x"3b65"),
(x"b93a",x"404d",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"3816",x"b931",x"404d",x"36da",x"b311",x"3bcd",x"0000",x"3b16",x"3819",x"b931",x"404d",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3820"),
(x"b116",x"4045",x"36da",x"3b51",x"b675",x"8000",x"3a50",x"3b75",x"b135",x"4043",x"36da",x"3822",x"bad9",x"8000",x"3a50",x"3b7a",x"b135",x"4043",x"3710",x"3934",x"ba13",x"0000",x"3a5a",x"3b7a"),
(x"b568",x"4037",x"36da",x"b919",x"ba29",x"0000",x"3a42",x"3b48",x"b575",x"4038",x"36da",x"bb97",x"b50d",x"0000",x"3a42",x"3b4c",x"b575",x"4038",x"3710",x"bab5",x"b85c",x"8000",x"3a4c",x"3b4c"),
(x"b5a1",x"404e",x"36da",x"b67b",x"3b50",x"0000",x"3a8b",x"3b65",x"b581",x"4050",x"36da",x"b89f",x"3a87",x"0000",x"3a8b",x"3b6c",x"b581",x"4050",x"3710",x"b794",x"3b0b",x"0000",x"3a96",x"3b6c"),
(x"b669",x"4042",x"36da",x"a65f",x"bbff",x"0000",x"3a42",x"3b89",x"b721",x"4042",x"36da",x"2560",x"bbff",x"8000",x"3a42",x"3bad",x"b721",x"4042",x"3710",x"0cea",x"bc00",x"0000",x"3a4c",x"3bad"),
(x"b581",x"4050",x"36da",x"b89f",x"3a87",x"0000",x"3a8b",x"3b6c",x"b568",x"4053",x"36da",x"bb03",x"37b2",x"868d",x"3a8b",x"3b72",x"b568",x"4053",x"3710",x"b9f3",x"3958",x"0000",x"3a96",x"3b72"),
(x"b8a3",x"4037",x"36da",x"2850",x"bbfe",x"8000",x"39fd",x"3b78",x"b906",x"4036",x"36da",x"2273",x"bbff",x"0000",x"39fd",x"3b9f",x"b906",x"4036",x"3710",x"2546",x"bbff",x"9624",x"3a07",x"3b9f"),
(x"b63d",x"4041",x"36da",x"affc",x"bbf0",x"8000",x"3a42",x"3b80",x"b669",x"4042",x"36da",x"a65f",x"bbff",x"0000",x"3a42",x"3b89",x"b669",x"4042",x"3710",x"abae",x"bbfc",x"0000",x"3a4c",x"3b89"),
(x"b568",x"4058",x"36da",x"b810",x"3ae4",x"8000",x"3a8b",x"3b7d",x"b558",x"4059",x"36da",x"b02d",x"3bee",x"0000",x"3a8b",x"3b80",x"b558",x"4059",x"3710",x"b3cc",x"3bc2",x"8000",x"3a96",x"3b80"),
(x"b62a",x"4041",x"36da",x"2fb9",x"bbf1",x"0000",x"3a42",x"3b7c",x"b63d",x"4041",x"36da",x"affc",x"bbf0",x"8000",x"3a42",x"3b80",x"b63d",x"4041",x"3710",x"ab45",x"bbfc",x"0000",x"3a4c",x"3b80"),
(x"b558",x"4059",x"36da",x"b02d",x"3bee",x"0000",x"3a8b",x"3b80",x"b544",x"4059",x"36da",x"b46b",x"3bb0",x"0000",x"3a8b",x"3b84",x"b544",x"4059",x"3710",x"b138",x"3be4",x"0000",x"3a96",x"3b84"),
(x"b575",x"4038",x"36da",x"bb97",x"b50d",x"0000",x"3a42",x"3b4c",x"b575",x"403a",x"36da",x"ba67",x"38cb",x"868d",x"3a42",x"3b4e",x"b575",x"403a",x"3710",x"bb59",x"3650",x"8000",x"3a4c",x"3b4e"),
(x"b544",x"4059",x"36da",x"b46b",x"3bb0",x"0000",x"3a8b",x"3b84",x"b52b",x"405a",x"36da",x"b237",x"3bd8",x"0000",x"3a8b",x"3b89",x"b52b",x"405a",x"3710",x"b472",x"3baf",x"0000",x"3a96",x"3b89"),
(x"b5ce",x"4043",x"36da",x"2f26",x"bbf3",x"0000",x"3a42",x"3b6a",x"b62a",x"4041",x"36da",x"2fb9",x"bbf1",x"0000",x"3a42",x"3b7c",x"b62a",x"4041",x"3710",x"303a",x"bbed",x"0000",x"3a4c",x"3b7c"),
(x"b52b",x"405a",x"36da",x"b237",x"3bd8",x"0000",x"3a8b",x"3b89",x"b50d",x"405b",x"36da",x"324a",x"3bd8",x"8000",x"3a8b",x"3b8f",x"b50d",x"405b",x"3710",x"253f",x"3bff",x"0000",x"3a96",x"3b8f"),
(x"b5bd",x"4043",x"36da",x"b559",x"bb8a",x"0000",x"3a42",x"3b66",x"b5ce",x"4043",x"36da",x"2f26",x"bbf3",x"0000",x"3a42",x"3b6a",x"b5ce",x"4043",x"3710",x"2ae9",x"bbfc",x"0000",x"3a4c",x"3b6a"),
(x"b50d",x"405b",x"36da",x"324a",x"3bd8",x"8000",x"3a8b",x"3b8f",x"b4f9",x"405a",x"36da",x"3a57",x"38e0",x"8000",x"3a8b",x"3b93",x"b4f9",x"405a",x"3710",x"38a5",x"3a82",x"068d",x"3a96",x"3b93"),
(x"b5a1",x"4041",x"36da",x"b72c",x"bb26",x"8000",x"3a42",x"3b60",x"b5bd",x"4043",x"36da",x"b559",x"bb8a",x"0000",x"3a42",x"3b66",x"b5bd",x"4043",x"3710",x"b6e1",x"bb38",x"0000",x"3a4c",x"3b66"),
(x"b4f9",x"405a",x"36da",x"3a57",x"38e0",x"8000",x"3a8b",x"3b93",x"b4f5",x"4058",x"36da",x"3bc4",x"33a2",x"0000",x"3a8b",x"3b96",x"b4f5",x"4058",x"3710",x"3bbb",x"341b",x"8000",x"3a96",x"3b96"),
(x"b581",x"403f",x"36da",x"b794",x"bb0b",x"0000",x"3a42",x"3b59",x"b5a1",x"4041",x"36da",x"b72c",x"bb26",x"8000",x"3a42",x"3b60",x"b5a1",x"4041",x"3710",x"b67b",x"bb50",x"8000",x"3a4c",x"3b60"),
(x"b4f5",x"4058",x"36da",x"3bc4",x"33a2",x"0000",x"3a8b",x"3b96",x"b4f2",x"4056",x"36da",x"3a46",x"38f6",x"0000",x"3a8b",x"3b98",x"b4f2",x"4056",x"3710",x"3aea",x"3805",x"8000",x"3a96",x"3b98"),
(x"b931",x"404d",x"36da",x"bbff",x"a4d0",x"0000",x"39d6",x"33f3",x"b931",x"4059",x"36da",x"bbff",x"a4d0",x"0000",x"39e9",x"33f9",x"b931",x"4059",x"3710",x"bbfe",x"a4d0",x"28c6",x"39ea",x"33c9"),
(x"b8ff",x"4059",x"36da",x"26a7",x"3bff",x"8000",x"3a2d",x"3b9f",x"b8a3",x"4058",x"36da",x"2a59",x"3bfd",x"0000",x"3a2d",x"3b7b",x"b8a3",x"4058",x"3710",x"286a",x"3bfe",x"8000",x"3a23",x"3b7b"),
(x"b568",x"403c",x"36da",x"b9f3",x"b958",x"0000",x"3a42",x"3b53",x"b581",x"403f",x"36da",x"b794",x"bb0b",x"0000",x"3a42",x"3b59",x"b581",x"403f",x"3710",x"b89f",x"ba87",x"0000",x"3a4c",x"3b59"),
(x"b4f2",x"4056",x"36da",x"3a46",x"38f6",x"0000",x"3a8b",x"3b98",x"b4da",x"4053",x"36da",x"3afc",x"37cc",x"0000",x"3a8b",x"3b9f",x"b4da",x"4053",x"3710",x"3a4b",x"38ef",x"0000",x"3a96",x"3b9f"),
(x"b8a3",x"4058",x"36da",x"2a59",x"3bfd",x"0000",x"3a2d",x"3b7b",x"b89e",x"4058",x"36da",x"380f",x"3ae4",x"068d",x"3a2d",x"3b79",x"b89e",x"4058",x"3710",x"36f0",x"3b35",x"0000",x"3a23",x"3b79"),
(x"b558",x"4036",x"36da",x"b3cc",x"bbc2",x"8000",x"3a42",x"3b44",x"b568",x"4037",x"36da",x"b919",x"ba29",x"0000",x"3a42",x"3b48",x"b568",x"4037",x"3710",x"b810",x"bae4",x"0000",x"3a4c",x"3b48"),
(x"b4da",x"4053",x"36da",x"3afc",x"37cc",x"0000",x"3a8b",x"3b9f",x"b4d8",x"4051",x"36da",x"3af9",x"b7d8",x"8000",x"3a8b",x"3ba1",x"b4d8",x"4051",x"3710",x"3be5",x"b11d",x"868d",x"3a96",x"3ba1"),
(x"b89e",x"4058",x"36da",x"380f",x"3ae4",x"068d",x"3a2d",x"3b79",x"b88f",x"4055",x"36da",x"377a",x"3b12",x"0000",x"3a2d",x"3b72",x"b88f",x"4055",x"3710",x"380a",x"3ae7",x"0000",x"3a23",x"3b72"),
(x"b544",x"4036",x"36da",x"b138",x"bbe4",x"0000",x"3a42",x"3b40",x"b558",x"4036",x"36da",x"b3cc",x"bbc2",x"8000",x"3a42",x"3b44",x"b558",x"4036",x"3710",x"b02d",x"bbee",x"0000",x"3a4c",x"3b44"),
(x"b4d8",x"4051",x"36da",x"3af9",x"b7d8",x"8000",x"3a8b",x"3ba1",x"b4e1",x"4050",x"36da",x"33d2",x"bbc1",x"8000",x"3a8b",x"3ba3",x"b4e1",x"4050",x"3710",x"3599",x"bb7e",x"0000",x"3a96",x"3ba3"),
(x"b88f",x"4055",x"36da",x"377a",x"3b12",x"0000",x"3a2d",x"3b72",x"b87d",x"4053",x"36da",x"3244",x"3bd8",x"0000",x"3a2d",x"3b6a",x"b87d",x"4053",x"3710",x"3541",x"3b8e",x"0000",x"3a23",x"3b6a"),
(x"b52b",x"4035",x"36da",x"b472",x"bbaf",x"0000",x"3a42",x"3b3b",x"b544",x"4036",x"36da",x"b138",x"bbe4",x"0000",x"3a42",x"3b40",x"b544",x"4036",x"3710",x"b46b",x"bbb0",x"0000",x"3a4c",x"3b40"),
(x"b4e1",x"4050",x"36da",x"33d2",x"bbc1",x"8000",x"3a8b",x"3ba3",x"b51a",x"404f",x"36da",x"347c",x"bbad",x"0000",x"3a8b",x"3bae",x"b51a",x"404f",x"3710",x"332b",x"bbcb",x"0000",x"3a96",x"3bae"),
(x"b87d",x"4053",x"36da",x"3244",x"3bd8",x"0000",x"3a2d",x"3b6a",x"b86e",x"4053",x"36da",x"b407",x"3bbe",x"8000",x"3a2d",x"3b64",x"b86e",x"4053",x"3710",x"ad02",x"3bf9",x"0000",x"3a23",x"3b64"),
(x"b50d",x"4034",x"36da",x"253f",x"bbff",x"8000",x"3a42",x"3b35",x"b52b",x"4035",x"36da",x"b472",x"bbaf",x"0000",x"3a42",x"3b3b",x"b52b",x"4035",x"3710",x"b237",x"bbd8",x"0000",x"3a4c",x"3b3b"),
(x"b51a",x"404f",x"36da",x"347c",x"bbad",x"0000",x"3a8b",x"3bae",x"b528",x"404e",x"36da",x"38ed",x"ba4d",x"8000",x"3a8b",x"3bb1",x"b528",x"404e",x"3710",x"37ff",x"baed",x"0000",x"3a96",x"3bb1"),
(x"b86e",x"4053",x"36da",x"b407",x"3bbe",x"8000",x"3a2d",x"3b64",x"b867",x"4054",x"36da",x"baa2",x"3877",x"0000",x"3a2d",x"3b61",x"b867",x"4054",x"3710",x"b975",x"39d8",x"0000",x"3a23",x"3b61"),
(x"b4f9",x"4035",x"36da",x"38a5",x"ba82",x"8000",x"3a42",x"3b31",x"b50d",x"4034",x"36da",x"253f",x"bbff",x"8000",x"3a42",x"3b35",x"b50d",x"4034",x"3710",x"324a",x"bbd8",x"8000",x"3a4c",x"3b35"),
(x"b528",x"404e",x"36da",x"38ed",x"ba4d",x"8000",x"3a8b",x"3bb1",x"b52c",x"404e",x"36da",x"3b0d",x"378c",x"0000",x"3a8b",x"3bb2",x"b52c",x"404e",x"3710",x"3bfc",x"ab69",x"0000",x"3a96",x"3bb2"),
(x"b867",x"4054",x"36da",x"baa2",x"3877",x"0000",x"3a2d",x"3b61",x"b865",x"4055",x"36da",x"baaf",x"3865",x"8000",x"3a2d",x"3b5e",x"b865",x"4055",x"3710",x"bb0e",x"378a",x"0000",x"3a23",x"3b5e"),
(x"b4f5",x"4037",x"36da",x"3bbb",x"b41b",x"8000",x"3a42",x"3b2e",x"b4f9",x"4035",x"36da",x"38a5",x"ba82",x"8000",x"3a42",x"3b31",x"b4f9",x"4035",x"3710",x"3a57",x"b8e0",x"0000",x"3a4c",x"3b31"),
(x"b52c",x"404e",x"36da",x"3b0d",x"378c",x"0000",x"3b11",x"39ae",x"b526",x"404d",x"36da",x"33bb",x"3bc3",x"0000",x"3b11",x"39af",x"b526",x"404d",x"3710",x"35f8",x"3b6b",x"0000",x"3b1c",x"39af"),
(x"b865",x"4055",x"36da",x"baaf",x"3865",x"8000",x"3a2d",x"3b5e",x"b85e",x"4058",x"36da",x"b5f3",x"3b6d",x"8000",x"3a2d",x"3b5a",x"b85e",x"4058",x"3710",x"b878",x"3aa2",x"0000",x"3a23",x"3b5a"),
(x"b4f2",x"4038",x"36da",x"3aea",x"b805",x"8000",x"3a42",x"3b2b",x"b4f5",x"4037",x"36da",x"3bbb",x"b41b",x"8000",x"3a42",x"3b2e",x"b4f5",x"4037",x"3710",x"3bc4",x"b3a1",x"8000",x"3a4c",x"3b2e"),
(x"b526",x"404d",x"36da",x"33bb",x"3bc3",x"0000",x"3b11",x"39af",x"b50c",x"404c",x"36da",x"236c",x"3bff",x"0000",x"3b11",x"39b4",x"b50c",x"404c",x"3710",x"292b",x"3bfe",x"8000",x"3b1c",x"39b4"),
(x"b116",x"404a",x"36da",x"3bdf",x"31b0",x"868d",x"3a50",x"3b6f",x"b116",x"4045",x"36da",x"3b51",x"b675",x"8000",x"3a50",x"3b75",x"b116",x"4045",x"3710",x"3bdf",x"b1b0",x"0000",x"3a5a",x"3b75"),
(x"b85e",x"4058",x"36da",x"b5f3",x"3b6d",x"8000",x"3a2d",x"3b5a",x"b84a",x"4059",x"36da",x"30e0",x"3be8",x"8000",x"3a2d",x"3b51",x"b84a",x"4059",x"3710",x"ac15",x"3bfb",x"868d",x"3a23",x"3b51"),
(x"b4da",x"403c",x"36da",x"3a4b",x"b8ef",x"068d",x"3a42",x"3b24",x"b4f2",x"4038",x"36da",x"3aea",x"b805",x"8000",x"3a42",x"3b2b",x"b4f2",x"4038",x"3710",x"3a46",x"b8f6",x"0000",x"3a4c",x"3b2b"),
(x"b451",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3b11",x"39d8",x"b441",x"404d",x"36da",x"b7a3",x"3b07",x"0000",x"3b11",x"39db",x"b441",x"404d",x"3710",x"b6f3",x"3b34",x"0000",x"3b1c",x"39db"),
(x"b89e",x"4037",x"36da",x"36f0",x"bb35",x"0000",x"39fd",x"3b76",x"b8a3",x"4037",x"36da",x"2850",x"bbfe",x"8000",x"39fd",x"3b78",x"b8a3",x"4037",x"3710",x"2a1e",x"bbfd",x"0000",x"3a07",x"3b78"),
(x"b84a",x"4059",x"36da",x"30e0",x"3be8",x"8000",x"3a2d",x"3b51",x"b83a",x"4057",x"36da",x"3953",x"39f7",x"8000",x"3a2d",x"3b4b",x"b83a",x"4057",x"3710",x"3890",x"3a92",x"0000",x"3a23",x"3b4b"),
(x"b4d8",x"403d",x"36da",x"3be5",x"311d",x"0000",x"3a42",x"3b22",x"b4da",x"403c",x"36da",x"3a4b",x"b8ef",x"068d",x"3a42",x"3b24",x"b4da",x"403c",x"3710",x"3afc",x"b7cc",x"8000",x"3a4c",x"3b24"),
(x"b50c",x"404c",x"36da",x"236c",x"3bff",x"0000",x"3b11",x"39b4",x"b451",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3b11",x"39d8",x"b451",x"404c",x"3710",x"a0dd",x"3c00",x"0000",x"3b1c",x"39d8"),
(x"b88f",x"403a",x"36da",x"380a",x"bae7",x"0000",x"39fd",x"3b6f",x"b89e",x"4037",x"36da",x"36f0",x"bb35",x"0000",x"39fd",x"3b76",x"b89e",x"4037",x"3710",x"380f",x"bae4",x"068d",x"3a07",x"3b76"),
(x"b568",x"4053",x"36da",x"bb03",x"37b2",x"868d",x"3a8b",x"3b72",x"b569",x"4054",x"36da",x"ba4b",x"b8f0",x"0000",x"3a8b",x"3b74",x"b569",x"4054",x"3710",x"bb2d",x"b70f",x"0000",x"3a96",x"3b74"),
(x"b4e1",x"403e",x"36da",x"3599",x"3b7e",x"0000",x"3a42",x"3b1f",x"b4d8",x"403d",x"36da",x"3be5",x"311d",x"0000",x"3a42",x"3b22",x"b4d8",x"403d",x"3710",x"3af9",x"37d7",x"868d",x"3a4c",x"3b22"),
(x"b441",x"404d",x"36da",x"b7a3",x"3b07",x"0000",x"3b11",x"39db",x"b40d",x"4051",x"36da",x"b8bf",x"3a70",x"068d",x"3b11",x"39e6",x"b40d",x"4051",x"3710",x"b83a",x"3aca",x"0000",x"3b1c",x"39e6"),
(x"b87d",x"403c",x"36da",x"3541",x"bb8e",x"0000",x"39fd",x"3b67",x"b88f",x"403a",x"36da",x"380a",x"bae7",x"0000",x"39fd",x"3b6f",x"b88f",x"403a",x"3710",x"377a",x"bb12",x"8000",x"3a07",x"3b6f"),
(x"b83a",x"4057",x"36da",x"3953",x"39f7",x"8000",x"3a2d",x"3b4b",x"b820",x"4051",x"36da",x"385c",x"3ab4",x"0000",x"3a2d",x"3b3c",x"b820",x"4051",x"3710",x"391f",x"3a25",x"0000",x"3a23",x"3b3c"),
(x"b51a",x"4040",x"36da",x"332b",x"3bcb",x"0000",x"3a42",x"3b14",x"b4e1",x"403e",x"36da",x"3599",x"3b7e",x"0000",x"3a42",x"3b1f",x"b4e1",x"403e",x"3710",x"33d2",x"3bc1",x"868d",x"3a4c",x"3b1f"),
(x"b40d",x"4051",x"36da",x"b8bf",x"3a70",x"068d",x"3b11",x"39e6",x"b407",x"4052",x"36da",x"bbf7",x"2ddc",x"0000",x"3b11",x"39e8",x"b407",x"4052",x"3710",x"bb61",x"362a",x"0000",x"3b1c",x"39e8"),
(x"b86e",x"403c",x"36da",x"ad01",x"bbf9",x"0000",x"39fd",x"3b61",x"b87d",x"403c",x"36da",x"3541",x"bb8e",x"0000",x"39fd",x"3b67",x"b87d",x"403c",x"3710",x"3244",x"bbd8",x"0000",x"3a07",x"3b67"),
(x"b569",x"4054",x"36da",x"ba4b",x"b8f0",x"0000",x"3a8b",x"3b74",x"b575",x"4055",x"36da",x"bb59",x"b650",x"8000",x"3a8b",x"3b77",x"b575",x"4055",x"3710",x"ba67",x"b8cb",x"0000",x"3a96",x"3b77"),
(x"b528",x"4041",x"36da",x"37fe",x"3aed",x"0000",x"3a42",x"3b11",x"b51a",x"4040",x"36da",x"332b",x"3bcb",x"0000",x"3a42",x"3b14",x"b51a",x"4040",x"3710",x"347c",x"3bad",x"8000",x"3a4c",x"3b14"),
(x"b407",x"4052",x"36da",x"bbf7",x"2ddc",x"0000",x"3b11",x"39e8",x"b409",x"4053",x"36da",x"bab5",x"b85b",x"0000",x"3b11",x"39e9",x"b409",x"4053",x"3710",x"bb1a",x"b75c",x"8000",x"3b1c",x"39e9"),
(x"b867",x"403b",x"36da",x"b975",x"b9d8",x"0000",x"39fd",x"3b5e",x"b86e",x"403c",x"36da",x"ad01",x"bbf9",x"0000",x"39fd",x"3b61",x"b86e",x"403c",x"3710",x"b406",x"bbbe",x"0000",x"3a07",x"3b61"),
(x"b820",x"4051",x"36da",x"385c",x"3ab4",x"0000",x"3a2d",x"3b3c",x"b801",x"404d",x"36da",x"3346",x"3bca",x"0000",x"3a2d",x"3b2e",x"b801",x"404d",x"3710",x"3561",x"3b88",x"0000",x"3a23",x"3b2e"),
(x"b52c",x"4041",x"36da",x"3bfc",x"2b6f",x"0000",x"3a42",x"3b10",x"b528",x"4041",x"36da",x"37fe",x"3aed",x"0000",x"3a42",x"3b11",x"b528",x"4041",x"3710",x"38ed",x"3a4d",x"8000",x"3a4c",x"3b11"),
(x"b409",x"4053",x"36da",x"bab5",x"b85b",x"0000",x"3b11",x"39e9",x"b413",x"4054",x"36da",x"bba9",x"b499",x"0000",x"3b11",x"39ed",x"b413",x"4054",x"3710",x"bb08",x"b7a1",x"868d",x"3b1c",x"39ed"),
(x"b865",x"4039",x"36da",x"bb0e",x"b78a",x"0000",x"39fd",x"3b5b",x"b867",x"403b",x"36da",x"b975",x"b9d8",x"0000",x"39fd",x"3b5e",x"b867",x"403b",x"3710",x"baa2",x"b877",x"0000",x"3a07",x"3b5e"),
(x"b801",x"404d",x"36da",x"3346",x"3bca",x"0000",x"3a2d",x"3b2e",x"b7c0",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3a2d",x"3b21",x"b7c0",x"404c",x"3710",x"29e3",x"3bfd",x"0000",x"3a23",x"3b21"),
(x"b526",x"4042",x"36da",x"35f9",x"bb6b",x"0000",x"3af0",x"3a0f",x"b52c",x"4041",x"36da",x"3bfc",x"2b6f",x"0000",x"3af0",x"3a11",x"b52c",x"4041",x"3710",x"3b0d",x"b78c",x"0000",x"3afb",x"3a11"),
(x"b413",x"4054",x"36da",x"bba9",x"b499",x"0000",x"3b11",x"39ed",x"b413",x"4055",x"36da",x"ba12",x"3935",x"8000",x"3b11",x"39ee",x"b413",x"4055",x"3710",x"bb8c",x"354a",x"868d",x"3b1c",x"39ee"),
(x"b85e",x"4037",x"36da",x"b878",x"baa2",x"0000",x"39fd",x"3b57",x"b865",x"4039",x"36da",x"bb0e",x"b78a",x"0000",x"39fd",x"3b5b",x"b865",x"4039",x"3710",x"baaf",x"b865",x"8000",x"3a07",x"3b5b"),
(x"b7c0",x"404c",x"36da",x"a984",x"3bfe",x"8000",x"3a2d",x"3b21",x"b794",x"404d",x"36da",x"b51c",x"3b94",x"0000",x"3a2d",x"3b18",x"b794",x"404d",x"3710",x"b357",x"3bc9",x"0000",x"3a23",x"3b18"),
(x"b50c",x"4042",x"36da",x"292b",x"bbfe",x"8000",x"3af0",x"3a0a",x"b526",x"4042",x"36da",x"35f9",x"bb6b",x"0000",x"3af0",x"3a0f",x"b526",x"4042",x"3710",x"33bc",x"bbc3",x"0000",x"3afb",x"3a0f"),
(x"b413",x"4055",x"36da",x"ba12",x"3935",x"8000",x"3b11",x"39ee",x"b40b",x"4056",x"36da",x"aabe",x"3bfd",x"868d",x"3b11",x"39f0",x"b40b",x"4056",x"3710",x"b3aa",x"3bc4",x"8000",x"3b1c",x"39f0"),
(x"b84a",x"4036",x"36da",x"ac15",x"bbfb",x"068d",x"39fd",x"3b4e",x"b85e",x"4037",x"36da",x"b878",x"baa2",x"0000",x"39fd",x"3b57",x"b85e",x"4037",x"3710",x"b5f3",x"bb6d",x"8000",x"3a07",x"3b57"),
(x"b794",x"404d",x"36da",x"b51c",x"3b94",x"0000",x"3a2d",x"3b18",x"b77a",x"404e",x"36da",x"b97c",x"39d2",x"0000",x"3a2d",x"3b13",x"b77a",x"404e",x"3710",x"b83f",x"3ac7",x"0000",x"3a23",x"3b13"),
(x"b441",x"4042",x"36da",x"b6f3",x"bb34",x"0000",x"3af0",x"39e4",x"b451",x"4042",x"36da",x"a0ea",x"bc00",x"0000",x"3af0",x"39e7",x"b451",x"4042",x"3710",x"a987",x"bbfe",x"8000",x"3afb",x"39e7"),
(x"b40b",x"4056",x"36da",x"aabe",x"3bfd",x"868d",x"3b11",x"39f0",x"b3f4",x"4056",x"36da",x"3408",x"3bbd",x"0000",x"3b11",x"39f3",x"b3f4",x"4056",x"3710",x"3148",x"3be3",x"8000",x"3b1c",x"39f3"),
(x"b83a",x"4037",x"36da",x"3890",x"ba92",x"0000",x"39fd",x"3b48",x"b84a",x"4036",x"36da",x"ac15",x"bbfb",x"068d",x"39fd",x"3b4e",x"b84a",x"4036",x"3710",x"30e0",x"bbe8",x"8000",x"3a07",x"3b4e"),
(x"b77a",x"404e",x"36da",x"b97c",x"39d2",x"0000",x"3a2d",x"3b13",x"b776",x"4050",x"36da",x"bbce",x"b2fb",x"0000",x"3a2d",x"3b10",x"b776",x"4050",x"3710",x"bbee",x"3037",x"0000",x"3a23",x"3b10"),
(x"b451",x"4042",x"36da",x"a0ea",x"bc00",x"0000",x"3af0",x"39e7",x"b50c",x"4042",x"36da",x"292b",x"bbfe",x"8000",x"3af0",x"3a0a",x"b50c",x"4042",x"3710",x"236c",x"bbff",x"0000",x"3afb",x"3a0a"),
(x"b3f4",x"4056",x"36da",x"3408",x"3bbd",x"0000",x"3b11",x"39f3",x"b3d2",x"4055",x"36da",x"abf9",x"3bfc",x"0000",x"3b11",x"39f7",x"b3d2",x"4055",x"3710",x"2ffb",x"3bf0",x"0000",x"3b1c",x"39f7"),
(x"b569",x"403b",x"36da",x"bb2d",x"370f",x"0000",x"3a42",x"3b51",x"b568",x"403c",x"36da",x"b9f3",x"b958",x"0000",x"3a42",x"3b53",x"b568",x"403c",x"3710",x"bb03",x"b7b1",x"868d",x"3a4c",x"3b53"),
(x"b776",x"4050",x"36da",x"bbce",x"b2fb",x"0000",x"3a2d",x"3b10",x"b77b",x"4051",x"36da",x"b853",x"baba",x"0000",x"3a2d",x"3b0f",x"b77b",x"4051",x"3710",x"b937",x"ba10",x"0000",x"3a23",x"3b0f"),
(x"b40d",x"403e",x"36da",x"b83a",x"baca",x"0000",x"3af0",x"39d8",x"b441",x"4042",x"36da",x"b6f3",x"bb34",x"0000",x"3af0",x"39e4",x"b441",x"4042",x"3710",x"b7a4",x"bb07",x"0000",x"3afb",x"39e4"),
(x"b3d2",x"4055",x"36da",x"abf9",x"3bfc",x"0000",x"3b11",x"39f7",x"b3a5",x"4056",x"36da",x"32b6",x"3bd2",x"068d",x"3b11",x"39fb",x"b3a5",x"4056",x"3710",x"24fd",x"3bff",x"0000",x"3b1c",x"39fb"),
(x"b820",x"403e",x"36da",x"391f",x"ba25",x"0000",x"39fd",x"3b39",x"b83a",x"4037",x"36da",x"3890",x"ba92",x"0000",x"39fd",x"3b48",x"b83a",x"4037",x"3710",x"3953",x"b9f7",x"068d",x"3a07",x"3b48"),
(x"b77b",x"4051",x"36da",x"b853",x"baba",x"0000",x"3a88",x"3ac5",x"b790",x"4052",x"36da",x"b461",x"bbb1",x"0000",x"3a88",x"3ac9",x"b790",x"4052",x"3710",x"b606",x"bb69",x"0000",x"3a93",x"3ac9"),
(x"b407",x"403d",x"36da",x"bb61",x"b629",x"0000",x"3af0",x"39d6",x"b40d",x"403e",x"36da",x"b83a",x"baca",x"0000",x"3af0",x"39d8",x"b40d",x"403e",x"3710",x"b8bf",x"ba70",x"8000",x"3afb",x"39d8"),
(x"b3a5",x"4056",x"36da",x"32b6",x"3bd2",x"068d",x"3b11",x"39fb",x"b368",x"4054",x"36da",x"3912",x"3a2f",x"8000",x"3b11",x"3a01",x"b368",x"4054",x"3710",x"37ea",x"3af3",x"8000",x"3b1c",x"3a01"),
(x"b575",x"403a",x"36da",x"ba67",x"38cb",x"868d",x"3a42",x"3b4e",x"b569",x"403b",x"36da",x"bb2d",x"370f",x"0000",x"3a42",x"3b51",x"b569",x"403b",x"3710",x"ba4b",x"38f0",x"0000",x"3a4c",x"3b51"),
(x"b790",x"4052",x"36da",x"b461",x"bbb1",x"0000",x"3a88",x"3ac9",x"b7a8",x"4053",x"36da",x"b4b8",x"bba4",x"8000",x"3a88",x"3ace",x"b7a8",x"4053",x"3710",x"b360",x"bbc8",x"0000",x"3a93",x"3ace"),
(x"b409",x"403c",x"36da",x"bb1a",x"375d",x"0000",x"3af0",x"39d5",x"b407",x"403d",x"36da",x"bb61",x"b629",x"0000",x"3af0",x"39d6",x"b407",x"403d",x"3710",x"bbf7",x"addb",x"0000",x"3afb",x"39d6"),
(x"b368",x"4054",x"36da",x"3912",x"3a2f",x"8000",x"3b11",x"3a01",x"b340",x"4051",x"36da",x"3b6b",x"35fb",x"8000",x"3b11",x"3a07",x"b340",x"4051",x"3710",x"3aba",x"3853",x"0000",x"3b1c",x"3a07"),
(x"b801",x"4042",x"36da",x"3561",x"bb88",x"0000",x"39fd",x"3b2b",x"b820",x"403e",x"36da",x"391f",x"ba25",x"0000",x"39fd",x"3b39",x"b820",x"403e",x"3710",x"385c",x"bab4",x"8000",x"3a07",x"3b39"),
(x"b7a8",x"4053",x"36da",x"b4b8",x"bba4",x"8000",x"3a88",x"3ace",x"b7bd",x"4054",x"36da",x"b821",x"bada",x"8000",x"3a88",x"3ad2",x"b7bd",x"4054",x"3710",x"b6d2",x"bb3c",x"0000",x"3a93",x"3ad2"),
(x"b413",x"403a",x"36da",x"bb07",x"37a1",x"8000",x"3af0",x"39d2",x"b409",x"403c",x"36da",x"bb1a",x"375d",x"0000",x"3af0",x"39d5",x"b409",x"403c",x"3710",x"bab5",x"385b",x"0000",x"3afb",x"39d5"),
(x"b340",x"4051",x"36da",x"3b6b",x"35fb",x"8000",x"3b11",x"3a07",x"b33a",x"404f",x"36da",x"3b88",x"b564",x"068d",x"3b11",x"3a0b",x"b33a",x"404f",x"3710",x"3bf6",x"ae02",x"8000",x"3b1c",x"3a0b"),
(x"b7c0",x"4043",x"36da",x"29e3",x"bbfd",x"0000",x"39fd",x"3b1e",x"b801",x"4042",x"36da",x"3561",x"bb88",x"0000",x"39fd",x"3b2b",x"b801",x"4042",x"3710",x"3346",x"bbca",x"0000",x"3a07",x"3b2b"),
(x"b7bd",x"4054",x"36da",x"b821",x"bada",x"8000",x"3a88",x"3ad2",x"b7c7",x"4055",x"36da",x"bb43",x"b6b4",x"0000",x"3a88",x"3ad5",x"b7c7",x"4055",x"3710",x"ba01",x"b948",x"0000",x"3a93",x"3ad5"),
(x"b931",x"4036",x"36da",x"bbff",x"26b5",x"0000",x"39b3",x"33fa",x"b930",x"4041",x"36da",x"bbff",x"26b5",x"0000",x"39c6",x"33f0",x"b930",x"4041",x"3710",x"bbeb",x"2604",x"3075",x"39c5",x"33c0"),
(x"b413",x"4039",x"36da",x"bb8c",x"b54a",x"868d",x"3af0",x"39d0",x"b413",x"403a",x"36da",x"bb07",x"37a1",x"8000",x"3af0",x"39d2",x"b413",x"403a",x"3710",x"bba9",x"3499",x"8000",x"3afb",x"39d2"),
(x"b33a",x"404f",x"36da",x"3b88",x"b564",x"068d",x"3b11",x"3a0b",x"b351",x"404d",x"36da",x"3bb2",x"b458",x"0000",x"3b11",x"3a0f",x"b351",x"404d",x"3710",x"3b23",x"b738",x"0000",x"3b1c",x"3a0f"),
(x"b794",x"4042",x"36da",x"b357",x"bbc9",x"0000",x"39fd",x"3b15",x"b7c0",x"4043",x"36da",x"29e3",x"bbfd",x"0000",x"39fd",x"3b1e",x"b7c0",x"4043",x"3710",x"a984",x"bbfe",x"0000",x"3a07",x"3b1e"),
(x"b7c7",x"4055",x"36da",x"bb43",x"b6b4",x"0000",x"3a88",x"3ad5",x"b7c7",x"4055",x"36da",x"b744",x"3b20",x"0cea",x"3a88",x"3ad6",x"b7c7",x"4055",x"3710",x"b8b7",x"3a76",x"0000",x"3a93",x"3ad6"),
(x"b40b",x"4039",x"36da",x"b3aa",x"bbc4",x"0000",x"3af0",x"39ce",x"b413",x"4039",x"36da",x"bb8c",x"b54a",x"868d",x"3af0",x"39d0",x"b413",x"4039",x"3710",x"ba12",x"b935",x"068d",x"3afb",x"39d0"),
(x"b351",x"404d",x"36da",x"3bb2",x"b458",x"0000",x"3b11",x"3a0f",x"b34f",x"404c",x"36da",x"3448",x"3bb5",x"0000",x"3b11",x"3a11",x"b34f",x"404c",x"3710",x"3913",x"3a2e",x"8000",x"3b1c",x"3a11"),
(x"b77a",x"4040",x"36da",x"b83f",x"bac7",x"0000",x"39fd",x"3b10",x"b794",x"4042",x"36da",x"b357",x"bbc9",x"0000",x"39fd",x"3b15",x"b794",x"4042",x"3710",x"b51c",x"bb94",x"0000",x"3a07",x"3b15"),
(x"b7c7",x"4055",x"36da",x"b744",x"3b20",x"0cea",x"3a88",x"3ad6",x"b7a4",x"4057",x"36da",x"b64b",x"3b5a",x"8000",x"3a88",x"3add",x"b7a4",x"4057",x"3710",x"b654",x"3b58",x"0000",x"3a93",x"3add"),
(x"b3f4",x"4039",x"36da",x"3148",x"bbe3",x"0000",x"3af0",x"39cb",x"b40b",x"4039",x"36da",x"b3aa",x"bbc4",x"0000",x"3af0",x"39ce",x"b40b",x"4039",x"3710",x"aabe",x"bbfd",x"8000",x"3afb",x"39ce"),
(x"b34f",x"404c",x"36da",x"3448",x"3bb5",x"0000",x"3a50",x"3b34",x"b326",x"404b",x"36da",x"ad8e",x"3bf8",x"0000",x"3a50",x"3b38",x"b326",x"404b",x"3710",x"a5e9",x"3bff",x"0000",x"3a5a",x"3b38"),
(x"b776",x"403f",x"36da",x"bbee",x"b037",x"0000",x"3b18",x"38a2",x"b77a",x"4040",x"36da",x"b83f",x"bac7",x"0000",x"3b16",x"38a2",x"b77a",x"4040",x"3710",x"b97c",x"b9d2",x"8000",x"3b16",x"38ac"),
(x"b7a4",x"4057",x"36da",x"b64b",x"3b5a",x"8000",x"3a88",x"3add",x"b783",x"4059",x"36da",x"afa0",x"3bf1",x"0000",x"3a88",x"3ae4",x"b783",x"4059",x"3710",x"b33d",x"3bca",x"0000",x"3a93",x"3ae4"),
(x"b3d2",x"403a",x"36da",x"2ffb",x"bbf0",x"0000",x"3af0",x"39c8",x"b3f4",x"4039",x"36da",x"3148",x"bbe3",x"0000",x"3af0",x"39cb",x"b3f4",x"4039",x"3710",x"3408",x"bbbd",x"0000",x"3afb",x"39cb"),
(x"b326",x"404b",x"36da",x"ad8e",x"3bf8",x"0000",x"3a50",x"3b38",x"b2d6",x"404c",x"36da",x"b4dd",x"3b9f",x"0000",x"3a50",x"3b3f",x"b2d6",x"404c",x"3710",x"b287",x"3bd4",x"0000",x"3a5a",x"3b3f"),
(x"b77b",x"403e",x"36da",x"b937",x"3a10",x"8000",x"3b1a",x"38a2",x"b776",x"403f",x"36da",x"bbee",x"b037",x"0000",x"3b18",x"38a2",x"b776",x"403f",x"3710",x"bbce",x"32fb",x"0000",x"3b18",x"38ac"),
(x"b783",x"4059",x"36da",x"afa0",x"3bf1",x"0000",x"3a88",x"3ae4",x"b73e",x"4059",x"36da",x"2f57",x"3bf2",x"8000",x"3a88",x"3af1",x"b73e",x"4059",x"3710",x"27ae",x"3bfe",x"0000",x"3a93",x"3af1"),
(x"b3a5",x"4039",x"36da",x"2504",x"bbff",x"0000",x"3af0",x"39c3",x"b3d2",x"403a",x"36da",x"2ffb",x"bbf0",x"0000",x"3af0",x"39c8",x"b3d2",x"403a",x"3710",x"abf9",x"bbfc",x"8000",x"3afb",x"39c8"),
(x"b2d6",x"404c",x"36da",x"b4dd",x"3b9f",x"0000",x"3a50",x"3b3f",x"b2aa",x"404d",x"36da",x"b7e2",x"3af5",x"0000",x"3a50",x"3b44",x"b2aa",x"404d",x"3710",x"b78b",x"3b0e",x"0000",x"3a5a",x"3b44"),
(x"b790",x"403d",x"36da",x"b606",x"3b69",x"0000",x"3b1e",x"38a2",x"b77b",x"403e",x"36da",x"b937",x"3a10",x"8000",x"3b1a",x"38a2",x"b77b",x"403e",x"3710",x"b853",x"3aba",x"0000",x"3b1a",x"38ac"),
(x"b73e",x"4059",x"36da",x"2f57",x"3bf2",x"8000",x"3a88",x"3af1",x"b705",x"4058",x"36da",x"36ee",x"3b35",x"0000",x"3a88",x"3afc",x"b705",x"4058",x"3710",x"34b8",x"3ba4",x"0000",x"3a93",x"3afc"),
(x"b368",x"403a",x"36da",x"37ea",x"baf3",x"8000",x"3af0",x"39bd",x"b3a5",x"4039",x"36da",x"2504",x"bbff",x"0000",x"3af0",x"39c3",x"b3a5",x"4039",x"3710",x"32b6",x"bbd2",x"0000",x"3afb",x"39c3"),
(x"b2aa",x"404d",x"36da",x"b7e2",x"3af5",x"0000",x"3a50",x"3b44",x"b261",x"4050",x"36da",x"b5e0",x"3b70",x"8000",x"3a50",x"3b4c",x"b261",x"4050",x"3710",x"b72e",x"3b26",x"8000",x"3a5a",x"3b4c"),
(x"b7a8",x"403c",x"36da",x"b360",x"3bc8",x"8000",x"3a72",x"3b0f",x"b790",x"403d",x"36da",x"b606",x"3b69",x"0000",x"3a72",x"3b13",x"b790",x"403d",x"3710",x"b461",x"3bb1",x"0000",x"3a7c",x"3b13"),
(x"b705",x"4058",x"36da",x"36ee",x"3b35",x"0000",x"3a88",x"3afc",x"b6f1",x"4056",x"36da",x"3b73",x"35d3",x"8000",x"3a88",x"3b01",x"b6f1",x"4056",x"3710",x"3a69",x"38c9",x"068d",x"3a93",x"3b01"),
(x"b340",x"403d",x"36da",x"3aba",x"b853",x"8000",x"3af0",x"39b7",x"b368",x"403a",x"36da",x"37ea",x"baf3",x"8000",x"3af0",x"39bd",x"b368",x"403a",x"3710",x"3912",x"ba2f",x"0000",x"3afb",x"39bd"),
(x"b261",x"4050",x"36da",x"b5e0",x"3b70",x"8000",x"3a50",x"3b4c",x"b22d",x"4051",x"36da",x"2c28",x"3bfb",x"0000",x"3a50",x"3b51",x"b22d",x"4051",x"3710",x"ae8a",x"3bf5",x"8000",x"3a5a",x"3b51"),
(x"b7bd",x"403b",x"36da",x"b6d2",x"3b3c",x"0000",x"3a72",x"3b0b",x"b7a8",x"403c",x"36da",x"b360",x"3bc8",x"8000",x"3a72",x"3b0f",x"b7a8",x"403c",x"3710",x"b4b8",x"3ba4",x"8000",x"3a7c",x"3b0f"),
(x"b6f1",x"4056",x"36da",x"3b73",x"35d3",x"8000",x"3a88",x"3b01",x"b6ef",x"4053",x"36da",x"3b57",x"b659",x"8000",x"3a88",x"3b05",x"b6ef",x"4053",x"3710",x"3be9",x"b0b7",x"0000",x"3a93",x"3b05"),
(x"b33a",x"4040",x"36da",x"3bf6",x"2e02",x"8000",x"3af0",x"39b3",x"b340",x"403d",x"36da",x"3aba",x"b853",x"8000",x"3af0",x"39b7",x"b340",x"403d",x"3710",x"3b6b",x"b5fb",x"0000",x"3afb",x"39b7"),
(x"b22d",x"4051",x"36da",x"2c28",x"3bfb",x"0000",x"3a50",x"3b51",x"b1fd",x"4050",x"36da",x"375d",x"3b1a",x"8000",x"3a50",x"3b56",x"b1fd",x"4050",x"3710",x"35da",x"3b72",x"0000",x"3a5a",x"3b56"),
(x"b7c7",x"403a",x"36da",x"ba01",x"3948",x"8000",x"3a72",x"3b08",x"b7bd",x"403b",x"36da",x"b6d2",x"3b3c",x"0000",x"3a72",x"3b0b",x"b7bd",x"403b",x"3710",x"b821",x"3ada",x"8000",x"3a7c",x"3b0b"),
(x"b6ef",x"4053",x"36da",x"3b57",x"b659",x"8000",x"3a88",x"3b05",x"b6fb",x"4051",x"36da",x"37ed",x"baf2",x"068d",x"3a88",x"3b08",x"b6fb",x"4051",x"3710",x"38e1",x"ba57",x"0000",x"3a93",x"3b08"),
(x"b351",x"4042",x"36da",x"3b23",x"3738",x"0000",x"3af0",x"39af",x"b33a",x"4040",x"36da",x"3bf6",x"2e02",x"8000",x"3af0",x"39b3",x"b33a",x"4040",x"3710",x"3b88",x"3564",x"0000",x"3afb",x"39b3"),
(x"b1fd",x"4050",x"36da",x"375d",x"3b1a",x"8000",x"3a50",x"3b56",x"b1c1",x"404e",x"36da",x"3680",x"3b4f",x"8000",x"3a50",x"3b5d",x"b1c1",x"404e",x"3710",x"37bd",x"3b00",x"0000",x"3a5a",x"3b5d"),
(x"b7c7",x"4039",x"36da",x"b8b7",x"ba76",x"0000",x"3a72",x"3b07",x"b7c7",x"403a",x"36da",x"ba01",x"3948",x"8000",x"3a72",x"3b08",x"b7c7",x"403a",x"3710",x"bb43",x"36b4",x"0000",x"3a7c",x"3b08"),
(x"b6fb",x"4051",x"36da",x"37ed",x"baf2",x"068d",x"3a88",x"3b08",x"b721",x"404f",x"36da",x"37a6",x"bb06",x"0000",x"3a88",x"3b10",x"b721",x"404f",x"3710",x"3711",x"bb2d",x"0000",x"3a93",x"3b10"),
(x"b34f",x"4043",x"36da",x"3913",x"ba2f",x"8000",x"3af0",x"39ae",x"b351",x"4042",x"36da",x"3b23",x"3738",x"0000",x"3af0",x"39af",x"b351",x"4042",x"3710",x"3bb3",x"3458",x"0000",x"3afb",x"39af"),
(x"b1c1",x"404e",x"36da",x"3680",x"3b4f",x"8000",x"3a50",x"3b5d",x"b1a1",x"404d",x"36da",x"2ede",x"3bf4",x"0000",x"3a50",x"3b60",x"b1a1",x"404d",x"3710",x"314c",x"3be3",x"0000",x"3a5a",x"3b60"),
(x"b7a4",x"4038",x"36da",x"b654",x"bb58",x"8000",x"3a72",x"3b00",x"b7c7",x"4039",x"36da",x"b8b7",x"ba76",x"0000",x"3a72",x"3b07",x"b7c7",x"4039",x"3710",x"b744",x"bb20",x"868d",x"3a7c",x"3b07"),
(x"b721",x"404f",x"36da",x"37a6",x"bb06",x"0000",x"3a88",x"3b10",x"b72e",x"404e",x"36da",x"3b4f",x"b67e",x"8000",x"3a88",x"3b13",x"b72e",x"404e",x"3710",x"39a7",x"b9a8",x"0000",x"3a93",x"3b13"),
(x"b326",x"4043",x"36da",x"a5e9",x"bbff",x"0000",x"3a50",x"3bac",x"b34f",x"4043",x"36da",x"3913",x"ba2f",x"8000",x"3a50",x"3bb0",x"b34f",x"4043",x"3710",x"3448",x"bbb5",x"0000",x"3a5a",x"3bb0"),
(x"b1a1",x"404d",x"36da",x"2ede",x"3bf4",x"0000",x"3a50",x"3b60",x"b161",x"404d",x"36da",x"3407",x"3bbe",x"0000",x"3a50",x"3b66",x"b161",x"404d",x"3710",x"30d8",x"3be8",x"8000",x"3a5a",x"3b66"),
(x"b783",x"4036",x"36da",x"b33d",x"bbca",x"8000",x"3a72",x"3af9",x"b7a4",x"4038",x"36da",x"b654",x"bb58",x"8000",x"3a72",x"3b00",x"b7a4",x"4038",x"3710",x"b64a",x"bb5a",x"8000",x"3a7c",x"3b00"),
(x"b72e",x"404e",x"36da",x"3b4f",x"b67e",x"8000",x"3a8b",x"3b18",x"b72d",x"404d",x"36da",x"3778",x"3b13",x"0000",x"3a8b",x"3b19",x"b72d",x"404d",x"3710",x"3a45",x"38f8",x"0000",x"3a96",x"3b19"),
(x"b2d6",x"4043",x"36da",x"b287",x"bbd4",x"0000",x"3a50",x"3ba5",x"b326",x"4043",x"36da",x"a5e9",x"bbff",x"0000",x"3a50",x"3bac",x"b326",x"4043",x"3710",x"ad8e",x"bbf8",x"0000",x"3a5a",x"3bac"),
(x"b161",x"404d",x"36da",x"3407",x"3bbe",x"0000",x"3a50",x"3b66",x"b135",x"404c",x"36da",x"3934",x"3a13",x"8000",x"3a50",x"3b6a",x"b135",x"404c",x"3710",x"3822",x"3ad9",x"0000",x"3a5a",x"3b6a"),
(x"b73e",x"4035",x"36da",x"27ae",x"bbff",x"0000",x"3a72",x"3aec",x"b783",x"4036",x"36da",x"b33d",x"bbca",x"8000",x"3a72",x"3af9",x"b783",x"4036",x"3710",x"afa0",x"bbf1",x"0000",x"3a7c",x"3af9"),
(x"b72d",x"404d",x"36da",x"3778",x"3b13",x"0000",x"3a8b",x"3b19",x"b721",x"404c",x"36da",x"0cea",x"3c00",x"0000",x"3a8b",x"3b1c",x"b721",x"404c",x"3710",x"2560",x"3bff",x"0000",x"3a96",x"3b1c"),
(x"b2aa",x"4041",x"36da",x"b78b",x"bb0e",x"0000",x"3a50",x"3ba0",x"b2d6",x"4043",x"36da",x"b287",x"bbd4",x"0000",x"3a50",x"3ba5",x"b2d6",x"4043",x"3710",x"b4dc",x"bb9f",x"0000",x"3a5a",x"3ba5"),
(x"b135",x"404c",x"36da",x"3934",x"3a13",x"8000",x"3a50",x"3b6a",x"b116",x"404a",x"36da",x"3bdf",x"31b0",x"868d",x"3a50",x"3b6f",x"b116",x"404a",x"3710",x"3b51",x"3675",x"0000",x"3a5a",x"3b6f"),
(x"b705",x"4037",x"36da",x"34b8",x"bba4",x"8000",x"3a72",x"3ae1",x"b73e",x"4035",x"36da",x"27ae",x"bbff",x"0000",x"3a72",x"3aec",x"b73e",x"4035",x"3710",x"2f55",x"bbf2",x"0000",x"3a7c",x"3aec"),
(x"b575",x"4056",x"36da",x"bab5",x"385c",x"8000",x"3a8b",x"3b79",x"b568",x"4058",x"36da",x"b810",x"3ae4",x"8000",x"3a8b",x"3b7d",x"b568",x"4058",x"3710",x"b919",x"3a29",x"0000",x"3a96",x"3b7d"),
(x"b938",x"4042",x"36da",x"bbfe",x"a8f0",x"0000",x"3bea",x"39c8",x"b93a",x"404d",x"36da",x"bbfe",x"a8f0",x"0000",x"3bfb",x"39c9",x"b93a",x"404d",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3bfb",x"39bf"),
(x"b261",x"403f",x"36da",x"b72e",x"bb26",x"0000",x"3a50",x"3b98",x"b2aa",x"4041",x"36da",x"b78b",x"bb0e",x"0000",x"3a50",x"3ba0",x"b2aa",x"4041",x"3710",x"b7e2",x"baf5",x"0000",x"3a5a",x"3ba0"),
(x"b931",x"4059",x"36da",x"23ae",x"3bff",x"0000",x"3a2d",x"3bb3",x"b8ff",x"4059",x"36da",x"26a7",x"3bff",x"8000",x"3a2d",x"3b9f",x"b8ff",x"4059",x"3710",x"2581",x"3bff",x"15bc",x"3a23",x"3b9f"),
(x"b6f1",x"4039",x"36da",x"3a69",x"b8c9",x"868d",x"3a72",x"3adc",x"b705",x"4037",x"36da",x"34b8",x"bba4",x"8000",x"3a72",x"3ae1",x"b705",x"4037",x"3710",x"36ee",x"bb35",x"0000",x"3a7c",x"3ae1"),
(x"b721",x"404c",x"36da",x"0cea",x"3c00",x"0000",x"3a8b",x"3b1c",x"b669",x"404d",x"36da",x"abae",x"3bfc",x"8000",x"3a8b",x"3b3e",x"b669",x"404d",x"3710",x"a666",x"3bff",x"0000",x"3a96",x"3b3e"),
(x"b22d",x"403e",x"36da",x"ae8a",x"bbf5",x"8000",x"3a50",x"3b93",x"b261",x"403f",x"36da",x"b72e",x"bb26",x"0000",x"3a50",x"3b98",x"b261",x"403f",x"3710",x"b5e0",x"bb70",x"8000",x"3a5a",x"3b98"),
(x"b6ef",x"403c",x"36da",x"3be9",x"30b7",x"868d",x"3a72",x"3ad8",x"b6f1",x"4039",x"36da",x"3a69",x"b8c9",x"868d",x"3a72",x"3adc",x"b6f1",x"4039",x"3710",x"3b73",x"b5d3",x"0000",x"3a7c",x"3adc"),
(x"b669",x"404d",x"36da",x"abae",x"3bfc",x"8000",x"3a8b",x"3b3e",x"b63d",x"404e",x"36da",x"ab45",x"3bfc",x"0000",x"3a8b",x"3b47",x"b63d",x"404e",x"3710",x"affc",x"3bf0",x"0000",x"3a96",x"3b47"),
(x"b930",x"4041",x"36da",x"b67a",x"bb50",x"0000",x"3b21",x"387e",x"b938",x"4042",x"36da",x"b67a",x"bb50",x"0000",x"3b1f",x"387c",x"b938",x"4042",x"3710",x"b678",x"bb4d",x"2af3",x"3b19",x"3884"),
(x"a379",x"3ee5",x"36eb",x"bba3",x"b453",x"2fdf",x"3919",x"31f6",x"a271",x"3ee5",x"3718",x"bbb8",x"b22d",x"31b0",x"390e",x"31e7",x"a1bd",x"3ee0",x"3715",x"bbf4",x"2da3",x"2b3e",x"390d",x"31fc"),
(x"a379",x"3ee5",x"36eb",x"bba3",x"b453",x"2fdf",x"3919",x"31f6",x"a3d0",x"3eed",x"36eb",x"bb7a",x"3531",x"30a8",x"391c",x"31d5",x"a303",x"3eed",x"3715",x"bbda",x"2e4f",x"312f",x"3911",x"31c8"),
(x"a3d0",x"3eed",x"36eb",x"bb7a",x"3531",x"30a8",x"391c",x"31d5",x"a133",x"3ef6",x"36eb",x"b8c7",x"3a49",x"310c",x"391e",x"31a8",x"a0f3",x"3ef4",x"3714",x"ba0a",x"3915",x"3126",x"3914",x"31a4"),
(x"a133",x"3ef6",x"36eb",x"b8c7",x"3a49",x"310c",x"391e",x"31a8",x"9725",x"3efa",x"36eb",x"a3ae",x"3bec",x"3065",x"391f",x"3181",x"96c5",x"3ef8",x"3714",x"b236",x"3bc0",x"30e1",x"3915",x"317d"),
(x"9725",x"3efa",x"36eb",x"a3ae",x"3bec",x"3065",x"391f",x"3181",x"22b9",x"3ef8",x"36eb",x"36e0",x"3b1c",x"3118",x"3920",x"313f",x"21e6",x"3ef7",x"3714",x"335f",x"3baf",x"30fd",x"3916",x"3143"),
(x"22b9",x"3ef8",x"36eb",x"36e0",x"3b1c",x"3118",x"3920",x"313f",x"2505",x"3ef2",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3920",x"3117",x"24a4",x"3ef1",x"3715",x"3a37",x"38de",x"311d",x"3915",x"311d"),
(x"2505",x"3ef2",x"36eb",x"3b2d",x"36c9",x"2ff1",x"3920",x"3117",x"256c",x"3eea",x"36eb",x"3bf7",x"2138",x"2dcf",x"391f",x"30f5",x"252e",x"3eea",x"3715",x"3bf2",x"2495",x"2f43",x"3914",x"30fc"),
(x"250e",x"3ee3",x"36eb",x"3b9a",x"b4b0",x"2eb3",x"391d",x"30d7",x"24bc",x"3ee3",x"3715",x"3b87",x"b537",x"2d81",x"3913",x"30de",x"252e",x"3eea",x"3715",x"3bf2",x"2495",x"2f43",x"3914",x"30fc"),
(x"2470",x"3ede",x"36eb",x"3bfd",x"212b",x"29e6",x"391c",x"30c1",x"2464",x"3ede",x"3717",x"3bff",x"2481",x"2487",x"3911",x"30ca",x"24bc",x"3ee3",x"3715",x"3b87",x"b537",x"2d81",x"3913",x"30de"),
(x"250d",x"3ec4",x"36eb",x"3b9b",x"34d2",x"2ca7",x"3917",x"3054",x"25ec",x"3ec3",x"36eb",x"3b76",x"3593",x"2dee",x"3917",x"3044",x"25c0",x"3ec2",x"3714",x"3b74",x"35a6",x"2d5e",x"390d",x"304b"),
(x"2066",x"3edf",x"36eb",x"bbf7",x"9e73",x"2dbc",x"392c",x"2cc6",x"2019",x"3ee5",x"36eb",x"bb95",x"3495",x"306c",x"3927",x"2cc6",x"20c8",x"3ee4",x"3716",x"bbad",x"3434",x"2e8a",x"3928",x"2d1c"),
(x"2029",x"3ec5",x"36eb",x"ba79",x"3840",x"3401",x"3948",x"2cc1",x"2066",x"3edf",x"36eb",x"bbf7",x"9e73",x"2dbc",x"392c",x"2cc6",x"20e0",x"3edf",x"3718",x"bbf1",x"95bc",x"2fb4",x"392d",x"2d20"),
(x"a50e",x"3eb9",x"36eb",x"b409",x"bbbc",x"27db",x"3905",x"32b4",x"a4fc",x"3ec4",x"36eb",x"bbc6",x"328d",x"2f71",x"390a",x"3287",x"a4b5",x"3ec3",x"3715",x"bbb4",x"33e8",x"2ed7",x"3900",x"3276"),
(x"262b",x"3eb8",x"36eb",x"36d0",x"bb39",x"2aae",x"3914",x"3017",x"25f4",x"3eb9",x"3714",x"2f03",x"bbf3",x"23ef",x"390b",x"3022",x"25c0",x"3ec2",x"3714",x"3b74",x"35a6",x"2d5e",x"390d",x"304b"),
(x"9909",x"3ee3",x"3715",x"3b88",x"3531",x"2dc2",x"38ff",x"2d27",x"95ed",x"3ee4",x"36ee",x"3b70",x"358e",x"2fc0",x"38ff",x"2cd9",x"9651",x"3ee0",x"36eb",x"3bd3",x"b208",x"2da6",x"38fa",x"2cd5"),
(x"9caa",x"3ee8",x"36ee",x"3b20",x"3725",x"2d51",x"3904",x"2cda",x"95ed",x"3ee4",x"36ee",x"3b70",x"358e",x"2fc0",x"38ff",x"2cd9",x"9909",x"3ee3",x"3715",x"3b88",x"3531",x"2dc2",x"38ff",x"2d27"),
(x"9cff",x"3eec",x"36ee",x"3b1d",x"b747",x"2911",x"3909",x"2cda",x"9caa",x"3ee8",x"36ee",x"3b20",x"3725",x"2d51",x"3904",x"2cda",x"9db7",x"3ee9",x"3717",x"3bd6",x"323b",x"2a8a",x"3905",x"2d2c"),
(x"219c",x"3eec",x"36ee",x"ba30",x"b90f",x"2921",x"391e",x"2cd4",x"1f13",x"3ef0",x"36ee",x"b188",x"bbe0",x"a53f",x"3917",x"2cd5",x"1f52",x"3ef0",x"3715",x"b638",x"bb5e",x"243f",x"3918",x"2d23"),
(x"9fcf",x"3ec6",x"36eb",x"3be6",x"2cac",x"3077",x"38de",x"2ce5",x"a069",x"3ec3",x"3718",x"398b",x"396b",x"33db",x"38db",x"2d41",x"993e",x"3edf",x"3716",x"3bce",x"b2bb",x"2b41",x"38fa",x"2d2d"),
(x"9909",x"3ee3",x"3715",x"28d3",x"a80e",x"3bfd",x"3988",x"31f3",x"993e",x"3edf",x"3716",x"a82f",x"2808",x"3bfd",x"3988",x"31ea",x"a1bd",x"3ee0",x"3715",x"a1a1",x"23fc",x"3bff",x"3983",x"31eb"),
(x"9db7",x"3ee9",x"3717",x"250b",x"281b",x"3bfe",x"3987",x"31ff",x"9909",x"3ee3",x"3715",x"28d3",x"a80e",x"3bfd",x"3988",x"31f3",x"a271",x"3ee5",x"3718",x"28fa",x"a4f7",x"3bfe",x"3983",x"31f6"),
(x"9cfd",x"3eed",x"3716",x"252b",x"2c96",x"3bfa",x"3987",x"3208",x"9db7",x"3ee9",x"3717",x"250b",x"281b",x"3bfe",x"3987",x"31ff",x"a303",x"3eed",x"3715",x"9ec2",x"2bd5",x"3bfc",x"3982",x"3208"),
(x"94d9",x"3eef",x"3713",x"184d",x"9cd0",x"3c00",x"3989",x"320d",x"9cfd",x"3eed",x"3716",x"252b",x"2c96",x"3bfa",x"3987",x"3208",x"a0f3",x"3ef4",x"3714",x"263f",x"27c8",x"3bfe",x"3984",x"3218"),
(x"1f52",x"3ef0",x"3715",x"9cb5",x"191e",x"3c00",x"398e",x"320f",x"94d9",x"3eef",x"3713",x"184d",x"9cd0",x"3c00",x"3989",x"320d",x"96c5",x"3ef8",x"3714",x"a194",x"a0dd",x"3bff",x"3989",x"3221"),
(x"21f4",x"3eec",x"3714",x"9da1",x"252b",x"3bff",x"3991",x"3205",x"1f52",x"3ef0",x"3715",x"9cb5",x"191e",x"3c00",x"398e",x"320f",x"21e6",x"3ef7",x"3714",x"1df0",x"2487",x"3bff",x"3990",x"321e"),
(x"21f4",x"3eec",x"3714",x"9da1",x"252b",x"3bff",x"3991",x"3205",x"24a4",x"3ef1",x"3715",x"a793",x"184d",x"3bff",x"3994",x"3211",x"252e",x"3eea",x"3715",x"9818",x"26bb",x"3bff",x"3995",x"3201"),
(x"2211",x"3ee8",x"3716",x"2338",x"267a",x"3bff",x"3991",x"31fe",x"252e",x"3eea",x"3715",x"9818",x"26bb",x"3bff",x"3995",x"3201",x"24bc",x"3ee3",x"3715",x"2645",x"29e0",x"3bfd",x"3994",x"31f1"),
(x"20e0",x"3edf",x"3718",x"2793",x"243f",x"3bfe",x"398f",x"31ea",x"20c8",x"3ee4",x"3716",x"24bc",x"2b17",x"3bfc",x"398f",x"31f4",x"24bc",x"3ee3",x"3715",x"2645",x"29e0",x"3bfd",x"3994",x"31f1"),
(x"24de",x"3ec4",x"3717",x"2984",x"a0c2",x"3bfd",x"3995",x"31ae",x"2116",x"3ec2",x"3718",x"23ae",x"ac2f",x"3bfb",x"398f",x"31a9",x"20e0",x"3edf",x"3718",x"2793",x"243f",x"3bfe",x"398f",x"31ea"),
(x"21cf",x"3ee8",x"36ee",x"bb7c",x"357c",x"2d58",x"3921",x"2cd1",x"219c",x"3eec",x"36ee",x"ba30",x"b90f",x"2921",x"391e",x"2cd4",x"21f4",x"3eec",x"3714",x"bb34",x"b6e6",x"2b2e",x"391f",x"2d20"),
(x"a46c",x"3ec5",x"36eb",x"bbaa",x"3475",x"2c25",x"390b",x"327d",x"a165",x"3ee0",x"36eb",x"bbf4",x"2d6d",x"ac2c",x"3917",x"3210",x"a1bd",x"3ee0",x"3715",x"bbf4",x"2da3",x"2b3e",x"390d",x"31fc"),
(x"a46c",x"3ec5",x"36eb",x"bbaa",x"3475",x"2c25",x"390b",x"327d",x"a3f1",x"3ec4",x"3718",x"bba4",x"33dc",x"313e",x"3900",x"3269",x"a4b5",x"3ec3",x"3715",x"bbb4",x"33e8",x"2ed7",x"3900",x"3276"),
(x"2116",x"3ec2",x"3718",x"23ae",x"ac2f",x"3bfb",x"398f",x"31a9",x"25f4",x"3eb9",x"3714",x"2745",x"ad9b",x"3bf7",x"3997",x"3194",x"a4d5",x"3eb8",x"3715",x"a081",x"ad9e",x"3bf8",x"397f",x"3194"),
(x"94d9",x"3eef",x"3713",x"3405",x"bbbe",x"a393",x"390f",x"2d21",x"9548",x"3ef0",x"36ee",x"34a7",x"bba3",x"ac10",x"390e",x"2cd7",x"9cff",x"3eec",x"36ee",x"3b1d",x"b747",x"2911",x"3909",x"2cda"),
(x"2470",x"3ede",x"36eb",x"3bfd",x"212b",x"29e6",x"391c",x"30c1",x"250d",x"3ec4",x"36eb",x"3b9b",x"34d2",x"2ca7",x"3917",x"3054",x"24de",x"3ec4",x"3717",x"3be8",x"30a2",x"2973",x"390d",x"305d"),
(x"1f13",x"3ef0",x"36ee",x"b188",x"bbe0",x"a53f",x"3917",x"2cd5",x"9548",x"3ef0",x"36ee",x"34a7",x"bba3",x"ac10",x"390e",x"2cd7",x"94d9",x"3eef",x"3713",x"3405",x"bbbe",x"a393",x"390f",x"2d21"),
(x"2029",x"3ec5",x"36eb",x"ba79",x"3840",x"3401",x"38cd",x"2cc1",x"2116",x"3ec2",x"3718",x"ba6d",x"3838",x"3468",x"38c8",x"2d16",x"a069",x"3ec3",x"3718",x"398b",x"396b",x"33db",x"38db",x"2d41"),
(x"a50e",x"3eb9",x"36eb",x"b409",x"bbbc",x"27db",x"3905",x"2ec4",x"a4d5",x"3eb8",x"3715",x"b3c8",x"bbc2",x"235f",x"38fc",x"2ee9",x"25f4",x"3eb9",x"3714",x"2f03",x"bbf3",x"23ef",x"390b",x"3022"),
(x"20c8",x"3ee4",x"3716",x"bbad",x"3434",x"2e8a",x"3928",x"2d1c",x"2019",x"3ee5",x"36eb",x"bb95",x"3495",x"306c",x"3927",x"2cc6",x"21cf",x"3ee8",x"36ee",x"bb7c",x"357c",x"2d58",x"3921",x"2cd1"),
(x"91f4",x"3fd4",x"3716",x"30f9",x"a8af",x"3be5",x"3ba8",x"3b0a",x"1aac",x"3fd4",x"3712",x"342b",x"2e69",x"3bae",x"3ba5",x"3b0a",x"20f7",x"3fcc",x"370e",x"2fd2",x"2717",x"3bef",x"3ba1",x"3b12"),
(x"a03c",x"3fc7",x"36eb",x"bb99",x"3315",x"330d",x"3b44",x"38e9",x"980d",x"3fd7",x"36eb",x"b996",x"395e",x"33ec",x"3b44",x"38e0",x"91f4",x"3fd4",x"3716",x"badd",x"375a",x"334d",x"3b3f",x"38e1"),
(x"8010",x"3f87",x"3714",x"ac39",x"29a5",x"3bf9",x"3bad",x"3b4b",x"a040",x"3f85",x"3713",x"a91b",x"2b55",x"3bfb",x"3bb4",x"3b4c",x"9d28",x"3f8f",x"3712",x"aa69",x"287e",x"3bfc",x"3bb1",x"3b44"),
(x"a34c",x"3f8d",x"3711",x"a481",x"2546",x"3bff",x"3bb8",x"3b46",x"a20d",x"3f91",x"3712",x"2a38",x"ad35",x"3bf6",x"3bb6",x"3b43",x"9ff6",x"3f91",x"3711",x"a994",x"2977",x"3bfc",x"3bb3",x"3b42"),
(x"9d28",x"3f8f",x"3712",x"aa69",x"287e",x"3bfc",x"3bb1",x"3b44",x"a040",x"3f85",x"3713",x"a91b",x"2b55",x"3bfb",x"3bb4",x"3b4c",x"a273",x"3f87",x"3712",x"aa73",x"2a97",x"3bfa",x"3bb7",x"3b4a"),
(x"9c36",x"3f82",x"3718",x"ae36",x"a160",x"3bf6",x"3bb0",x"3b4f",x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53",x"a17b",x"3f81",x"3711",x"afec",x"ac2c",x"3beb",x"3bb6",x"3b4f"),
(x"a035",x"3f6a",x"3713",x"ae9c",x"3366",x"3bbd",x"3bb5",x"3b64",x"a289",x"3f6b",x"370f",x"9df0",x"a631",x"3bff",x"3bb9",x"3b62",x"9c56",x"3f71",x"370e",x"26d5",x"25c2",x"3bfe",x"3bb1",x"3b5e"),
(x"9f72",x"3f76",x"3713",x"a538",x"ac79",x"3bfa",x"3bb4",x"3b59",x"9c56",x"3f71",x"370e",x"26d5",x"25c2",x"3bfe",x"3bb1",x"3b5e",x"a289",x"3f6b",x"370f",x"9df0",x"a631",x"3bff",x"3bb9",x"3b62"),
(x"a407",x"3f79",x"370f",x"aec5",x"1a59",x"3bf4",x"3bba",x"3b56",x"9f87",x"3f78",x"3713",x"a7e9",x"2849",x"3bfd",x"3bb4",x"3b58",x"9f72",x"3f76",x"3713",x"a538",x"ac79",x"3bfa",x"3bb4",x"3b59"),
(x"9f87",x"3f78",x"3713",x"a7e9",x"2849",x"3bfd",x"3bb4",x"3b58",x"a407",x"3f79",x"370f",x"aec5",x"1a59",x"3bf4",x"3bba",x"3b56",x"a17b",x"3f81",x"3711",x"afec",x"ac2c",x"3beb",x"3bb6",x"3b4f"),
(x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53",x"9476",x"3f7b",x"3713",x"25b5",x"b7de",x"3af6",x"3bae",x"3b55",x"9d1a",x"3f7a",x"3710",x"ac5b",x"b0a5",x"3be5",x"3bb1",x"3b56"),
(x"9d1a",x"3f7a",x"3710",x"ac5b",x"b0a5",x"3be5",x"3bb1",x"3b56",x"9f87",x"3f78",x"3713",x"a7e9",x"2849",x"3bfd",x"3bb4",x"3b58",x"a17b",x"3f81",x"3711",x"afec",x"ac2c",x"3beb",x"3bb6",x"3b4f"),
(x"1e77",x"3f4b",x"3715",x"a6c2",x"ac63",x"3bfa",x"3ba8",x"3b7e",x"990c",x"3f4b",x"3712",x"af67",x"a981",x"3bf0",x"3baf",x"3b7e",x"19fe",x"3f52",x"3717",x"aff2",x"aa7d",x"3bed",x"3bab",x"3b78"),
(x"a38f",x"3f55",x"3712",x"b163",x"a345",x"3be2",x"3bb9",x"3b75",x"a2d9",x"3f59",x"3714",x"a860",x"af8b",x"3bf0",x"3bb8",x"3b72",x"a13d",x"3f5b",x"3716",x"acd8",x"a7e2",x"3bf9",x"3bb5",x"3b70"),
(x"9e62",x"3f5a",x"3716",x"2818",x"ad04",x"3bf8",x"3bb2",x"3b71",x"9d1e",x"3f4e",x"3711",x"240b",x"ad5c",x"3bf8",x"3bb1",x"3b7b",x"a2cb",x"3f51",x"3714",x"1553",x"ab62",x"3bfc",x"3bb8",x"3b78"),
(x"9d1e",x"3f4e",x"3711",x"240b",x"ad5c",x"3bf8",x"3bb1",x"3b7b",x"987a",x"3f57",x"3714",x"a4fd",x"ada9",x"3bf7",x"3baf",x"3b74",x"0e53",x"3f54",x"3714",x"b036",x"a73e",x"3bed",x"3bad",x"3b76"),
(x"19fe",x"3f52",x"3717",x"aff2",x"aa7d",x"3bed",x"3bab",x"3b78",x"990c",x"3f4b",x"3712",x"af67",x"a981",x"3bf0",x"3baf",x"3b7e",x"9a71",x"3f4c",x"3711",x"b27d",x"16f6",x"3bd5",x"3bb0",x"3b7c"),
(x"9a71",x"3f4c",x"3711",x"b27d",x"16f6",x"3bd5",x"3bb0",x"3b7c",x"9d1e",x"3f4e",x"3711",x"240b",x"ad5c",x"3bf8",x"3bb1",x"3b7b",x"0e53",x"3f54",x"3714",x"b036",x"a73e",x"3bed",x"3bad",x"3b76"),
(x"9ae8",x"3f45",x"3712",x"b146",x"2c91",x"3bde",x"3bb0",x"3b82",x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f"),
(x"1f1f",x"3f39",x"3718",x"2138",x"ae95",x"3bf4",x"3ba8",x"3b8c",x"21d8",x"3f39",x"3719",x"a3bb",x"27ae",x"3bfe",x"3ba5",x"3b8c",x"21e0",x"3f38",x"3719",x"a90e",x"af00",x"3bf2",x"3ba5",x"3b8d"),
(x"1e5a",x"3f3a",x"3718",x"2b4f",x"2525",x"3bfc",x"3ba9",x"3b8b",x"1f1f",x"3f39",x"3718",x"2138",x"ae95",x"3bf4",x"3ba8",x"3b8c",x"8dee",x"3f36",x"3718",x"ae3b",x"1fae",x"3bf6",x"3bae",x"3b8f"),
(x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"20ca",x"3f3e",x"3715",x"2d65",x"ac5a",x"3bf3",x"3ba6",x"3b89",x"1e5a",x"3f3a",x"3718",x"2b4f",x"2525",x"3bfc",x"3ba9",x"3b8b"),
(x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"2091",x"3f49",x"3717",x"2d2f",x"2ecb",x"3bed",x"3ba6",x"3b80",x"2288",x"3f43",x"3718",x"2cf2",x"18ea",x"3bf9",x"3ba3",x"3b85"),
(x"22dc",x"3f47",x"3712",x"359c",x"336a",x"3b42",x"3ba3",x"3b81",x"2288",x"3f43",x"3718",x"2cf2",x"18ea",x"3bf9",x"3ba3",x"3b85",x"2091",x"3f49",x"3717",x"2d2f",x"2ecb",x"3bed",x"3ba6",x"3b80"),
(x"1b8e",x"3f42",x"3718",x"abb4",x"28d3",x"3bfa",x"3bab",x"3b85",x"9ae8",x"3f45",x"3712",x"b146",x"2c91",x"3bde",x"3bb0",x"3b82",x"1f4b",x"3f49",x"3716",x"b009",x"2da6",x"3be7",x"3ba8",x"3b7f"),
(x"1f4b",x"3f49",x"3716",x"b009",x"2da6",x"3be7",x"3ba8",x"3b7f",x"9ae8",x"3f45",x"3712",x"b146",x"2c91",x"3bde",x"3bb0",x"3b82",x"990c",x"3f4b",x"3712",x"af67",x"a981",x"3bf0",x"3baf",x"3b7e"),
(x"1d4c",x"3f53",x"3717",x"97c8",x"9f79",x"3c00",x"3ba9",x"3b76",x"2147",x"3f51",x"3718",x"ac00",x"290e",x"3bfa",x"3ba5",x"3b79",x"1f29",x"3f4d",x"3714",x"a57a",x"ae8a",x"3bf4",x"3ba8",x"3b7c"),
(x"1d4c",x"3f53",x"3717",x"97c8",x"9f79",x"3c00",x"3ba9",x"3b76",x"20ef",x"3f58",x"3715",x"a51e",x"2d06",x"3bf9",x"3ba6",x"3b73",x"2147",x"3f51",x"3718",x"ac00",x"290e",x"3bfa",x"3ba5",x"3b79"),
(x"20ef",x"3f58",x"3715",x"a51e",x"2d06",x"3bf9",x"3ba6",x"3b73",x"2308",x"3f60",x"3714",x"2dba",x"2266",x"3bf7",x"3ba3",x"3b6c",x"2442",x"3f5d",x"3714",x"175f",x"2c2c",x"3bfb",x"3ba0",x"3b6f"),
(x"2308",x"3f60",x"3714",x"2dba",x"2266",x"3bf7",x"3ba3",x"3b6c",x"2365",x"3f6b",x"3715",x"3468",x"247a",x"3bb0",x"3ba2",x"3b63",x"24cc",x"3f69",x"3712",x"3106",x"273e",x"3be5",x"3b9f",x"3b64"),
(x"2365",x"3f6b",x"3715",x"3468",x"247a",x"3bb0",x"3ba2",x"3b63",x"22bc",x"3f73",x"3717",x"3273",x"2f43",x"3bc8",x"3ba3",x"3b5c",x"243c",x"3f75",x"3710",x"3550",x"2e33",x"3b81",x"3ba0",x"3b5a"),
(x"22bc",x"3f73",x"3717",x"3273",x"2f43",x"3bc8",x"3ba3",x"3b5c",x"1f35",x"3f7a",x"3711",x"ae24",x"2a2b",x"3bf4",x"3ba8",x"3b56",x"21ba",x"3f7d",x"3712",x"2b5c",x"2345",x"3bfc",x"3ba5",x"3b54"),
(x"1a19",x"3f7b",x"3712",x"2dd2",x"b04b",x"3be4",x"3bab",x"3b55",x"08f2",x"3f83",x"3716",x"2f4b",x"aa5f",x"3bf0",x"3bad",x"3b4f",x"21ba",x"3f7d",x"3712",x"2b5c",x"2345",x"3bfc",x"3ba5",x"3b54"),
(x"1a19",x"3f7b",x"3712",x"2dd2",x"b04b",x"3be4",x"3bab",x"3b55",x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53",x"08f2",x"3f83",x"3716",x"2f4b",x"aa5f",x"3bf0",x"3bad",x"3b4f"),
(x"1a19",x"3f7b",x"3712",x"2dd2",x"b04b",x"3be4",x"3bab",x"3b55",x"9476",x"3f7b",x"3713",x"25b5",x"b7de",x"3af6",x"3bae",x"3b55",x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53"),
(x"08f2",x"3f83",x"3716",x"2f4b",x"aa5f",x"3bf0",x"3bad",x"3b4f",x"91dd",x"3f7e",x"3718",x"ac13",x"b1c4",x"3bda",x"3bae",x"3b53",x"9c36",x"3f82",x"3718",x"ae36",x"a160",x"3bf6",x"3bb0",x"3b4f"),
(x"9e8d",x"3f84",x"3716",x"af14",x"329b",x"3bc7",x"3bb2",x"3b4e",x"8010",x"3f87",x"3714",x"ac39",x"29a5",x"3bf9",x"3bad",x"3b4b",x"9588",x"3f84",x"3716",x"a559",x"32c7",x"3bd1",x"3bae",x"3b4d"),
(x"9e8d",x"3f84",x"3716",x"af14",x"329b",x"3bc7",x"3bb2",x"3b4e",x"a040",x"3f85",x"3713",x"a91b",x"2b55",x"3bfb",x"3bb4",x"3b4c",x"8010",x"3f87",x"3714",x"ac39",x"29a5",x"3bf9",x"3bad",x"3b4b"),
(x"9a85",x"3f8f",x"3713",x"ada3",x"2f15",x"3beb",x"3baf",x"3b45",x"1820",x"3f93",x"370f",x"aedc",x"2cd0",x"3bee",x"3bab",x"3b41",x"1f40",x"3f8e",x"3717",x"b0e7",x"3057",x"3bd4",x"3ba7",x"3b45"),
(x"1820",x"3f93",x"370f",x"aedc",x"2cd0",x"3bee",x"3bab",x"3b41",x"1d56",x"3f9e",x"3716",x"aadf",x"a6b5",x"3bfc",x"3ba8",x"3b38",x"221f",x"3f9c",x"3713",x"a9b8",x"a6e9",x"3bfd",x"3ba3",x"3b3a"),
(x"2312",x"3fb8",x"370d",x"3809",x"2e09",x"3add",x"3b9f",x"3b23",x"2386",x"3fb5",x"370f",x"36ca",x"2fac",x"3b2e",x"3b9e",x"3b26",x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21"),
(x"21a5",x"3fc1",x"3712",x"29f0",x"2b1d",x"3bfa",x"3ba1",x"3b1b",x"9cbb",x"3fba",x"3715",x"19bc",x"a6cf",x"3bff",x"3bae",x"3b20",x"9df1",x"3fc7",x"3715",x"2d56",x"20d0",x"3bf8",x"3bad",x"3b15"),
(x"1882",x"3fa8",x"370e",x"bb5f",x"b5f1",x"2f4f",x"3b3c",x"38f9",x"1737",x"3fa7",x"36eb",x"bb4a",x"b677",x"2cfa",x"3b40",x"38fa",x"9f02",x"3fb9",x"36eb",x"bb89",x"b473",x"31fc",x"3b43",x"38f0"),
(x"a175",x"3f1a",x"3710",x"3bfd",x"a997",x"a0a8",x"3b8a",x"3a03",x"a0d2",x"3f23",x"3713",x"3ba5",x"b497",x"ac28",x"3b8a",x"39fe",x"a122",x"3f23",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3b85",x"39fe"),
(x"a167",x"3f14",x"36eb",x"3bf5",x"2e59",x"2467",x"3b86",x"3a06",x"a140",x"3f12",x"3714",x"3beb",x"308b",x"98b5",x"3b8b",x"3a07",x"a175",x"3f1a",x"3710",x"3bfd",x"a997",x"a0a8",x"3b8a",x"3a03"),
(x"9c3a",x"3f30",x"3714",x"3b1c",x"b754",x"223f",x"3b8a",x"39f7",x"8dee",x"3f36",x"3718",x"b9e5",x"b968",x"0000",x"3b8b",x"39f3",x"8dee",x"3f36",x"36eb",x"b469",x"bb91",x"316a",x"3b85",x"39f3"),
(x"a122",x"3f23",x"36eb",x"3ba1",x"b4cc",x"1f45",x"3b85",x"39fe",x"a0d2",x"3f23",x"3713",x"3ba5",x"b497",x"ac28",x"3b8a",x"39fe",x"9c3a",x"3f30",x"3714",x"3b1c",x"b754",x"223f",x"3b8a",x"39f7"),
(x"a099",x"3f0e",x"3712",x"3b76",x"35c5",x"204d",x"3b8a",x"3a09",x"a140",x"3f12",x"3714",x"3beb",x"308b",x"98b5",x"3b8b",x"3a07",x"a167",x"3f14",x"36eb",x"3bf5",x"2e59",x"2467",x"3b86",x"3a06"),
(x"a051",x"3f0c",x"36eb",x"3ab1",x"3862",x"21e3",x"3b86",x"3a0a",x"9ecc",x"3f0b",x"3714",x"395a",x"39f1",x"2025",x"3b8b",x"3a0b",x"a099",x"3f0e",x"3712",x"3b76",x"35c5",x"204d",x"3b8a",x"3a09"),
(x"9b3f",x"3f08",x"36eb",x"37e1",x"3af5",x"269a",x"3b86",x"3a0d",x"9aa8",x"3f08",x"3714",x"35bf",x"3b76",x"27db",x"3b8b",x"3a0d",x"9ecc",x"3f0b",x"3714",x"395a",x"39f1",x"2025",x"3b8b",x"3a0b"),
(x"197e",x"3f07",x"36eb",x"303c",x"3beb",x"299e",x"3b86",x"3a11",x"1a1e",x"3f06",x"3715",x"a836",x"3bfd",x"294f",x"3b8b",x"3a11",x"9aa8",x"3f08",x"3714",x"35bf",x"3b76",x"27db",x"3b8b",x"3a0d"),
(x"20a0",x"3f08",x"36eb",x"b868",x"3aab",x"296a",x"3b86",x"3a14",x"20b2",x"3f08",x"3716",x"b86f",x"3aa7",x"2604",x"3b8b",x"3a14",x"1a1e",x"3f06",x"3715",x"a836",x"3bfd",x"294f",x"3b8b",x"3a11"),
(x"20a0",x"3f08",x"36eb",x"b868",x"3aab",x"296a",x"3b86",x"3a14",x"2300",x"3f0e",x"36eb",x"baf3",x"37df",x"2b38",x"3b86",x"3a18",x"2335",x"3f0e",x"3714",x"bb01",x"37b5",x"2839",x"3b8b",x"3a18"),
(x"23d0",x"3f13",x"36eb",x"bbf9",x"2d11",x"2511",x"3b85",x"3a1b",x"23d3",x"3f13",x"3714",x"bbe6",x"b10f",x"9bfc",x"3b8b",x"3a1b",x"2335",x"3f0e",x"3714",x"bb01",x"37b5",x"2839",x"3b8b",x"3a18"),
(x"2300",x"3f18",x"36eb",x"b90c",x"ba34",x"2532",x"3b85",x"3a1e",x"22d3",x"3f18",x"3715",x"b928",x"ba1d",x"1553",x"3b8b",x"3a1e",x"23d3",x"3f13",x"3714",x"bbe6",x"b10f",x"9bfc",x"3b8b",x"3a1b"),
(x"2300",x"3f18",x"36eb",x"b90c",x"ba34",x"2532",x"3a68",x"3a42",x"20b2",x"3f18",x"36eb",x"35dd",x"bb6d",x"2be9",x"3a68",x"3a3f",x"20d5",x"3f18",x"3714",x"2fe4",x"bbee",x"2901",x"3a63",x"3a3f"),
(x"20b2",x"3f18",x"36eb",x"35dd",x"bb6d",x"2be9",x"3a68",x"3a3f",x"1ead",x"3f15",x"36eb",x"32b1",x"bbc8",x"2e54",x"3a68",x"3a3d",x"1e4f",x"3f16",x"3711",x"364f",x"bb52",x"2d1b",x"3a64",x"3a3d"),
(x"13e1",x"3f25",x"36eb",x"bbf6",x"2a70",x"2d61",x"3a69",x"3a31",x"15a0",x"3f25",x"3713",x"bbc2",x"33a4",x"298a",x"3a64",x"3a32",x"3d81",x"3f23",x"3711",x"ba7a",x"38b0",x"2839",x"3a64",x"3a33"),
(x"1ead",x"3f15",x"36eb",x"32b1",x"bbc8",x"2e54",x"3a68",x"3a3d",x"0f13",x"3f15",x"36eb",x"b37e",x"bbba",x"2ef6",x"3a69",x"3a3a",x"14bb",x"3f16",x"3710",x"b416",x"bbad",x"2f8d",x"3a64",x"3a3b"),
(x"9f83",x"3f68",x"36eb",x"35e4",x"bb4d",x"31a2",x"3b2b",x"3927",x"a035",x"3f6a",x"3713",x"3583",x"bb63",x"3153",x"3b29",x"3922",x"9c14",x"3f6f",x"370f",x"3a9b",x"b854",x"30fa",x"3b26",x"3924"),
(x"9f02",x"3fb9",x"36eb",x"bb89",x"b473",x"31fc",x"3b43",x"38f0",x"a03c",x"3fc7",x"36eb",x"bb99",x"3315",x"330d",x"3b44",x"38e9",x"9df1",x"3fc7",x"3715",x"bbc5",x"2b9a",x"3358",x"3b3e",x"38e9"),
(x"983c",x"3f20",x"3710",x"a856",x"a9ab",x"3bfc",x"3bb0",x"3ba1",x"3d81",x"3f23",x"3711",x"b40c",x"26bb",x"3bbc",x"3bae",x"3b9f",x"1f0f",x"3f25",x"3718",x"ab65",x"b528",x"3b8f",x"3ba8",x"3b9d"),
(x"210e",x"3fbb",x"36eb",x"3be3",x"2ce8",x"30c3",x"3b3c",x"38cf",x"21a5",x"3fc1",x"3712",x"3bcf",x"b081",x"3141",x"3b3a",x"38d5",x"229f",x"3fc1",x"36eb",x"3bdb",x"1c67",x"320a",x"3b3e",x"38d2"),
(x"210e",x"3fbb",x"36eb",x"3be3",x"2ce8",x"30c3",x"3b3c",x"38cf",x"20d5",x"3fbc",x"3715",x"3bd7",x"b1f9",x"2c2a",x"3b38",x"38d3",x"21a5",x"3fc1",x"3712",x"3bcf",x"b081",x"3141",x"3b3a",x"38d5"),
(x"2267",x"3f7e",x"36eb",x"3958",x"39de",x"2fdf",x"3b35",x"3b43",x"2469",x"3f76",x"36eb",x"3b75",x"35a2",x"2d46",x"3b35",x"3b3e",x"243c",x"3f75",x"3710",x"3b6a",x"35bb",x"2efe",x"3b31",x"3b3e"),
(x"9889",x"3f18",x"36eb",x"baa4",x"b859",x"2fe5",x"3a69",x"3a38",x"951c",x"3f19",x"3711",x"ba7e",x"b887",x"3089",x"3a64",x"3a39",x"14bb",x"3f16",x"3710",x"b416",x"bbad",x"2f8d",x"3a64",x"3a3b"),
(x"1e52",x"3f28",x"36eb",x"3be6",x"308f",x"2c41",x"3a31",x"3a5e",x"1d9c",x"3f28",x"3718",x"3be6",x"309e",x"2baa",x"3a2c",x"3a5c",x"1d4f",x"3f31",x"3715",x"3bfa",x"a710",x"2c48",x"3a2b",x"3a61"),
(x"9889",x"3f18",x"36eb",x"baa4",x"b859",x"2fe5",x"3a69",x"3a38",x"9b9c",x"3f1c",x"36eb",x"bbf4",x"9edc",x"2ebb",x"3a69",x"3a36",x"99ac",x"3f1c",x"3710",x"bbcc",x"b228",x"2f2f",x"3a64",x"3a37"),
(x"998f",x"3f6e",x"36eb",x"3b7d",x"b521",x"3095",x"3b28",x"3928",x"9c14",x"3f6f",x"370f",x"3a9b",x"b854",x"30fa",x"3b26",x"3924",x"9c56",x"3f71",x"370e",x"3b25",x"370d",x"2d68",x"3b25",x"3924"),
(x"a30f",x"3f4f",x"36eb",x"b6fe",x"bb25",x"2ea4",x"3b1f",x"3b1f",x"a2cb",x"3f51",x"3714",x"b972",x"b9bb",x"30de",x"3b1a",x"3b1d",x"9d1e",x"3f4e",x"3711",x"b4dc",x"bb97",x"2d61",x"3b19",x"3b22"),
(x"865b",x"3f23",x"36eb",x"b9db",x"396c",x"2c1a",x"3a69",x"3a32",x"3d81",x"3f23",x"3711",x"ba7a",x"38b0",x"2839",x"3a64",x"3a33",x"983c",x"3f20",x"3710",x"bb2f",x"36d9",x"2e52",x"3a64",x"3a35"),
(x"8d14",x"3f84",x"36eb",x"3776",x"3b0b",x"2d41",x"3b34",x"3b4b",x"2267",x"3f7e",x"36eb",x"3958",x"39de",x"2fdf",x"3b35",x"3b43",x"21ba",x"3f7d",x"3712",x"384e",x"3ab0",x"2ec8",x"3b30",x"3b43"),
(x"1e6c",x"3f33",x"36eb",x"39df",x"b964",x"2d28",x"3a2f",x"3a63",x"1e18",x"3f31",x"36eb",x"3bfa",x"a0b5",x"2cb4",x"3a30",x"3a63",x"1d4f",x"3f31",x"3715",x"3bfa",x"a710",x"2c48",x"3a2b",x"3a61"),
(x"9f02",x"3f76",x"36eb",x"3ad3",x"3822",x"2c4d",x"3b24",x"392a",x"9aca",x"3f71",x"36eb",x"3b19",x"3744",x"2cf7",x"3b27",x"3929",x"9c56",x"3f71",x"370e",x"3b25",x"370d",x"2d68",x"3b25",x"3924"),
(x"1d3a",x"3f9d",x"36eb",x"bbfe",x"1e8d",x"2828",x"3b3f",x"3900",x"1737",x"3fa7",x"36eb",x"bb4a",x"b677",x"2cfa",x"3b40",x"38fa",x"1882",x"3fa8",x"370e",x"bb5f",x"b5f1",x"2f4f",x"3b3c",x"38f9"),
(x"8d14",x"3f84",x"36eb",x"3776",x"3b0b",x"2d41",x"3b34",x"3b4b",x"08f2",x"3f83",x"3716",x"37e9",x"3af1",x"2aa7",x"3b2f",x"3b4a",x"9588",x"3f84",x"3716",x"3bde",x"31b5",x"2825",x"3b2e",x"3b4b"),
(x"22d4",x"3f38",x"36eb",x"39ed",x"b94b",x"2f45",x"3a2e",x"3a68",x"1e6c",x"3f33",x"36eb",x"39df",x"b964",x"2d28",x"3a2f",x"3a63",x"1e3f",x"3f34",x"3715",x"395d",x"b9e3",x"2de3",x"3a2a",x"3a62"),
(x"9a71",x"3f4c",x"3711",x"bb12",x"b763",x"2ca3",x"3a28",x"3a14",x"990c",x"3f4b",x"3712",x"bbf7",x"283f",x"2d8f",x"3a28",x"3a15",x"9acb",x"3f4a",x"36eb",x"bbf8",x"a379",x"2d44",x"3a2d",x"3a14"),
(x"9c70",x"3f4d",x"36eb",x"b7d8",x"baf6",x"2a35",x"3a2c",x"3a12",x"9d1e",x"3f4e",x"3711",x"b4dc",x"bb97",x"2d61",x"3a28",x"3a13",x"9a71",x"3f4c",x"3711",x"bb12",x"b763",x"2ca3",x"3a28",x"3a14"),
(x"9f11",x"3f77",x"36eb",x"39e9",x"b955",x"2e31",x"3b23",x"392a",x"9f02",x"3f76",x"36eb",x"3ad3",x"3822",x"2c4d",x"3b24",x"392a",x"9f72",x"3f76",x"3713",x"3b5b",x"3634",x"2c03",x"3b22",x"3925"),
(x"1d3a",x"3f9d",x"36eb",x"bbfe",x"1e8d",x"2828",x"3b3f",x"3900",x"1d56",x"3f9e",x"3716",x"bbff",x"20c2",x"2138",x"3b3a",x"38ff",x"1820",x"3f93",x"370f",x"bad7",x"3821",x"29e6",x"3b3a",x"3904"),
(x"9427",x"3f84",x"36eb",x"3b23",x"b71d",x"2cde",x"3b25",x"38b9",x"9588",x"3f84",x"3716",x"3bde",x"31b5",x"2825",x"3b21",x"38bd",x"8010",x"3f87",x"3714",x"39e8",x"b951",x"2f27",x"3b23",x"38be"),
(x"22d4",x"3f38",x"36eb",x"39ed",x"b94b",x"2f45",x"3a2e",x"3a68",x"21e0",x"3f38",x"3719",x"39a6",x"b994",x"2fc6",x"3a29",x"3a66",x"21d8",x"3f39",x"3719",x"3250",x"3bca",x"2f22",x"3a29",x"3a66"),
(x"9acb",x"3f4a",x"36eb",x"bbf8",x"a379",x"2d44",x"3a2d",x"3a14",x"990c",x"3f4b",x"3712",x"bbf7",x"283f",x"2d8f",x"3a28",x"3a15",x"9ae8",x"3f45",x"3712",x"bb92",x"3509",x"2cb0",x"3a29",x"3a18"),
(x"9d1a",x"3f7a",x"3710",x"3833",x"bac7",x"2d1d",x"3b1b",x"3aef",x"9476",x"3f7b",x"3713",x"30a8",x"bbe9",x"22dc",x"3b1a",x"3af1",x"9096",x"3f7b",x"36eb",x"3046",x"bbe8",x"2cb7",x"3b1f",x"3af2"),
(x"9f11",x"3f77",x"36eb",x"39e9",x"b955",x"2e31",x"3b1f",x"3aee",x"9f87",x"3f78",x"3713",x"3b09",x"b791",x"2ab8",x"3b1a",x"3aed",x"9d1a",x"3f7a",x"3710",x"3833",x"bac7",x"2d1d",x"3b1b",x"3aef"),
(x"9bdf",x"3f8f",x"36eb",x"b73f",x"3b1a",x"2d3c",x"3b3e",x"3909",x"173f",x"3f94",x"36eb",x"bab4",x"3859",x"2a66",x"3b3e",x"3905",x"1820",x"3f93",x"370f",x"bad7",x"3821",x"29e6",x"3b3a",x"3904"),
(x"141e",x"3f86",x"36eb",x"397a",x"b9b6",x"309a",x"3b26",x"38b9",x"8010",x"3f87",x"3714",x"39e8",x"b951",x"2f27",x"3b23",x"38be",x"1f40",x"3f8e",x"3717",x"3a77",x"b889",x"310e",x"3b27",x"38c1"),
(x"1e72",x"3f3a",x"36eb",x"3b01",x"3745",x"3141",x"3a2c",x"3a6c",x"2283",x"3f3b",x"36eb",x"32cb",x"3bc1",x"2fc5",x"3a2e",x"3a69",x"21d8",x"3f39",x"3719",x"3250",x"3bca",x"2f22",x"3a29",x"3a66"),
(x"9bea",x"3f46",x"36eb",x"bb57",x"3625",x"2e99",x"3a2d",x"3a16",x"9ae8",x"3f45",x"3712",x"bb92",x"3509",x"2cb0",x"3a29",x"3a18",x"a16d",x"3f34",x"3711",x"bb70",x"3585",x"3014",x"3a2c",x"3a21"),
(x"1a19",x"3f7b",x"3712",x"b2e8",x"bbcb",x"2c10",x"3b1a",x"3af3",x"1f35",x"3f7a",x"3711",x"b934",x"ba0d",x"2c16",x"3b1a",x"3af5",x"1ecc",x"3f79",x"36eb",x"b74a",x"bb15",x"2de4",x"3b1f",x"3af6"),
(x"9096",x"3f7b",x"36eb",x"3046",x"bbe8",x"2cb7",x"3b1f",x"3af2",x"9476",x"3f7b",x"3713",x"30a8",x"bbe9",x"22dc",x"3b1a",x"3af1",x"1a19",x"3f7b",x"3712",x"b2e8",x"bbcb",x"2c10",x"3b1a",x"3af3"),
(x"9bdf",x"3f8f",x"36eb",x"b73f",x"3b1a",x"2d3c",x"3b3e",x"3909",x"9a85",x"3f8f",x"3713",x"b7c3",x"3af3",x"2e28",x"3b39",x"3908",x"9d28",x"3f8f",x"3712",x"3721",x"3b24",x"2bf9",x"3b39",x"3909"),
(x"2078",x"3f8e",x"36eb",x"3aff",x"b73c",x"3197",x"3b2a",x"38bd",x"1f40",x"3f8e",x"3717",x"3a77",x"b889",x"310e",x"3b27",x"38c1",x"221f",x"3f9c",x"3713",x"3bc6",x"b1be",x"30de",x"3b2c",x"38c6"),
(x"a25f",x"3f33",x"36eb",x"bb99",x"345f",x"30d6",x"3a30",x"3a21",x"a16d",x"3f34",x"3711",x"bb70",x"3585",x"3014",x"3a2c",x"3a21",x"a2e9",x"3f24",x"3711",x"bbe4",x"2d1d",x"308c",x"3a2e",x"3a2a"),
(x"2284",x"3f73",x"36eb",x"baaf",x"b860",x"2a70",x"3b1f",x"3afa",x"1ecc",x"3f79",x"36eb",x"b74a",x"bb15",x"2de4",x"3b1f",x"3af6",x"1f35",x"3f7a",x"3711",x"b934",x"ba0d",x"2c16",x"3b1a",x"3af5"),
(x"9d97",x"3f90",x"36eb",x"38ae",x"3a73",x"2d47",x"3b3d",x"390a",x"9d28",x"3f8f",x"3712",x"3721",x"3b24",x"2bf9",x"3b39",x"3909",x"9ff6",x"3f91",x"3711",x"35dd",x"3b65",x"2eae",x"3b39",x"390b"),
(x"22be",x"3fa9",x"36eb",x"3bea",x"ae0a",x"2f10",x"3b35",x"38c7",x"231e",x"3f9c",x"36eb",x"3bbf",x"b113",x"322d",x"3b30",x"38c2",x"221f",x"3f9c",x"3713",x"3bc6",x"b1be",x"30de",x"3b2c",x"38c6"),
(x"1e72",x"3f3a",x"36eb",x"3b01",x"3745",x"3141",x"3b34",x"3b18",x"20ca",x"3f3e",x"3715",x"39d1",x"b974",x"2cc6",x"3b2f",x"3b1c",x"21d1",x"3f3e",x"36eb",x"3a0e",x"b929",x"2e76",x"3b35",x"3b1c"),
(x"1e72",x"3f3a",x"36eb",x"3b01",x"3745",x"3141",x"3b34",x"3b18",x"1e5a",x"3f3a",x"3718",x"3af6",x"b7e0",x"2460",x"3b2f",x"3b1a",x"20ca",x"3f3e",x"3715",x"39d1",x"b974",x"2cc6",x"3b2f",x"3b1c"),
(x"a382",x"3f13",x"36eb",x"bbe8",x"ad68",x"3010",x"3a34",x"3a31",x"a397",x"3f24",x"36eb",x"bbe6",x"2c77",x"308c",x"3a32",x"3a28",x"a2e9",x"3f24",x"3711",x"bbe4",x"2d1d",x"308c",x"3a2e",x"3a2a"),
(x"234c",x"3f6b",x"36eb",x"bbfa",x"ac62",x"2617",x"3b1f",x"3afe",x"2284",x"3f73",x"36eb",x"baaf",x"b860",x"2a70",x"3b1f",x"3afa",x"22bc",x"3f73",x"3717",x"bb6f",x"b5e5",x"261e",x"3b19",x"3afa"),
(x"9f8c",x"3f92",x"36eb",x"2e29",x"3be6",x"3005",x"3b3d",x"390b",x"9ff6",x"3f91",x"3711",x"35dd",x"3b65",x"2eae",x"3b39",x"390b",x"a20d",x"3f91",x"3712",x"b5a5",x"3b63",x"30cc",x"3b38",x"390d"),
(x"22be",x"3fa9",x"36eb",x"3bea",x"ae0a",x"2f10",x"3b35",x"38c7",x"2273",x"3faa",x"3717",x"3bf0",x"af10",x"2aec",x"3b31",x"38cb",x"2386",x"3fb5",x"370f",x"3bdd",x"b0de",x"2e6c",x"3b36",x"38ce"),
(x"21d1",x"3f3e",x"36eb",x"3a0e",x"b929",x"2e76",x"3b35",x"3b1c",x"20ca",x"3f3e",x"3715",x"39d1",x"b974",x"2cc6",x"3b2f",x"3b1c",x"2288",x"3f43",x"3718",x"3b13",x"b732",x"2fec",x"3b2f",x"3b1f"),
(x"a382",x"3f13",x"36eb",x"bbe8",x"ad68",x"3010",x"3a34",x"3a31",x"a2ee",x"3f13",x"3714",x"bbec",x"ad02",x"2f4a",x"3a2f",x"3a32",x"a1ea",x"3f0b",x"3712",x"bb45",x"b640",x"30a6",x"3a30",x"3a36"),
(x"9b9c",x"3f1c",x"36eb",x"bbf4",x"9edc",x"2ebb",x"3a69",x"3a36",x"9a2a",x"3f21",x"36eb",x"bb02",x"3776",x"2fc8",x"3a69",x"3a34",x"983c",x"3f20",x"3710",x"bb2f",x"36d9",x"2e52",x"3a64",x"3a35"),
(x"22be",x"3f61",x"36eb",x"bbcf",x"32aa",x"2bc5",x"3b1e",x"3b04",x"234c",x"3f6b",x"36eb",x"bbfa",x"ac62",x"2617",x"3b1f",x"3afe",x"2365",x"3f6b",x"3715",x"bbfe",x"2412",x"2867",x"3b19",x"3aff"),
(x"a2ba",x"3f92",x"36eb",x"b913",x"3a0d",x"310f",x"3b3d",x"390e",x"a20d",x"3f91",x"3712",x"b5a5",x"3b63",x"30cc",x"3b38",x"390d",x"a34c",x"3f8d",x"3711",x"bbb2",x"332f",x"30f4",x"3b38",x"390f"),
(x"2414",x"3fb4",x"36eb",x"3be4",x"aadf",x"30ee",x"3b39",x"38ca",x"2386",x"3fb5",x"370f",x"3bdd",x"b0de",x"2e6c",x"3b36",x"38ce",x"2312",x"3fb8",x"370d",x"3b0d",x"370c",x"3169",x"3b37",x"38cf"),
(x"2349",x"3f43",x"36eb",x"3bbf",x"b333",x"2ed0",x"3b35",x"3b1f",x"2288",x"3f43",x"3718",x"3b13",x"b732",x"2fec",x"3b2f",x"3b1f",x"22dc",x"3f47",x"3712",x"3bf0",x"2c20",x"2e95",x"3b30",x"3b22"),
(x"a269",x"3f0a",x"36eb",x"bab2",x"b834",x"30cb",x"3a35",x"3a36",x"a1ea",x"3f0b",x"3712",x"bb45",x"b640",x"30a6",x"3a30",x"3a36",x"9d7f",x"3f04",x"3715",x"b93c",x"b9e9",x"3110",x"3a31",x"3a3c"),
(x"207d",x"3f59",x"36eb",x"bac2",x"3833",x"2e8a",x"3b1f",x"3b09",x"22be",x"3f61",x"36eb",x"bbcf",x"32aa",x"2bc5",x"3b1e",x"3b04",x"2308",x"3f60",x"3714",x"bb81",x"3558",x"2da5",x"3b19",x"3b04"),
(x"a3f7",x"3f8d",x"36eb",x"bbe5",x"adbc",x"3036",x"3b3c",x"3911",x"a34c",x"3f8d",x"3711",x"bbb2",x"332f",x"30f4",x"3b38",x"390f",x"a273",x"3f87",x"3712",x"bae4",x"b7c3",x"30c9",x"3b36",x"3912"),
(x"226e",x"3fbb",x"36eb",x"3571",x"3b6d",x"30cc",x"3b3b",x"38ce",x"23bf",x"3fba",x"36eb",x"3af6",x"3714",x"32f0",x"3b3b",x"38cd",x"2312",x"3fb8",x"370d",x"3b0d",x"370c",x"3169",x"3b37",x"38cf"),
(x"2324",x"3f48",x"36eb",x"3bbf",x"3371",x"2dad",x"3b35",x"3b21",x"22dc",x"3f47",x"3712",x"3bf0",x"2c20",x"2e95",x"3b30",x"3b22",x"2257",x"3f49",x"3712",x"3297",x"3bcc",x"2d84",x"3b30",x"3b23"),
(x"9dfd",x"3f02",x"36eb",x"b7cb",x"bae6",x"3068",x"3a36",x"3a3b",x"9d7f",x"3f04",x"3715",x"b93c",x"b9e9",x"3110",x"3a31",x"3a3c",x"17a2",x"3f01",x"3715",x"9ef6",x"bbee",x"302a",x"3a31",x"3a40"),
(x"1ce6",x"3f54",x"36eb",x"b9cd",x"3979",x"2caa",x"3b1f",x"3b0c",x"207d",x"3f59",x"36eb",x"bac2",x"3833",x"2e8a",x"3b1f",x"3b09",x"20ef",x"3f58",x"3715",x"ba65",x"38c1",x"2d9c",x"3b19",x"3b09"),
(x"a2c3",x"3f85",x"36eb",x"b902",x"ba23",x"306a",x"3b3a",x"3915",x"a273",x"3f87",x"3712",x"bae4",x"b7c3",x"30c9",x"3b36",x"3912",x"a040",x"3f85",x"3713",x"b607",x"bb5e",x"2e4f",x"3b35",x"3914"),
(x"210e",x"3fbb",x"36eb",x"3be3",x"2ce8",x"30c3",x"3b3c",x"38cf",x"226e",x"3fbb",x"36eb",x"3571",x"3b6d",x"30cc",x"3b3b",x"38ce",x"2243",x"3fba",x"3713",x"3451",x"3bac",x"2d81",x"3b37",x"38d1"),
(x"2058",x"3f49",x"36eb",x"2c56",x"3bf7",x"2bc1",x"3b35",x"3b25",x"22c6",x"3f49",x"36eb",x"2eda",x"3bea",x"2e47",x"3b35",x"3b22",x"2257",x"3f49",x"3712",x"3297",x"3bcc",x"2d84",x"3b30",x"3b23"),
(x"20e4",x"3f02",x"36eb",x"366a",x"bb44",x"2f81",x"3a36",x"3a44",x"17aa",x"3f00",x"36eb",x"96f6",x"bbf5",x"2e97",x"3a36",x"3a3f",x"17a2",x"3f01",x"3715",x"9ef6",x"bbee",x"302a",x"3a31",x"3a40"),
(x"1a1b",x"3f52",x"36eb",x"35a6",x"3b74",x"2d53",x"3b1f",x"3b0d",x"1ce6",x"3f54",x"36eb",x"b9cd",x"3979",x"2caa",x"3b1f",x"3b0c",x"1d4c",x"3f53",x"3717",x"b939",x"3a0b",x"29e0",x"3b19",x"3b0c"),
(x"9efd",x"3f84",x"36eb",x"b94d",x"39f2",x"2dc5",x"3b38",x"3918",x"9ff8",x"3f85",x"36eb",x"b3f1",x"bbbc",x"2b5c",x"3b39",x"3917",x"a040",x"3f85",x"3713",x"b607",x"bb5e",x"2e4f",x"3b35",x"3914"),
(x"20d5",x"3fbc",x"3715",x"a587",x"307a",x"3beb",x"3ba2",x"3b1f",x"9cbb",x"3fba",x"3715",x"19bc",x"a6cf",x"3bff",x"3bae",x"3b20",x"21a5",x"3fc1",x"3712",x"29f0",x"2b1d",x"3bfa",x"3ba1",x"3b1b"),
(x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21",x"1882",x"3fa8",x"370e",x"b004",x"a71d",x"3bef",x"3baa",x"3b2f",x"9cbb",x"3fba",x"3715",x"19bc",x"a6cf",x"3bff",x"3bae",x"3b20"),
(x"20f8",x"3fba",x"3716",x"a0ea",x"a780",x"3bfe",x"3ba2",x"3b21",x"9cbb",x"3fba",x"3715",x"19bc",x"a6cf",x"3bff",x"3bae",x"3b20",x"20d5",x"3fbc",x"3715",x"a587",x"307a",x"3beb",x"3ba2",x"3b1f"),
(x"2273",x"3faa",x"3717",x"abf6",x"25ae",x"3bfb",x"3ba1",x"3b2f",x"1d56",x"3f9e",x"3716",x"aadf",x"a6b5",x"3bfc",x"3ba8",x"3b38",x"1882",x"3fa8",x"370e",x"b004",x"a71d",x"3bef",x"3baa",x"3b2f"),
(x"2058",x"3f49",x"36eb",x"2c56",x"3bf7",x"2bc1",x"3b35",x"3b25",x"2091",x"3f49",x"3717",x"2a07",x"3bfc",x"284d",x"3b2f",x"3b24",x"1f4b",x"3f49",x"3716",x"38f4",x"3a42",x"2c09",x"3b30",x"3b25"),
(x"24bd",x"3f09",x"36eb",x"39f2",x"b938",x"30b5",x"3a36",x"3a4a",x"20e4",x"3f02",x"36eb",x"366a",x"bb44",x"2f81",x"3a36",x"3a44",x"210b",x"3f04",x"3713",x"382e",x"baba",x"306c",x"3a31",x"3a44"),
(x"0e53",x"3f54",x"3714",x"39a7",x"399f",x"2d1e",x"3b1a",x"3b0f",x"987a",x"3f57",x"3714",x"397e",x"39c5",x"2dbf",x"3b1a",x"3b12",x"98cf",x"3f58",x"36eb",x"3976",x"39cc",x"2dcc",x"3b1f",x"3b12"),
(x"1a1b",x"3f52",x"36eb",x"35a6",x"3b74",x"2d53",x"3b1f",x"3b0d",x"19fe",x"3f52",x"3717",x"2c95",x"3bf9",x"2918",x"3b19",x"3b0e",x"0e53",x"3f54",x"3714",x"39a7",x"399f",x"2d1e",x"3b1a",x"3b0f"),
(x"9efd",x"3f84",x"36eb",x"b94d",x"39f2",x"2dc5",x"3b38",x"3918",x"9e8d",x"3f84",x"3716",x"bac7",x"383c",x"283f",x"3b34",x"3915",x"a17b",x"3f81",x"3711",x"b8c8",x"3a4e",x"30a8",x"3b33",x"3917"),
(x"2585",x"3f12",x"36eb",x"3bc4",x"b27a",x"3012",x"3a35",x"3a4f",x"24bd",x"3f09",x"36eb",x"39f2",x"b938",x"30b5",x"3a36",x"3a4a",x"2466",x"3f0a",x"3715",x"3ae0",x"b7cf",x"30d4",x"3a31",x"3a49"),
(x"98cf",x"3f58",x"36eb",x"3976",x"39cc",x"2dcc",x"3b1f",x"3b12",x"987a",x"3f57",x"3714",x"397e",x"39c5",x"2dbf",x"3b1a",x"3b12",x"9e62",x"3f5a",x"3716",x"37d5",x"3af0",x"2d8e",x"3b1a",x"3b14"),
(x"a282",x"3f82",x"36eb",x"b9ec",x"392b",x"31e4",x"3b37",x"391b",x"a17b",x"3f81",x"3711",x"b8c8",x"3a4e",x"30a8",x"3b33",x"3917",x"a407",x"3f79",x"370f",x"bb4b",x"35cc",x"3223",x"3b30",x"391b"),
(x"229f",x"3fc1",x"36eb",x"3bdb",x"1c67",x"320a",x"3b3e",x"38d2",x"21a5",x"3fc1",x"3712",x"3bcf",x"b081",x"3141",x"3b3a",x"38d5",x"20f7",x"3fcc",x"370e",x"3b7b",x"34a9",x"3270",x"3b3d",x"38d9"),
(x"1e77",x"3f4b",x"3715",x"3ac2",x"b812",x"3146",x"3b30",x"3b26",x"1f29",x"3f4d",x"3714",x"b879",x"347b",x"3a3d",x"3b2f",x"3b28",x"2147",x"3f51",x"3718",x"3ac6",x"b7dc",x"3286",x"3b2f",x"3b2a"),
(x"255d",x"3f1c",x"36eb",x"3b6e",x"3575",x"309e",x"3a34",x"3a54",x"2585",x"3f12",x"36eb",x"3bc4",x"b27a",x"3012",x"3a35",x"3a4f",x"253f",x"3f13",x"3715",x"3bec",x"abe2",x"2fce",x"3a30",x"3a4e"),
(x"9c3a",x"3f30",x"3714",x"b05e",x"21a1",x"3bec",x"3bb1",x"3b94",x"a2e9",x"3f24",x"3711",x"acd1",x"250b",x"3bf9",x"3bb9",x"3b9d",x"a16d",x"3f34",x"3711",x"b115",x"27d5",x"3be4",x"3bb6",x"3b90"),
(x"9c3a",x"3f30",x"3714",x"b05e",x"21a1",x"3bec",x"3bb1",x"3b94",x"a0d2",x"3f23",x"3713",x"b0f4",x"19bc",x"3be7",x"3bb5",x"3b9f",x"a2e9",x"3f24",x"3711",x"acd1",x"250b",x"3bf9",x"3bb9",x"3b9d"),
(x"9e13",x"3f5b",x"36eb",x"353f",x"3b87",x"2d28",x"3b20",x"3b14",x"9e62",x"3f5a",x"3716",x"37d5",x"3af0",x"2d8e",x"3b1a",x"3b14",x"a13d",x"3f5b",x"3716",x"a345",x"3bf7",x"2dcc",x"3b1a",x"3b17"),
(x"a471",x"3f79",x"36eb",x"bbbc",x"3212",x"3175",x"3b34",x"391f",x"a407",x"3f79",x"370f",x"bb4b",x"35cc",x"3223",x"3b30",x"391b",x"a425",x"3f70",x"370f",x"bbd3",x"af46",x"3182",x"3b2d",x"391f"),
(x"22bc",x"3f52",x"36eb",x"3adb",x"b7e7",x"30ac",x"3b35",x"3b2b",x"2147",x"3f51",x"3718",x"3ac6",x"b7dc",x"3286",x"3b2f",x"3b2a",x"2442",x"3f5d",x"3714",x"3b6b",x"b587",x"3095",x"3b30",x"3b31"),
(x"255d",x"3f1c",x"36eb",x"3b6e",x"3575",x"309e",x"3a34",x"3a54",x"24fc",x"3f1b",x"3717",x"3b55",x"35fd",x"307e",x"3a2f",x"3a53",x"2375",x"3f22",x"3711",x"38a4",x"3a69",x"309a",x"3a2f",x"3a57"),
(x"a172",x"3f5c",x"36eb",x"b3e5",x"3bb4",x"2ec2",x"3b20",x"3b17",x"a13d",x"3f5b",x"3716",x"a345",x"3bf7",x"2dcc",x"3b1a",x"3b17",x"a2d9",x"3f59",x"3714",x"b976",x"39c0",x"3024",x"3b1b",x"3b19"),
(x"a482",x"3f6f",x"36eb",x"bb61",x"b5a0",x"3119",x"3b30",x"3922",x"a425",x"3f70",x"370f",x"bbd3",x"af46",x"3182",x"3b2d",x"391f",x"a289",x"3f6b",x"370f",x"b891",x"ba72",x"30f5",x"3b2b",x"3921"),
(x"21ae",x"3fcd",x"36eb",x"3ade",x"37ab",x"31d3",x"3b41",x"38d7",x"20f7",x"3fcc",x"370e",x"3b7b",x"34a9",x"3270",x"3b3d",x"38d9",x"1aac",x"3fd4",x"3712",x"38b5",x"3a3e",x"32bd",x"3b3f",x"38df"),
(x"2496",x"3f5d",x"36eb",x"3bba",x"b376",x"2f14",x"3b35",x"3b31",x"2442",x"3f5d",x"3714",x"3b6b",x"b587",x"3095",x"3b30",x"3b31",x"24cc",x"3f69",x"3712",x"3bf0",x"aa00",x"2f46",x"3b31",x"3b38"),
(x"1fad",x"3f26",x"36eb",x"360d",x"3b5a",x"2ef4",x"3a31",x"3a5d",x"2409",x"3f24",x"36eb",x"3884",x"3a69",x"324a",x"3a33",x"3a59",x"2375",x"3f22",x"3711",x"38a4",x"3a69",x"309a",x"3a2f",x"3a57"),
(x"a38b",x"3f5a",x"36eb",x"bacc",x"3812",x"3065",x"3b20",x"3b19",x"a2d9",x"3f59",x"3714",x"b976",x"39c0",x"3024",x"3b1b",x"3b19",x"a38f",x"3f55",x"3712",x"bbe0",x"2e5e",x"30a3",x"3b1b",x"3b1b"),
(x"9f83",x"3f68",x"36eb",x"35e4",x"bb4d",x"31a2",x"3b2b",x"3927",x"a2ad",x"3f6a",x"36eb",x"b86e",x"ba87",x"313e",x"3b2e",x"3925",x"a289",x"3f6b",x"370f",x"b891",x"ba72",x"30f5",x"3b2b",x"3921"),
(x"980d",x"3fd7",x"36eb",x"b996",x"395e",x"33ec",x"3b44",x"38e0",x"1a0c",x"3fd7",x"36eb",x"38a6",x"3a54",x"3207",x"3b44",x"38de",x"1aac",x"3fd4",x"3712",x"38b5",x"3a3e",x"32bd",x"3b3f",x"38df"),
(x"250f",x"3f6a",x"36eb",x"3bef",x"2d0b",x"2e69",x"3b35",x"3b38",x"24cc",x"3f69",x"3712",x"3bf0",x"aa00",x"2f46",x"3b31",x"3b38",x"243c",x"3f75",x"3710",x"3b6a",x"35bb",x"2efe",x"3b31",x"3b3e"),
(x"1e52",x"3f28",x"36eb",x"3be6",x"308f",x"2c41",x"3a31",x"3a5e",x"1fad",x"3f26",x"36eb",x"360d",x"3b5a",x"2ef4",x"3a31",x"3a5d",x"1f0f",x"3f25",x"3718",x"38ae",x"3a78",x"2b7c",x"3a2c",x"3a5b"),
(x"a422",x"3f54",x"36eb",x"bbcf",x"b174",x"303e",x"3b1f",x"3b1c",x"a38f",x"3f55",x"3712",x"bbe0",x"2e5e",x"30a3",x"3b1b",x"3b1b",x"a2cb",x"3f51",x"3714",x"b972",x"b9bb",x"30de",x"3b1a",x"3b1d"),
(x"a2e9",x"3f24",x"3711",x"acd1",x"250b",x"3bf9",x"3bb9",x"3b9d",x"a0d2",x"3f23",x"3713",x"b0f4",x"19bc",x"3be7",x"3bb5",x"3b9f",x"a175",x"3f1a",x"3710",x"2828",x"260a",x"3bfe",x"3bb7",x"3ba6"),
(x"a175",x"3f1a",x"3710",x"2828",x"260a",x"3bfe",x"3bb7",x"3ba6",x"a2ee",x"3f13",x"3714",x"2eb0",x"28fa",x"3bf3",x"3bb9",x"3bab",x"a2e9",x"3f24",x"3711",x"acd1",x"250b",x"3bf9",x"3bb9",x"3b9d"),
(x"a1ea",x"3f0b",x"3712",x"a587",x"208e",x"3bff",x"3bb8",x"3bb2",x"a140",x"3f12",x"3714",x"2946",x"1ffc",x"3bfe",x"3bb7",x"3bac",x"a099",x"3f0e",x"3712",x"2953",x"27ae",x"3bfd",x"3bb6",x"3bb0"),
(x"a1ea",x"3f0b",x"3712",x"a587",x"208e",x"3bff",x"3bb8",x"3bb2",x"a2ee",x"3f13",x"3714",x"2eb0",x"28fa",x"3bf3",x"3bb9",x"3bab",x"a140",x"3f12",x"3714",x"2946",x"1ffc",x"3bfe",x"3bb7",x"3bac"),
(x"9d7f",x"3f04",x"3715",x"a0ea",x"2b00",x"3bfc",x"3bb3",x"3bb9",x"a1ea",x"3f0b",x"3712",x"a587",x"208e",x"3bff",x"3bb8",x"3bb2",x"9ecc",x"3f0b",x"3714",x"a8bf",x"2c22",x"3bfa",x"3bb4",x"3bb3"),
(x"17a2",x"3f01",x"3715",x"27e2",x"29b5",x"3bfc",x"3bae",x"3bbb",x"9d7f",x"3f04",x"3715",x"a0ea",x"2b00",x"3bfc",x"3bb3",x"3bb9",x"9aa8",x"3f08",x"3714",x"231d",x"2b5f",x"3bfc",x"3bb2",x"3bb5"),
(x"210b",x"3f04",x"3713",x"2b1d",x"aee4",x"3bf0",x"3ba7",x"3bb9",x"17a2",x"3f01",x"3715",x"27e2",x"29b5",x"3bfc",x"3bae",x"3bbb",x"1a1e",x"3f06",x"3715",x"270a",x"a779",x"3bfe",x"3bad",x"3bb7"),
(x"2466",x"3f0a",x"3715",x"a266",x"9d87",x"3bff",x"3ba1",x"3bb4",x"210b",x"3f04",x"3713",x"2b1d",x"aee4",x"3bf0",x"3ba7",x"3bb9",x"20b2",x"3f08",x"3716",x"24bc",x"aceb",x"3bf9",x"3ba8",x"3bb6"),
(x"253f",x"3f13",x"3715",x"a891",x"a7ce",x"3bfd",x"3b9e",x"3bad",x"2466",x"3f0a",x"3715",x"a266",x"9d87",x"3bff",x"3ba1",x"3bb4",x"2335",x"3f0e",x"3714",x"a8e0",x"299e",x"3bfc",x"3ba4",x"3bb1"),
(x"22d3",x"3f18",x"3715",x"ac67",x"28a5",x"3bf9",x"3ba4",x"3ba9",x"24fc",x"3f1b",x"3717",x"ad06",x"2793",x"3bf8",x"3b9f",x"3ba6",x"253f",x"3f13",x"3715",x"a891",x"a7ce",x"3bfd",x"3b9e",x"3bad"),
(x"2375",x"3f22",x"3711",x"a8d9",x"a52b",x"3bfe",x"3ba2",x"3ba0",x"24fc",x"3f1b",x"3717",x"ad06",x"2793",x"3bf8",x"3b9f",x"3ba6",x"22d3",x"3f18",x"3715",x"ac67",x"28a5",x"3bf9",x"3ba4",x"3ba9"),
(x"951c",x"3f19",x"3711",x"abef",x"a8a8",x"3bfa",x"3baf",x"3ba7",x"20d5",x"3f18",x"3714",x"aa45",x"2b10",x"3bfa",x"3ba7",x"3ba8",x"1e4f",x"3f16",x"3711",x"aa66",x"b31a",x"3bca",x"3baa",x"3baa"),
(x"1f0f",x"3f25",x"3718",x"ab65",x"b528",x"3b8f",x"3ba8",x"3b9d",x"3d81",x"3f23",x"3711",x"b40c",x"26bb",x"3bbc",x"3bae",x"3b9f",x"15a0",x"3f25",x"3713",x"b41f",x"ac3a",x"3bb6",x"3bad",x"3b9d"),
(x"16c6",x"3f29",x"3714",x"ade0",x"a4c2",x"3bf6",x"3bad",x"3b99",x"1d9c",x"3f28",x"3718",x"b420",x"1418",x"3bba",x"3ba9",x"3b9b",x"15a0",x"3f25",x"3713",x"b41f",x"ac3a",x"3bb6",x"3bad",x"3b9d"),
(x"16c6",x"3f29",x"3714",x"ade0",x"a4c2",x"3bf6",x"3bad",x"3b99",x"1d4f",x"3f31",x"3715",x"a7ae",x"a4ea",x"3bfe",x"3baa",x"3b93",x"1d9c",x"3f28",x"3718",x"b420",x"1418",x"3bba",x"3ba9",x"3b9b"),
(x"20d5",x"3f18",x"3714",x"aa45",x"2b10",x"3bfa",x"3ba7",x"3ba8",x"983c",x"3f20",x"3710",x"a856",x"a9ab",x"3bfc",x"3bb0",x"3ba1",x"2375",x"3f22",x"3711",x"a8d9",x"a52b",x"3bfe",x"3ba2",x"3ba0"),
(x"951c",x"3f19",x"3711",x"abef",x"a8a8",x"3bfa",x"3baf",x"3ba7",x"99ac",x"3f1c",x"3710",x"aa8d",x"2973",x"3bfb",x"3bb0",x"3ba5",x"983c",x"3f20",x"3710",x"a856",x"a9ab",x"3bfc",x"3bb0",x"3ba1"),
(x"a1bd",x"3ee0",x"3715",x"a1a1",x"23fc",x"3bff",x"3983",x"31eb",x"993e",x"3edf",x"3716",x"a82f",x"2808",x"3bfd",x"3988",x"31ea",x"a069",x"3ec3",x"3718",x"a24c",x"a379",x"3bff",x"3985",x"31ab"),
(x"16c6",x"3f29",x"3714",x"bbf3",x"ae23",x"2b27",x"3a63",x"3a30",x"15a0",x"3f25",x"3713",x"bbc2",x"33a4",x"298a",x"3a64",x"3a32",x"13e1",x"3f25",x"36eb",x"bbf6",x"2a70",x"2d61",x"3a69",x"3a31"),
(x"8dee",x"3f36",x"36eb",x"b469",x"bb91",x"316a",x"3a68",x"3a28",x"8dee",x"3f36",x"3718",x"b9e5",x"b968",x"0000",x"3a62",x"3a29",x"16c6",x"3f29",x"3714",x"bbf3",x"ae23",x"2b27",x"3a63",x"3a30"),
(x"1c89",x"3ddc",x"3716",x"b0f9",x"28af",x"3be5",x"3b6a",x"3b03",x"0f4a",x"3ddc",x"3712",x"b42b",x"ae69",x"3bae",x"3b66",x"3b03",x"9e24",x"3de5",x"370e",x"afd2",x"a717",x"3bef",x"3b62",x"3b0b"),
(x"2222",x"3de9",x"36eb",x"3b99",x"b315",x"330d",x"3b91",x"3a3c",x"1dd1",x"3dd9",x"36eb",x"3996",x"b95e",x"33ec",x"3b92",x"3a33",x"1c89",x"3ddc",x"3716",x"3add",x"b75a",x"334d",x"3b8c",x"3a34"),
(x"1ba5",x"3e29",x"3714",x"2c39",x"a9a5",x"3bf9",x"3b6e",x"3b46",x"2226",x"3e2b",x"3713",x"291b",x"ab55",x"3bfb",x"3b75",x"3b47",x"2079",x"3e21",x"3712",x"2a69",x"a87e",x"3bfc",x"3b72",x"3b3e"),
(x"2498",x"3e24",x"3711",x"2481",x"a546",x"3bff",x"3b7a",x"3b40",x"23f2",x"3e20",x"3712",x"aa38",x"2d35",x"3bf6",x"3b77",x"3b3d",x"21e0",x"3e1f",x"3711",x"2994",x"a977",x"3bfc",x"3b74",x"3b3d"),
(x"2079",x"3e21",x"3712",x"2a69",x"a87e",x"3bfc",x"3b72",x"3b3e",x"2226",x"3e2b",x"3713",x"291b",x"ab55",x"3bfb",x"3b75",x"3b47",x"242c",x"3e29",x"3712",x"2a73",x"aa97",x"3bfa",x"3b78",x"3b45"),
(x"2000",x"3e2e",x"3718",x"2e36",x"2160",x"3bf6",x"3b72",x"3b49",x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d",x"2360",x"3e2f",x"3711",x"2fec",x"2c2c",x"3beb",x"3b77",x"3b4a"),
(x"221a",x"3e47",x"3713",x"2e9c",x"b366",x"3bbd",x"3b76",x"3b5f",x"2437",x"3e45",x"370f",x"1df0",x"2631",x"3bff",x"3b7a",x"3b5d",x"2010",x"3e3f",x"370e",x"a6d5",x"a5c2",x"3bfe",x"3b73",x"3b59"),
(x"219e",x"3e3b",x"3713",x"2538",x"2c79",x"3bfa",x"3b75",x"3b54",x"2010",x"3e3f",x"370e",x"a6d5",x"a5c2",x"3bfe",x"3b73",x"3b59",x"2437",x"3e45",x"370f",x"1df0",x"2631",x"3bff",x"3b7a",x"3b5d"),
(x"24fa",x"3e37",x"370f",x"2ec5",x"9a24",x"3bf4",x"3b7c",x"3b51",x"21a8",x"3e39",x"3713",x"27ef",x"a84d",x"3bfd",x"3b75",x"3b53",x"219e",x"3e3b",x"3713",x"2538",x"2c79",x"3bfa",x"3b75",x"3b54"),
(x"21a8",x"3e39",x"3713",x"27ef",x"a84d",x"3bfd",x"3b75",x"3b53",x"24fa",x"3e37",x"370f",x"2ec5",x"9a24",x"3bf4",x"3b7c",x"3b51",x"2360",x"3e2f",x"3711",x"2fec",x"2c2c",x"3beb",x"3b77",x"3b4a"),
(x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d",x"1ce8",x"3e35",x"3713",x"a5bc",x"37de",x"3af6",x"3b70",x"3b50",x"2072",x"3e36",x"3710",x"2c5b",x"30a5",x"3be5",x"3b73",x"3b51"),
(x"2072",x"3e36",x"3710",x"2c5b",x"30a5",x"3be5",x"3b73",x"3b51",x"21a8",x"3e39",x"3713",x"27ef",x"a84d",x"3bfd",x"3b75",x"3b53",x"2360",x"3e2f",x"3711",x"2fec",x"2c2c",x"3beb",x"3b77",x"3b4a"),
(x"9959",x"3e66",x"3715",x"26c2",x"2c63",x"3bfa",x"3b6a",x"3b7a",x"1e50",x"3e66",x"3712",x"2f67",x"2981",x"3bf0",x"3b71",x"3b7a",x"125b",x"3e5e",x"3717",x"2ff2",x"2a7d",x"3bed",x"3b6c",x"3b73"),
(x"24ba",x"3e5b",x"3712",x"3163",x"2345",x"3be2",x"3b7b",x"3b71",x"245f",x"3e57",x"3714",x"2860",x"2f8b",x"3bf0",x"3b79",x"3b6d",x"2323",x"3e55",x"3716",x"2cd8",x"27e2",x"3bf9",x"3b77",x"3b6c"),
(x"2116",x"3e56",x"3716",x"a818",x"2d04",x"3bf8",x"3b74",x"3b6c",x"2074",x"3e62",x"3711",x"a40b",x"2d5c",x"3bf8",x"3b73",x"3b77",x"2458",x"3e5f",x"3714",x"9553",x"2b62",x"3bfc",x"3b79",x"3b74"),
(x"2074",x"3e62",x"3711",x"a40b",x"2d5c",x"3bf8",x"3b73",x"3b77",x"1e07",x"3e59",x"3714",x"2504",x"2da9",x"3bf7",x"3b70",x"3b6f",x"1acb",x"3e5c",x"3714",x"3036",x"273e",x"3bed",x"3b6e",x"3b72"),
(x"125b",x"3e5e",x"3717",x"2ff2",x"2a7d",x"3bed",x"3b6c",x"3b73",x"1e50",x"3e66",x"3712",x"2f67",x"2981",x"3bf0",x"3b71",x"3b7a",x"1f03",x"3e64",x"3711",x"327d",x"975f",x"3bd5",x"3b71",x"3b78"),
(x"1f03",x"3e64",x"3711",x"327d",x"975f",x"3bd5",x"3b71",x"3b78",x"2074",x"3e62",x"3711",x"a40b",x"2d5c",x"3bf8",x"3b73",x"3b77",x"1acb",x"3e5c",x"3714",x"3036",x"273e",x"3bed",x"3b6e",x"3b72"),
(x"1f3f",x"3e6b",x"3712",x"3146",x"ac91",x"3bde",x"3b71",x"3b7e",x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c"),
(x"9aa8",x"3e77",x"3718",x"a138",x"2e95",x"3bf4",x"3b69",x"3b89",x"9fe7",x"3e77",x"3719",x"23bb",x"a7ae",x"3bfe",x"3b66",x"3b89",x"9ff6",x"3e78",x"3719",x"290e",x"2f00",x"3bf2",x"3b66",x"3b89"),
(x"9920",x"3e76",x"3718",x"ab4f",x"a525",x"3bfc",x"3b6a",x"3b88",x"9aa8",x"3e77",x"3718",x"a138",x"2e95",x"3bf4",x"3b69",x"3b89",x"1c29",x"3e7b",x"3718",x"2e3b",x"9fae",x"3bf6",x"3b6f",x"3b8c"),
(x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"9dca",x"3e73",x"3715",x"ad65",x"2c5a",x"3bf3",x"3b67",x"3b85",x"9920",x"3e76",x"3718",x"ab4f",x"a525",x"3bfc",x"3b6a",x"3b88"),
(x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"9d58",x"3e68",x"3717",x"ad2d",x"aecb",x"3bed",x"3b67",x"3b7c",x"a0a3",x"3e6e",x"3718",x"acf2",x"991e",x"3bf9",x"3b64",x"3b81"),
(x"a0f6",x"3e69",x"3712",x"b59c",x"b36a",x"3b42",x"3b64",x"3b7d",x"a0a3",x"3e6e",x"3718",x"acf2",x"991e",x"3bf9",x"3b64",x"3b81",x"9d58",x"3e68",x"3717",x"ad2d",x"aecb",x"3bed",x"3b67",x"3b7c"),
(x"3b57",x"3e6e",x"3718",x"2bb4",x"a8d3",x"3bfa",x"3b6c",x"3b81",x"1f3f",x"3e6b",x"3712",x"3146",x"ac91",x"3bde",x"3b71",x"3b7e",x"9b02",x"3e67",x"3716",x"3009",x"ada6",x"3be7",x"3b69",x"3b7b"),
(x"9b02",x"3e67",x"3716",x"3009",x"ada6",x"3be7",x"3b69",x"3b7b",x"1f3f",x"3e6b",x"3712",x"3146",x"ac91",x"3bde",x"3b71",x"3b7e",x"1e50",x"3e66",x"3712",x"2f67",x"2981",x"3bf0",x"3b71",x"3b7a"),
(x"9607",x"3e5d",x"3717",x"17c8",x"1f79",x"3c00",x"3b6a",x"3b72",x"9ec5",x"3e5f",x"3718",x"2c00",x"a90e",x"3bfa",x"3b66",x"3b75",x"9abe",x"3e63",x"3714",x"257a",x"2e8a",x"3bf4",x"3b69",x"3b78"),
(x"9607",x"3e5d",x"3717",x"17c8",x"1f79",x"3c00",x"3b6a",x"3b72",x"9e13",x"3e58",x"3715",x"251e",x"ad06",x"3bf9",x"3b67",x"3b6e",x"9ec5",x"3e5f",x"3718",x"2c00",x"a90e",x"3bfa",x"3b66",x"3b75"),
(x"9e13",x"3e58",x"3715",x"251e",x"ad06",x"3bf9",x"3b67",x"3b6e",x"a123",x"3e50",x"3714",x"adba",x"a266",x"3bf7",x"3b63",x"3b68",x"a29f",x"3e53",x"3714",x"975f",x"ac2c",x"3bfb",x"3b61",x"3b6a"),
(x"a123",x"3e50",x"3714",x"adba",x"a266",x"3bf7",x"3b63",x"3b68",x"a180",x"3e45",x"3715",x"b468",x"a47a",x"3bb0",x"3b63",x"3b5e",x"a3b3",x"3e47",x"3712",x"b106",x"a73e",x"3be5",x"3b5f",x"3b60"),
(x"a180",x"3e45",x"3715",x"b468",x"a47a",x"3bb0",x"3b63",x"3b5e",x"a0d7",x"3e3d",x"3717",x"b273",x"af43",x"3bc8",x"3b64",x"3b57",x"a294",x"3e3b",x"3710",x"b550",x"ae33",x"3b81",x"3b61",x"3b55"),
(x"a0d7",x"3e3d",x"3717",x"b273",x"af43",x"3bc8",x"3b64",x"3b57",x"9ad5",x"3e36",x"3711",x"2e24",x"aa2b",x"3bf4",x"3b69",x"3b51",x"9faa",x"3e33",x"3712",x"ab5c",x"a345",x"3bfc",x"3b65",x"3b4f"),
(x"11f0",x"3e35",x"3712",x"add2",x"304b",x"3be4",x"3b6c",x"3b50",x"1b46",x"3e2e",x"3716",x"af4b",x"2a5f",x"3bf0",x"3b6e",x"3b49",x"9faa",x"3e33",x"3712",x"ab5c",x"a345",x"3bfc",x"3b65",x"3b4f"),
(x"11f0",x"3e35",x"3712",x"add2",x"304b",x"3be4",x"3b6c",x"3b50",x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d",x"1b46",x"3e2e",x"3716",x"af4b",x"2a5f",x"3bf0",x"3b6e",x"3b49"),
(x"11f0",x"3e35",x"3712",x"add2",x"304b",x"3be4",x"3b6c",x"3b50",x"1ce8",x"3e35",x"3713",x"a5bc",x"37de",x"3af6",x"3b70",x"3b50",x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d"),
(x"1b46",x"3e2e",x"3716",x"af4b",x"2a5f",x"3bf0",x"3b6e",x"3b49",x"1c86",x"3e32",x"3718",x"2c13",x"31c5",x"3bda",x"3b6f",x"3b4d",x"2000",x"3e2e",x"3718",x"2e36",x"2160",x"3bf6",x"3b72",x"3b49"),
(x"212c",x"3e2d",x"3716",x"2f15",x"b29c",x"3bc6",x"3b73",x"3b48",x"1ba5",x"3e29",x"3714",x"2c39",x"a9a5",x"3bf9",x"3b6e",x"3b46",x"1d2c",x"3e2c",x"3716",x"2553",x"b2c7",x"3bd1",x"3b6f",x"3b48"),
(x"212c",x"3e2d",x"3716",x"2f15",x"b29c",x"3bc6",x"3b73",x"3b48",x"2226",x"3e2b",x"3713",x"291b",x"ab55",x"3bfb",x"3b75",x"3b47",x"1ba5",x"3e29",x"3714",x"2c39",x"a9a5",x"3bf9",x"3b6e",x"3b46"),
(x"1f0d",x"3e22",x"3713",x"2da3",x"af14",x"3beb",x"3b70",x"3b3f",x"16e7",x"3e1d",x"370f",x"2edc",x"acd0",x"3bee",x"3b6c",x"3b3b",x"9aec",x"3e22",x"3717",x"30e7",x"b057",x"3bd4",x"3b68",x"3b3f"),
(x"16e7",x"3e1d",x"370f",x"2edc",x"acd0",x"3bee",x"3b6c",x"3b3b",x"9631",x"3e13",x"3716",x"2adf",x"26b5",x"3bfc",x"3b69",x"3b32",x"a039",x"3e14",x"3713",x"29b8",x"26e9",x"3bfd",x"3b64",x"3b34"),
(x"a12d",x"3df8",x"370d",x"b809",x"ae09",x"3add",x"3b5f",x"3b1c",x"a1a0",x"3dfc",x"370f",x"b6ca",x"afac",x"3b2e",x"3b5f",x"3b1f",x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a"),
(x"9f80",x"3def",x"3712",x"a9f0",x"ab1d",x"3bfa",x"3b61",x"3b14",x"2043",x"3df7",x"3715",x"99bc",x"26cf",x"3bff",x"3b6f",x"3b19",x"20de",x"3dea",x"3715",x"ad56",x"a0d0",x"3bf8",x"3b6f",x"3b0e"),
(x"1624",x"3e08",x"370e",x"3b5f",x"35f1",x"2f4d",x"3b89",x"3a4c",x"17f3",x"3e09",x"36eb",x"3b4a",x"3677",x"2cf9",x"3b8e",x"3a4d",x"2166",x"3df7",x"36eb",x"3b89",x"3473",x"31fc",x"3b90",x"3a43"),
(x"235a",x"3e97",x"3710",x"bbfd",x"2997",x"a0a8",x"3b38",x"3b56",x"22b8",x"3e8e",x"3713",x"bba5",x"3497",x"ac28",x"3b38",x"3b5a",x"2307",x"3e8d",x"36eb",x"bba1",x"34cc",x"1f45",x"3b3d",x"3b5a"),
(x"234d",x"3e9c",x"36eb",x"bbf5",x"ae59",x"2467",x"3b3d",x"3b53",x"2325",x"3e9e",x"3714",x"bbeb",x"b08a",x"98b5",x"3b38",x"3b52",x"235a",x"3e97",x"3710",x"bbfd",x"2997",x"a0a8",x"3b38",x"3b56"),
(x"2002",x"3e80",x"3714",x"bb1c",x"3754",x"223f",x"3b37",x"3b62",x"1c29",x"3e7b",x"3718",x"39e5",x"3968",x"0000",x"3b37",x"3b65",x"1c29",x"3e7b",x"36eb",x"346a",x"3b91",x"316a",x"3b3c",x"3b66"),
(x"2307",x"3e8d",x"36eb",x"bba1",x"34cc",x"1f45",x"3b3d",x"3b5a",x"22b8",x"3e8e",x"3713",x"bba5",x"3497",x"ac28",x"3b38",x"3b5a",x"2002",x"3e80",x"3714",x"bb1c",x"3754",x"223f",x"3b37",x"3b62"),
(x"227e",x"3ea3",x"3712",x"bb76",x"b5c5",x"204d",x"3b38",x"3b4f",x"2325",x"3e9e",x"3714",x"bbeb",x"b08a",x"98b5",x"3b38",x"3b52",x"234d",x"3e9c",x"36eb",x"bbf5",x"ae59",x"2467",x"3b3d",x"3b53"),
(x"2237",x"3ea4",x"36eb",x"bab1",x"b862",x"21f0",x"3b3d",x"3b4f",x"214b",x"3ea6",x"3714",x"b95a",x"b9f1",x"2025",x"3b38",x"3b4d",x"227e",x"3ea3",x"3712",x"bb76",x"b5c5",x"204d",x"3b38",x"3b4f"),
(x"1f6a",x"3ea8",x"36eb",x"b7e1",x"baf5",x"269a",x"3b3d",x"3b4b",x"1f1f",x"3ea8",x"3714",x"b5bf",x"bb76",x"27db",x"3b38",x"3b4b",x"214b",x"3ea6",x"3714",x"b95a",x"b9f1",x"2025",x"3b38",x"3b4d"),
(x"142d",x"3eaa",x"36eb",x"b03c",x"bbeb",x"299b",x"3b3d",x"3b48",x"11db",x"3eaa",x"3715",x"2836",x"bbfd",x"294f",x"3b38",x"3b47",x"1f1f",x"3ea8",x"3714",x"b5bf",x"bb76",x"27db",x"3b38",x"3b4b"),
(x"9d76",x"3ea9",x"36eb",x"3868",x"baab",x"296a",x"3b3d",x"3b44",x"9d99",x"3ea9",x"3716",x"386f",x"baa7",x"2604",x"3b38",x"3b44",x"11db",x"3eaa",x"3715",x"2836",x"bbfd",x"294f",x"3b38",x"3b47"),
(x"9d76",x"3ea9",x"36eb",x"3868",x"baab",x"296a",x"3b3d",x"3b44",x"a11a",x"3ea2",x"36eb",x"3af3",x"b7df",x"2b38",x"3b3e",x"3b40",x"a14f",x"3ea3",x"3714",x"3b01",x"b7b5",x"2839",x"3b39",x"3b40"),
(x"a1ea",x"3e9d",x"36eb",x"3bf9",x"ad11",x"2511",x"3b3e",x"3b3d",x"a1ee",x"3e9d",x"3714",x"3be6",x"310f",x"9bfc",x"3b39",x"3b3d",x"a14f",x"3ea3",x"3714",x"3b01",x"b7b5",x"2839",x"3b39",x"3b40"),
(x"a11a",x"3e99",x"36eb",x"390c",x"3a34",x"2532",x"3b3e",x"3b3b",x"a0ed",x"3e98",x"3715",x"3928",x"3a1d",x"1553",x"3b39",x"3b3a",x"a1ee",x"3e9d",x"3714",x"3be6",x"310f",x"9bfc",x"3b39",x"3b3d"),
(x"a11a",x"3e99",x"36eb",x"390c",x"3a34",x"2532",x"3b3e",x"3b3b",x"9d99",x"3e98",x"36eb",x"b5dd",x"3b6d",x"2be9",x"3b3e",x"3b38",x"9ddf",x"3e98",x"3714",x"afe4",x"3bee",x"28fd",x"3b39",x"3b38"),
(x"9d99",x"3e98",x"36eb",x"b5dd",x"3b6d",x"2be9",x"3b3e",x"3b38",x"99c6",x"3e9b",x"36eb",x"b2b1",x"3bc8",x"2e54",x"3b3f",x"3b37",x"9908",x"3e9a",x"3711",x"b64f",x"3b52",x"2d1b",x"3b3a",x"3b36"),
(x"199d",x"3e8c",x"36eb",x"3bf6",x"aa70",x"2d61",x"3b3e",x"3b29",x"18c5",x"3e8c",x"3713",x"3bc2",x"b3a4",x"298a",x"3b39",x"3b2a",x"1b8a",x"3e8e",x"3711",x"3a7a",x"b8af",x"2839",x"3b39",x"3b2c"),
(x"99c6",x"3e9b",x"36eb",x"b2b1",x"3bc8",x"2e54",x"3b3f",x"3b37",x"1ab2",x"3e9b",x"36eb",x"337e",x"3bba",x"2ef6",x"3b3f",x"3b33",x"1937",x"3e9a",x"3710",x"3416",x"3bad",x"2f8d",x"3b3a",x"3b33"),
(x"21a6",x"3e48",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b1f",x"3b51",x"221a",x"3e47",x"3713",x"b583",x"3b63",x"3153",x"3b1a",x"3b4f",x"1fdf",x"3e42",x"370f",x"ba9b",x"3854",x"30fa",x"3b19",x"3b52"),
(x"2166",x"3df7",x"36eb",x"3b89",x"3473",x"31fc",x"3b90",x"3a43",x"2222",x"3de9",x"36eb",x"3b99",x"b315",x"330d",x"3b91",x"3a3c",x"20de",x"3dea",x"3715",x"3bc5",x"ab9a",x"3358",x"3b8c",x"3a3c"),
(x"1de8",x"3e90",x"3710",x"2856",x"29ab",x"3bfc",x"3b71",x"3b9e",x"1b8a",x"3e8e",x"3711",x"340c",x"a6c2",x"3bbc",x"3b6f",x"3b9c",x"9a89",x"3e8b",x"3718",x"2b65",x"3528",x"3b8f",x"3b69",x"3b9a"),
(x"9e52",x"3df5",x"36eb",x"bbe3",x"ace8",x"30c3",x"3b8a",x"3a22",x"9f80",x"3def",x"3712",x"bbcf",x"3082",x"3141",x"3b88",x"3a28",x"a0ba",x"3def",x"36eb",x"bbdb",x"9c67",x"320a",x"3b8c",x"3a25"),
(x"9e52",x"3df5",x"36eb",x"bbe3",x"ace8",x"30c3",x"3b8a",x"3a22",x"9de0",x"3df4",x"3715",x"bbd7",x"31f9",x"2c2a",x"3b86",x"3a26",x"9f80",x"3def",x"3712",x"bbcf",x"3082",x"3141",x"3b88",x"3a28"),
(x"a081",x"3e33",x"36eb",x"b958",x"b9de",x"2fdf",x"3a3f",x"3a41",x"a2ed",x"3e3a",x"36eb",x"bb75",x"b5a2",x"2d46",x"3a3f",x"3a3c",x"a294",x"3e3b",x"3710",x"bb6a",x"b5bb",x"2efe",x"3a3b",x"3a3c"),
(x"1e0f",x"3e99",x"36eb",x"3aa4",x"3859",x"2fe4",x"3b3f",x"3b31",x"1d11",x"3e98",x"3711",x"3a7e",x"3887",x"3089",x"3b3a",x"3b31",x"1937",x"3e9a",x"3710",x"3416",x"3bad",x"2f8d",x"3b3a",x"3b33"),
(x"990f",x"3e89",x"36eb",x"bbe6",x"b08f",x"2c41",x"3b3a",x"38ac",x"9747",x"3e88",x"3718",x"bbe6",x"b09f",x"2baa",x"3b35",x"38aa",x"9613",x"3e7f",x"3715",x"bbfa",x"2710",x"2c48",x"3b33",x"38ae"),
(x"1e0f",x"3e99",x"36eb",x"3aa4",x"3859",x"2fe4",x"3b3f",x"3b31",x"1f98",x"3e94",x"36eb",x"3bf4",x"1edc",x"2ebb",x"3b3f",x"3b2f",x"1ea1",x"3e94",x"3710",x"3bcc",x"3228",x"2f2f",x"3b3a",x"3b30"),
(x"1e92",x"3e42",x"36eb",x"bb7d",x"3521",x"3096",x"3b1d",x"3b54",x"1fdf",x"3e42",x"370f",x"ba9b",x"3854",x"30fa",x"3b19",x"3b52",x"2010",x"3e3f",x"370e",x"bb25",x"b70d",x"2d6a",x"3b19",x"3b53"),
(x"247a",x"3e61",x"36eb",x"36fe",x"3b25",x"2ea4",x"3b42",x"385c",x"2458",x"3e5f",x"3714",x"3972",x"39bb",x"30de",x"3b3d",x"385c",x"2074",x"3e62",x"3711",x"34dc",x"3b97",x"2d61",x"3b3e",x"3861"),
(x"1bc8",x"3e8d",x"36eb",x"39db",x"b96c",x"2c1a",x"3b3e",x"3b2b",x"1b8a",x"3e8e",x"3711",x"3a7a",x"b8af",x"2839",x"3b39",x"3b2c",x"1de8",x"3e90",x"3710",x"3b2f",x"b6d9",x"2e52",x"3b3a",x"3b2d"),
(x"1c1b",x"3e2d",x"36eb",x"b776",x"bb0b",x"2d41",x"3a3f",x"3a49",x"a081",x"3e33",x"36eb",x"b958",x"b9de",x"2fdf",x"3a3f",x"3a41",x"9faa",x"3e33",x"3712",x"b84e",x"bab0",x"2ec8",x"3a3a",x"3a41"),
(x"9943",x"3e7e",x"36eb",x"b9df",x"3964",x"2d28",x"3b37",x"38b2",x"989a",x"3e7f",x"36eb",x"bbfa",x"20b5",x"2cb4",x"3b37",x"38b1",x"9613",x"3e7f",x"3715",x"bbfa",x"2710",x"2c48",x"3b33",x"38ae"),
(x"2166",x"3e3a",x"36eb",x"bad3",x"b822",x"2c4d",x"3b1b",x"3b58",x"1f2f",x"3e3f",x"36eb",x"bb19",x"b744",x"2cf7",x"3b1c",x"3b55",x"2010",x"3e3f",x"370e",x"bb25",x"b70d",x"2d6a",x"3b19",x"3b53"),
(x"95be",x"3e13",x"36eb",x"3bfe",x"9ea7",x"2828",x"3b8c",x"3a53",x"17f3",x"3e09",x"36eb",x"3b4a",x"3677",x"2cf9",x"3b8e",x"3a4d",x"1624",x"3e08",x"370e",x"3b5f",x"35f1",x"2f4d",x"3b89",x"3a4c"),
(x"1c1b",x"3e2d",x"36eb",x"b776",x"bb0b",x"2d41",x"3a3f",x"3a49",x"1b46",x"3e2e",x"3716",x"b7e9",x"baf1",x"2aa7",x"3a3a",x"3a48",x"1d2c",x"3e2c",x"3716",x"bbde",x"b1b6",x"2825",x"3a3a",x"3a49"),
(x"a0ef",x"3e78",x"36eb",x"b9ed",x"394b",x"2f45",x"3b35",x"38b6",x"9943",x"3e7e",x"36eb",x"b9df",x"3964",x"2d28",x"3b37",x"38b2",x"98e9",x"3e7d",x"3715",x"b95d",x"39e3",x"2de3",x"3b32",x"38af"),
(x"1f03",x"3e64",x"3711",x"3b12",x"3763",x"2ca3",x"3b3e",x"3862",x"1e50",x"3e66",x"3712",x"3bf7",x"a83f",x"2d8f",x"3b3e",x"3863",x"1f30",x"3e66",x"36eb",x"3bf8",x"2379",x"2d44",x"3b43",x"3863"),
(x"201d",x"3e63",x"36eb",x"37d8",x"3af6",x"2a35",x"3b42",x"3861",x"2074",x"3e62",x"3711",x"34dc",x"3b97",x"2d61",x"3b3e",x"3861",x"1f03",x"3e64",x"3711",x"3b12",x"3763",x"2ca3",x"3b3e",x"3862"),
(x"216e",x"3e39",x"36eb",x"b9e9",x"3955",x"2e31",x"3b34",x"382e",x"2166",x"3e3a",x"36eb",x"bad3",x"b822",x"2c4d",x"3b33",x"382d",x"219e",x"3e3b",x"3713",x"bb5b",x"b634",x"2c03",x"3b2f",x"382e"),
(x"95be",x"3e13",x"36eb",x"3bfe",x"9ea7",x"2828",x"3b8c",x"3a53",x"9631",x"3e13",x"3716",x"3bff",x"a0c2",x"2138",x"3b87",x"3a51",x"16e7",x"3e1d",x"370f",x"3ad7",x"b821",x"29e6",x"3b87",x"3a57"),
(x"1cd4",x"3e2c",x"36eb",x"bb24",x"371c",x"2cde",x"3a3f",x"3a49",x"1d2c",x"3e2c",x"3716",x"bbde",x"b1b6",x"2825",x"3a3a",x"3a49",x"1ba5",x"3e29",x"3714",x"b9e8",x"3951",x"2f27",x"3a3a",x"3a4a"),
(x"a0ef",x"3e78",x"36eb",x"b9ed",x"394b",x"2f45",x"3b35",x"38b6",x"9ff6",x"3e78",x"3719",x"b9a6",x"3994",x"2fc6",x"3b30",x"38b3",x"9fe7",x"3e77",x"3719",x"b250",x"bbca",x"2f22",x"3b30",x"38b3"),
(x"1f30",x"3e66",x"36eb",x"3bf8",x"2379",x"2d44",x"3b43",x"3863",x"1e50",x"3e66",x"3712",x"3bf7",x"a83f",x"2d8f",x"3b3e",x"3863",x"1f3f",x"3e6b",x"3712",x"3b92",x"b509",x"2cb0",x"3b3e",x"3866"),
(x"2072",x"3e36",x"3710",x"b833",x"3ac7",x"2d1d",x"3b2f",x"3831",x"1ce8",x"3e35",x"3713",x"b0a8",x"3bea",x"22dc",x"3b30",x"3833",x"1c5d",x"3e35",x"36eb",x"b046",x"3be8",x"2cb7",x"3b34",x"3832"),
(x"216e",x"3e39",x"36eb",x"b9e9",x"3955",x"2e31",x"3b34",x"382e",x"21a8",x"3e39",x"3713",x"bb09",x"3791",x"2ab8",x"3b2f",x"382f",x"2072",x"3e36",x"3710",x"b833",x"3ac7",x"2d1d",x"3b2f",x"3831"),
(x"1fba",x"3e21",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b8a",x"3a5c",x"17ea",x"3e1d",x"36eb",x"3ab4",x"b859",x"2a66",x"3b8b",x"3a58",x"16e7",x"3e1d",x"370f",x"3ad7",x"b821",x"29e6",x"3b87",x"3a57"),
(x"1986",x"3e2a",x"36eb",x"b97a",x"39b6",x"309a",x"3a3f",x"3a4b",x"1ba5",x"3e29",x"3714",x"b9e8",x"3951",x"2f27",x"3a3a",x"3a4a",x"9aec",x"3e22",x"3717",x"ba77",x"3889",x"310e",x"3a3a",x"3a50"),
(x"9950",x"3e76",x"36eb",x"bb01",x"b745",x"3141",x"3b32",x"38b9",x"a09e",x"3e76",x"36eb",x"b2cb",x"bbc1",x"2fc5",x"3b35",x"38b7",x"9fe7",x"3e77",x"3719",x"b250",x"bbca",x"2f22",x"3b30",x"38b3"),
(x"1fbf",x"3e6a",x"36eb",x"3b57",x"b625",x"2e99",x"3b43",x"3865",x"1f3f",x"3e6b",x"3712",x"3b92",x"b509",x"2cb0",x"3b3e",x"3866",x"2353",x"3e7c",x"3711",x"3b70",x"b585",x"3014",x"3b3f",x"3870"),
(x"11f0",x"3e35",x"3712",x"32e8",x"3bcb",x"2c10",x"3b30",x"3835",x"9ad5",x"3e36",x"3711",x"3934",x"3a0d",x"2c18",x"3b31",x"3837",x"9a03",x"3e37",x"36eb",x"374a",x"3b15",x"2de4",x"3b35",x"3836"),
(x"1c5d",x"3e35",x"36eb",x"b046",x"3be8",x"2cb7",x"3b34",x"3832",x"1ce8",x"3e35",x"3713",x"b0a8",x"3bea",x"22dc",x"3b30",x"3833",x"11f0",x"3e35",x"3712",x"32e8",x"3bcb",x"2c10",x"3b30",x"3835"),
(x"1fba",x"3e21",x"36eb",x"373f",x"bb1a",x"2d3c",x"3b1b",x"3b2d",x"1f0d",x"3e22",x"3713",x"37c3",x"baf3",x"2e28",x"3b17",x"3b30",x"2079",x"3e21",x"3712",x"b721",x"bb24",x"2bf9",x"3b17",x"3b30"),
(x"9d26",x"3e23",x"36eb",x"baff",x"373c",x"3197",x"3a3f",x"3a50",x"9aec",x"3e22",x"3717",x"ba77",x"3889",x"310e",x"3a3a",x"3a50",x"a039",x"3e14",x"3713",x"bbc6",x"31be",x"30de",x"3a3a",x"3a57"),
(x"2422",x"3e7d",x"36eb",x"3b99",x"b45f",x"30d6",x"3b44",x"3870",x"2353",x"3e7c",x"3711",x"3b70",x"b585",x"3014",x"3b3f",x"3870",x"2467",x"3e8c",x"3711",x"3be4",x"ad1e",x"308c",x"3b40",x"3878"),
(x"a09f",x"3e3d",x"36eb",x"3aaf",x"3860",x"2a70",x"3b37",x"383a",x"9a03",x"3e37",x"36eb",x"374a",x"3b15",x"2de4",x"3b35",x"3836",x"9ad5",x"3e36",x"3711",x"3934",x"3a0d",x"2c18",x"3b31",x"3837"),
(x"20b1",x"3e20",x"36eb",x"b8ae",x"ba73",x"2d47",x"3b1b",x"3b2e",x"2079",x"3e21",x"3712",x"b721",x"bb24",x"2bf9",x"3b17",x"3b30",x"21e0",x"3e1f",x"3711",x"b5dd",x"bb65",x"2eae",x"3b18",x"3b32"),
(x"a0d9",x"3e07",x"36eb",x"bbea",x"2e09",x"2f12",x"3a3e",x"3a5f",x"a139",x"3e14",x"36eb",x"bbbf",x"3113",x"322d",x"3a3f",x"3a58",x"a039",x"3e14",x"3713",x"bbc6",x"31be",x"30de",x"3a3a",x"3a57"),
(x"9950",x"3e76",x"36eb",x"bb01",x"b745",x"3141",x"3b82",x"396a",x"9dca",x"3e73",x"3715",x"b9d1",x"3974",x"2cc6",x"3b84",x"396f",x"9fd8",x"3e72",x"36eb",x"ba0e",x"3929",x"2e76",x"3b85",x"396a"),
(x"9950",x"3e76",x"36eb",x"bb01",x"b745",x"3141",x"3b82",x"396a",x"9920",x"3e76",x"3718",x"baf6",x"37e1",x"2460",x"3b82",x"3970",x"9dca",x"3e73",x"3715",x"b9d1",x"3974",x"2cc6",x"3b84",x"396f"),
(x"24b3",x"3e9d",x"36eb",x"3be8",x"2d66",x"3010",x"3b45",x"3881",x"24be",x"3e8c",x"36eb",x"3be6",x"ac77",x"308c",x"3b44",x"3878",x"2467",x"3e8c",x"3711",x"3be4",x"ad1e",x"308c",x"3b40",x"3878"),
(x"a166",x"3e45",x"36eb",x"3bfa",x"2c62",x"2617",x"3b38",x"383e",x"a09f",x"3e3d",x"36eb",x"3aaf",x"3860",x"2a70",x"3b37",x"383a",x"a0d7",x"3e3d",x"3717",x"3b6f",x"35e5",x"261e",x"3b32",x"383c"),
(x"21ab",x"3e1e",x"36eb",x"ae29",x"bbe6",x"3005",x"3b1c",x"3b2f",x"21e0",x"3e1f",x"3711",x"b5dd",x"bb65",x"2eae",x"3b18",x"3b32",x"23f2",x"3e20",x"3712",x"35a5",x"bb63",x"30cc",x"3b19",x"3b34"),
(x"a0d9",x"3e07",x"36eb",x"bbea",x"2e09",x"2f12",x"3a3e",x"3a5f",x"a08e",x"3e07",x"3717",x"bbf0",x"2f10",x"2aec",x"3a39",x"3a5e",x"a1a0",x"3dfc",x"370f",x"bbdd",x"30de",x"2e6c",x"3a39",x"3a64"),
(x"9fd8",x"3e72",x"36eb",x"ba0e",x"3929",x"2e76",x"3b85",x"396a",x"9dca",x"3e73",x"3715",x"b9d1",x"3974",x"2cc6",x"3b84",x"396f",x"a0a3",x"3e6e",x"3718",x"bb13",x"3732",x"2fec",x"3b87",x"396f"),
(x"24b3",x"3e9d",x"36eb",x"3be8",x"2d66",x"3010",x"3b45",x"3881",x"2469",x"3e9d",x"3714",x"3bec",x"2d02",x"2f48",x"3b40",x"3881",x"23cf",x"3ea5",x"3712",x"3b45",x"3640",x"30a6",x"3b40",x"3885"),
(x"1f98",x"3e94",x"36eb",x"3bf4",x"1edc",x"2ebb",x"3b3f",x"3b2f",x"1edf",x"3e90",x"36eb",x"3b02",x"b776",x"2fc8",x"3b3e",x"3b2c",x"1de8",x"3e90",x"3710",x"3b2f",x"b6d9",x"2e52",x"3b3a",x"3b2d"),
(x"a0d8",x"3e4f",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"3b3a",x"3843",x"a166",x"3e45",x"36eb",x"3bfa",x"2c62",x"2617",x"3b38",x"383e",x"a180",x"3e45",x"3715",x"3bfe",x"a412",x"2867",x"3b33",x"3840"),
(x"244f",x"3e1f",x"36eb",x"3913",x"ba0d",x"310f",x"3b1e",x"3b32",x"23f2",x"3e20",x"3712",x"35a5",x"bb63",x"30cc",x"3b19",x"3b34",x"2498",x"3e24",x"3711",x"3bb2",x"b32f",x"30f4",x"3b1a",x"3b36"),
(x"a243",x"3dfc",x"36eb",x"bbe4",x"2adf",x"30ee",x"3a3d",x"3a65",x"a1a0",x"3dfc",x"370f",x"bbdd",x"30de",x"2e6c",x"3a39",x"3a64",x"a12d",x"3df8",x"370d",x"bb0d",x"b70c",x"3169",x"3a39",x"3a66"),
(x"a164",x"3e6e",x"36eb",x"bbbf",x"3333",x"2ed0",x"3b87",x"3969",x"a0a3",x"3e6e",x"3718",x"bb13",x"3732",x"2fec",x"3b87",x"396f",x"a0f6",x"3e69",x"3712",x"bbf0",x"ac20",x"2e95",x"3b8a",x"396e"),
(x"2427",x"3ea6",x"36eb",x"3ab2",x"3834",x"30cb",x"3b45",x"3886",x"23cf",x"3ea5",x"3712",x"3b45",x"3640",x"30a6",x"3b40",x"3885",x"20a5",x"3eac",x"3715",x"393c",x"39e9",x"3110",x"3b40",x"388b"),
(x"9d2f",x"3e57",x"36eb",x"3ac2",x"b833",x"2e8a",x"3b3b",x"3848",x"a0d8",x"3e4f",x"36eb",x"3bcf",x"b2aa",x"2bc5",x"3b3a",x"3843",x"a123",x"3e50",x"3714",x"3b81",x"b558",x"2da5",x"3b35",x"3845"),
(x"24ee",x"3e23",x"36eb",x"3be5",x"2dbc",x"3036",x"3b1f",x"3b34",x"2498",x"3e24",x"3711",x"3bb2",x"b32f",x"30f4",x"3b1a",x"3b36",x"242c",x"3e29",x"3712",x"3ae4",x"37c3",x"30c9",x"3b1b",x"3b39"),
(x"a088",x"3df5",x"36eb",x"b571",x"bb6d",x"30cc",x"3a3d",x"3a69",x"a1da",x"3df6",x"36eb",x"baf6",x"b714",x"32f0",x"3a3d",x"3a68",x"a12d",x"3df8",x"370d",x"bb0d",x"b70c",x"3169",x"3a39",x"3a66"),
(x"a13e",x"3e68",x"36eb",x"bbbf",x"b370",x"2dad",x"3b8a",x"3969",x"a0f6",x"3e69",x"3712",x"bbf0",x"ac20",x"2e95",x"3b8a",x"396e",x"a072",x"3e68",x"3712",x"b297",x"bbcc",x"2d84",x"3b8b",x"396f"),
(x"20e4",x"3eae",x"36eb",x"37cb",x"3ae6",x"3068",x"3b45",x"388b",x"20a5",x"3eac",x"3715",x"393c",x"39e9",x"3110",x"3b40",x"388b",x"1788",x"3eaf",x"3715",x"1ef6",x"3bee",x"302a",x"3b3f",x"388f"),
(x"9470",x"3e5c",x"36eb",x"39cd",x"b979",x"2caa",x"3b3c",x"384b",x"9d2f",x"3e57",x"36eb",x"3ac2",x"b833",x"2e8a",x"3b3b",x"3848",x"9e13",x"3e58",x"3715",x"3a65",x"b8c1",x"2d9c",x"3b36",x"384a"),
(x"2454",x"3e2b",x"36eb",x"3902",x"3a23",x"306a",x"3b20",x"3b38",x"242c",x"3e29",x"3712",x"3ae4",x"37c3",x"30c9",x"3b1b",x"3b39",x"2226",x"3e2b",x"3713",x"3607",x"3b5e",x"2e4f",x"3b1b",x"3b3b"),
(x"9e52",x"3df5",x"36eb",x"bbe3",x"ace8",x"30c3",x"3a3c",x"3a6b",x"a088",x"3df5",x"36eb",x"b571",x"bb6d",x"30cc",x"3a3d",x"3a69",x"a05e",x"3df6",x"3713",x"b451",x"bbac",x"2d81",x"3a38",x"3a67"),
(x"9ce6",x"3e67",x"36eb",x"ac58",x"bbf7",x"2bc5",x"3b8d",x"396a",x"a0e1",x"3e67",x"36eb",x"aeda",x"bbea",x"2e47",x"3b8b",x"3969",x"a072",x"3e68",x"3712",x"b297",x"bbcc",x"2d84",x"3b8b",x"396f"),
(x"9dfd",x"3eae",x"36eb",x"b66a",x"3b44",x"2f81",x"3b43",x"3894",x"177f",x"3eb0",x"36eb",x"175f",x"3bf5",x"2e99",x"3b44",x"3890",x"1788",x"3eaf",x"3715",x"1ef6",x"3bee",x"302a",x"3b3f",x"388f"),
(x"11e3",x"3e5e",x"36eb",x"b5a6",x"bb74",x"2d53",x"3b3d",x"384c",x"9470",x"3e5c",x"36eb",x"39cd",x"b979",x"2caa",x"3b3c",x"384b",x"9607",x"3e5d",x"3717",x"3939",x"ba0b",x"29e0",x"3b38",x"384d"),
(x"2164",x"3e2d",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b20",x"3b3c",x"21e1",x"3e2c",x"36eb",x"33f1",x"3bbc",x"2b5c",x"3b20",x"3b3b",x"2226",x"3e2b",x"3713",x"3607",x"3b5e",x"2e4f",x"3b1b",x"3b3b"),
(x"9de0",x"3df4",x"3715",x"2587",x"b07a",x"3beb",x"3b63",x"3b19",x"2043",x"3df7",x"3715",x"99bc",x"26cf",x"3bff",x"3b6f",x"3b19",x"9f80",x"3def",x"3712",x"a9f0",x"ab1d",x"3bfa",x"3b61",x"3b14"),
(x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a",x"1624",x"3e08",x"370e",x"3004",x"271d",x"3bef",x"3b6b",x"3b29",x"2043",x"3df7",x"3715",x"99bc",x"26cf",x"3bff",x"3b6f",x"3b19"),
(x"9e25",x"3df6",x"3716",x"20ea",x"2786",x"3bfe",x"3b63",x"3b1a",x"2043",x"3df7",x"3715",x"99bc",x"26cf",x"3bff",x"3b6f",x"3b19",x"9de0",x"3df4",x"3715",x"2587",x"b07a",x"3beb",x"3b63",x"3b19"),
(x"a08e",x"3e07",x"3717",x"2bf6",x"a5ae",x"3bfb",x"3b62",x"3b29",x"9631",x"3e13",x"3716",x"2adf",x"26b5",x"3bfc",x"3b69",x"3b32",x"1624",x"3e08",x"370e",x"3004",x"271d",x"3bef",x"3b6b",x"3b29"),
(x"9ce6",x"3e67",x"36eb",x"ac58",x"bbf7",x"2bc5",x"3b8d",x"396a",x"9d58",x"3e68",x"3717",x"aa07",x"bbfc",x"284d",x"3b8c",x"3970",x"9b02",x"3e67",x"3716",x"b8f4",x"ba42",x"2c09",x"3b8d",x"3970"),
(x"a395",x"3ea8",x"36eb",x"b9f2",x"3938",x"30b5",x"3b42",x"389a",x"9dfd",x"3eae",x"36eb",x"b66a",x"3b44",x"2f81",x"3b43",x"3894",x"9e4d",x"3ead",x"3713",x"b82e",x"3aba",x"306c",x"3b3f",x"3893"),
(x"1acb",x"3e5c",x"3714",x"b9a7",x"b99e",x"2d1e",x"3b39",x"3850",x"1e07",x"3e59",x"3714",x"b97e",x"b9c5",x"2dbf",x"3b3a",x"3852",x"1e32",x"3e58",x"36eb",x"b976",x"b9cc",x"2dcc",x"3b3f",x"3850"),
(x"11e3",x"3e5e",x"36eb",x"b5a6",x"bb74",x"2d53",x"3b3d",x"384c",x"125b",x"3e5e",x"3717",x"ac95",x"bbf9",x"2918",x"3b38",x"384e",x"1acb",x"3e5c",x"3714",x"b9a7",x"b99e",x"2d1e",x"3b39",x"3850"),
(x"2164",x"3e2d",x"36eb",x"394d",x"b9f2",x"2dc5",x"3b20",x"3b3c",x"212c",x"3e2d",x"3716",x"3ac7",x"b83c",x"283f",x"3b1b",x"3b3d",x"2360",x"3e2f",x"3711",x"38c8",x"ba4e",x"30a8",x"3b1c",x"3b3f"),
(x"a493",x"3e9e",x"36eb",x"bbc4",x"327a",x"3012",x"3b40",x"389e",x"a395",x"3ea8",x"36eb",x"b9f2",x"3938",x"30b5",x"3b42",x"389a",x"a2e7",x"3ea6",x"3715",x"bae0",x"37cf",x"30d4",x"3b3d",x"3898"),
(x"1e32",x"3e58",x"36eb",x"b976",x"b9cc",x"2dcc",x"3b3f",x"3850",x"1e07",x"3e59",x"3714",x"b97e",x"b9c5",x"2dbf",x"3b3a",x"3852",x"2116",x"3e56",x"3716",x"b7d5",x"baf0",x"2d8e",x"3b3b",x"3854"),
(x"2433",x"3e2e",x"36eb",x"39ec",x"b92b",x"31e4",x"3b20",x"3b3f",x"2360",x"3e2f",x"3711",x"38c8",x"ba4e",x"30a8",x"3b1c",x"3b3f",x"24fa",x"3e37",x"370f",x"3b4b",x"b5cc",x"3223",x"3b1c",x"3b44"),
(x"a0ba",x"3def",x"36eb",x"bbdb",x"9c67",x"320a",x"3b8c",x"3a25",x"9f80",x"3def",x"3712",x"bbcf",x"3082",x"3141",x"3b88",x"3a28",x"9e24",x"3de5",x"370e",x"bb7b",x"b4a9",x"3270",x"3b8b",x"3a2c"),
(x"9959",x"3e66",x"3715",x"ba5f",x"3874",x"3388",x"3a37",x"3a24",x"9abe",x"3e63",x"3714",x"387a",x"b47b",x"3a3d",x"3a37",x"3a25",x"9ec5",x"3e5f",x"3718",x"bac6",x"37dc",x"3286",x"3a38",x"3a28"),
(x"a46a",x"3e94",x"36eb",x"bb6e",x"b575",x"309e",x"3b3f",x"38a3",x"a493",x"3e9e",x"36eb",x"bbc4",x"327a",x"3012",x"3b40",x"389e",x"a44d",x"3e9d",x"3715",x"bbec",x"2be2",x"2fce",x"3b3c",x"389d"),
(x"2002",x"3e80",x"3714",x"305e",x"a194",x"3bec",x"3b72",x"3b90",x"2467",x"3e8c",x"3711",x"2cd1",x"a504",x"3bf9",x"3b7a",x"3b9a",x"2353",x"3e7c",x"3711",x"3115",x"a7d5",x"3be4",x"3b78",x"3b8d"),
(x"2002",x"3e80",x"3714",x"305e",x"a194",x"3bec",x"3b72",x"3b90",x"22b8",x"3e8e",x"3713",x"30f4",x"99bc",x"3be7",x"3b77",x"3b9b",x"2467",x"3e8c",x"3711",x"2cd1",x"a504",x"3bf9",x"3b7a",x"3b9a"),
(x"20ef",x"3e55",x"36eb",x"b53f",x"bb87",x"2d28",x"3b40",x"3852",x"2116",x"3e56",x"3716",x"b7d5",x"baf0",x"2d8e",x"3b3b",x"3854",x"2323",x"3e55",x"3716",x"2345",x"bbf7",x"2dcc",x"3b3c",x"3856"),
(x"2563",x"3e37",x"36eb",x"3bbc",x"b212",x"3175",x"3b20",x"3b44",x"24fa",x"3e37",x"370f",x"3b4b",x"b5cc",x"3223",x"3b1c",x"3b44",x"2517",x"3e40",x"370f",x"3bd3",x"2f46",x"3182",x"3b1c",x"3b49"),
(x"a0d7",x"3e5f",x"36eb",x"bafe",x"375c",x"30f4",x"3a3d",x"3a29",x"9ec5",x"3e5f",x"3718",x"bac6",x"37dc",x"3286",x"3a38",x"3a28",x"a29f",x"3e53",x"3714",x"bb6b",x"3587",x"3096",x"3a39",x"3a2f"),
(x"a46a",x"3e94",x"36eb",x"bb6e",x"b575",x"309e",x"3b3f",x"38a3",x"a409",x"3e95",x"3717",x"bb55",x"b5fd",x"307e",x"3b3a",x"38a1",x"a18f",x"3e8e",x"3711",x"b8a4",x"ba69",x"309a",x"3b39",x"38a5"),
(x"2357",x"3e54",x"36eb",x"33e5",x"bbb4",x"2ec2",x"3b41",x"3854",x"2323",x"3e55",x"3716",x"2345",x"bbf7",x"2dcc",x"3b3c",x"3856",x"245f",x"3e57",x"3714",x"3976",x"b9c0",x"3023",x"3b3c",x"3858"),
(x"2574",x"3e41",x"36eb",x"3b61",x"35a0",x"3119",x"3b20",x"3b4a",x"2517",x"3e40",x"370f",x"3bd3",x"2f46",x"3182",x"3b1c",x"3b49",x"2437",x"3e45",x"370f",x"3891",x"3a72",x"30f5",x"3b1b",x"3b4c"),
(x"9f92",x"3de3",x"36eb",x"bade",x"b7ab",x"31d3",x"3b8f",x"3a2a",x"9e24",x"3de5",x"370e",x"bb7b",x"b4a9",x"3270",x"3b8b",x"3a2c",x"0f4a",x"3ddc",x"3712",x"b8b5",x"ba3e",x"32bd",x"3b8d",x"3a32"),
(x"a348",x"3e53",x"36eb",x"bbba",x"3376",x"2f14",x"3a3e",x"3a2f",x"a29f",x"3e53",x"3714",x"bb6b",x"3587",x"3096",x"3a39",x"3a2f",x"a3b3",x"3e47",x"3712",x"bbf0",x"2a00",x"2f46",x"3a3a",x"3a36"),
(x"9bc5",x"3e8b",x"36eb",x"b60d",x"bb5a",x"2ef3",x"3b3a",x"38ab",x"a22e",x"3e8d",x"36eb",x"b884",x"ba69",x"324a",x"3b3d",x"38a8",x"a18f",x"3e8e",x"3711",x"b8a4",x"ba69",x"309a",x"3b39",x"38a5"),
(x"24b8",x"3e56",x"36eb",x"3acc",x"b812",x"3064",x"3b41",x"3856",x"245f",x"3e57",x"3714",x"3976",x"b9c0",x"3023",x"3b3c",x"3858",x"24ba",x"3e5b",x"3712",x"3be0",x"ae5e",x"30a3",x"3b3d",x"385a"),
(x"21a6",x"3e48",x"36eb",x"b5e4",x"3b4d",x"31a2",x"3b1f",x"3b51",x"2449",x"3e47",x"36eb",x"386e",x"3a87",x"313e",x"3b20",x"3b4e",x"2437",x"3e45",x"370f",x"3891",x"3a72",x"30f5",x"3b1b",x"3b4c"),
(x"1dd1",x"3dd9",x"36eb",x"3996",x"b95e",x"33ec",x"3b92",x"3a33",x"1222",x"3dd9",x"36eb",x"b8a6",x"ba54",x"3207",x"3b91",x"3a31",x"0f4a",x"3ddc",x"3712",x"b8b5",x"ba3e",x"32bd",x"3b8d",x"3a32"),
(x"a41c",x"3e46",x"36eb",x"bbef",x"ad09",x"2e69",x"3a3f",x"3a36",x"a3b3",x"3e47",x"3712",x"bbf0",x"2a00",x"2f46",x"3a3a",x"3a36",x"a294",x"3e3b",x"3710",x"bb6a",x"b5bb",x"2efe",x"3a3b",x"3a3c"),
(x"990f",x"3e89",x"36eb",x"bbe6",x"b08f",x"2c41",x"3b3a",x"38ac",x"9bc5",x"3e8b",x"36eb",x"b60d",x"bb5a",x"2ef3",x"3b3a",x"38ab",x"9a89",x"3e8b",x"3718",x"b8ae",x"ba78",x"2b7c",x"3b36",x"38a8"),
(x"2515",x"3e5c",x"36eb",x"3bcf",x"3174",x"303e",x"3b42",x"3859",x"24ba",x"3e5b",x"3712",x"3be0",x"ae5e",x"30a3",x"3b3d",x"385a",x"2458",x"3e5f",x"3714",x"3972",x"39bb",x"30de",x"3b3d",x"385c"),
(x"2467",x"3e8c",x"3711",x"2cd1",x"a504",x"3bf9",x"3b7a",x"3b9a",x"22b8",x"3e8e",x"3713",x"30f4",x"99bc",x"3be7",x"3b77",x"3b9b",x"235a",x"3e97",x"3710",x"a828",x"a60a",x"3bfe",x"3b78",x"3ba3"),
(x"235a",x"3e97",x"3710",x"a828",x"a60a",x"3bfe",x"3b78",x"3ba3",x"2469",x"3e9d",x"3714",x"aeb0",x"a8fa",x"3bf3",x"3b7b",x"3ba9",x"2467",x"3e8c",x"3711",x"2cd1",x"a504",x"3bf9",x"3b7a",x"3b9a"),
(x"23cf",x"3ea5",x"3712",x"2587",x"a09b",x"3bff",x"3b79",x"3baf",x"2325",x"3e9e",x"3714",x"a946",x"9ffc",x"3bfe",x"3b78",x"3baa",x"227e",x"3ea3",x"3712",x"a953",x"a7b4",x"3bfd",x"3b77",x"3bad"),
(x"23cf",x"3ea5",x"3712",x"2587",x"a09b",x"3bff",x"3b79",x"3baf",x"2469",x"3e9d",x"3714",x"aeb0",x"a8fa",x"3bf3",x"3b7b",x"3ba9",x"2325",x"3e9e",x"3714",x"a946",x"9ffc",x"3bfe",x"3b78",x"3baa"),
(x"20a5",x"3eac",x"3715",x"20ea",x"aafd",x"3bfc",x"3b75",x"3bb6",x"23cf",x"3ea5",x"3712",x"2587",x"a09b",x"3bff",x"3b79",x"3baf",x"214b",x"3ea6",x"3714",x"28bf",x"ac22",x"3bfa",x"3b76",x"3bb0"),
(x"1788",x"3eaf",x"3715",x"a7e2",x"a9b5",x"3bfc",x"3b6f",x"3bb9",x"20a5",x"3eac",x"3715",x"20ea",x"aafd",x"3bfc",x"3b75",x"3bb6",x"1f1f",x"3ea8",x"3714",x"a31d",x"ab5f",x"3bfc",x"3b73",x"3bb3"),
(x"9e4d",x"3ead",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3b69",x"3bb7",x"1788",x"3eaf",x"3715",x"a7e2",x"a9b5",x"3bfc",x"3b6f",x"3bb9",x"11db",x"3eaa",x"3715",x"a70a",x"2773",x"3bfe",x"3b6e",x"3bb4"),
(x"a2e7",x"3ea6",x"3715",x"2266",x"1d87",x"3bff",x"3b62",x"3bb2",x"9e4d",x"3ead",x"3713",x"ab1d",x"2ee4",x"3bf0",x"3b69",x"3bb7",x"9d99",x"3ea9",x"3716",x"a4bc",x"2ceb",x"3bf9",x"3b69",x"3bb4"),
(x"a44d",x"3e9d",x"3715",x"2891",x"27ce",x"3bfd",x"3b5f",x"3baa",x"a2e7",x"3ea6",x"3715",x"2266",x"1d87",x"3bff",x"3b62",x"3bb2",x"a14f",x"3ea3",x"3714",x"28e0",x"a99e",x"3bfc",x"3b65",x"3baf"),
(x"a0ed",x"3e98",x"3715",x"2c67",x"a8a5",x"3bf9",x"3b65",x"3ba6",x"a409",x"3e95",x"3717",x"2d06",x"a793",x"3bf8",x"3b60",x"3ba3",x"a44d",x"3e9d",x"3715",x"2891",x"27ce",x"3bfd",x"3b5f",x"3baa"),
(x"a18f",x"3e8e",x"3711",x"28d9",x"252b",x"3bfe",x"3b63",x"3b9d",x"a409",x"3e95",x"3717",x"2d06",x"a793",x"3bf8",x"3b60",x"3ba3",x"a0ed",x"3e98",x"3715",x"2c67",x"a8a5",x"3bf9",x"3b65",x"3ba6"),
(x"1d11",x"3e98",x"3711",x"2bef",x"28a8",x"3bfa",x"3b71",x"3ba4",x"9ddf",x"3e98",x"3714",x"2a45",x"ab10",x"3bfa",x"3b68",x"3ba5",x"9908",x"3e9a",x"3711",x"2a66",x"331a",x"3bca",x"3b6b",x"3ba7"),
(x"9a89",x"3e8b",x"3718",x"2b65",x"3528",x"3b8f",x"3b69",x"3b9a",x"1b8a",x"3e8e",x"3711",x"340c",x"a6c2",x"3bbc",x"3b6f",x"3b9c",x"18c5",x"3e8c",x"3713",x"341f",x"2c3a",x"3bb6",x"3b6e",x"3b9a"),
(x"1832",x"3e87",x"3714",x"2de0",x"24c2",x"3bf6",x"3b6e",x"3b96",x"9747",x"3e88",x"3718",x"3420",x"9418",x"3bba",x"3b6a",x"3b97",x"18c5",x"3e8c",x"3713",x"341f",x"2c3a",x"3bb6",x"3b6e",x"3b9a"),
(x"1832",x"3e87",x"3714",x"2de0",x"24c2",x"3bf6",x"3b6e",x"3b96",x"9613",x"3e7f",x"3715",x"27ae",x"24ea",x"3bfe",x"3b6b",x"3b8f",x"9747",x"3e88",x"3718",x"3420",x"9418",x"3bba",x"3b6a",x"3b97"),
(x"9ddf",x"3e98",x"3714",x"2a45",x"ab10",x"3bfa",x"3b68",x"3ba5",x"1de8",x"3e90",x"3710",x"2856",x"29ab",x"3bfc",x"3b71",x"3b9e",x"a18f",x"3e8e",x"3711",x"28d9",x"252b",x"3bfe",x"3b63",x"3b9d"),
(x"1d11",x"3e98",x"3711",x"2bef",x"28a8",x"3bfa",x"3b71",x"3ba4",x"1ea1",x"3e94",x"3710",x"2a8d",x"a973",x"3bfb",x"3b72",x"3ba2",x"1de8",x"3e90",x"3710",x"2856",x"29ab",x"3bfc",x"3b71",x"3b9e"),
(x"1832",x"3e87",x"3714",x"3bf3",x"2e23",x"2b27",x"3b38",x"3b28",x"18c5",x"3e8c",x"3713",x"3bc2",x"b3a4",x"298a",x"3b39",x"3b2a",x"199d",x"3e8c",x"36eb",x"3bf6",x"aa70",x"2d61",x"3b3e",x"3b29"),
(x"1c29",x"3e7b",x"36eb",x"346a",x"3b91",x"316a",x"3b3c",x"3b21",x"1c29",x"3e7b",x"3718",x"39e5",x"3968",x"0000",x"3b37",x"3b22",x"1832",x"3e87",x"3714",x"3bf3",x"2e23",x"2b27",x"3b38",x"3b28"),
(x"b930",x"3d5c",x"3710",x"bbeb",x"2604",x"3075",x"3a49",x"33c0",x"b92a",x"3d5c",x"3733",x"bb1e",x"251e",x"3748",x"3a49",x"339f",x"b92b",x"3d45",x"3732",x"bb64",x"243f",x"361b",x"3a35",x"33aa"),
(x"b92a",x"3d5c",x"3733",x"bb1e",x"251e",x"3748",x"3a49",x"339f",x"b922",x"3d5c",x"3748",x"b86c",x"29d9",x"3aa7",x"3a48",x"3388",x"b924",x"3d45",x"3749",x"ba3b",x"267a",x"3902",x"3a35",x"3392"),
(x"b922",x"3d5c",x"3748",x"b86c",x"29d9",x"3aa7",x"3a48",x"3388",x"b91b",x"3d5c",x"3749",x"3594",x"2b76",x"3b7b",x"3a48",x"337b",x"b91f",x"3d45",x"374e",x"ac96",x"29b2",x"3bf8",x"3a34",x"3387"),
(x"b91b",x"3d5c",x"3749",x"3594",x"2b76",x"3b7b",x"3a48",x"337b",x"b913",x"3d5c",x"373b",x"3aa1",x"2559",x"3879",x"3a48",x"3369",x"b918",x"3d45",x"374b",x"38f0",x"29d6",x"3a48",x"3a34",x"337b"),
(x"b913",x"3d5c",x"373b",x"381d",x"3a67",x"34eb",x"3bbd",x"39cf",x"b913",x"3d5e",x"373a",x"3ae3",x"2b4f",x"380a",x"3bbc",x"39cf",x"b90e",x"3d5d",x"370e",x"3754",x"3ae5",x"32eb",x"3bc0",x"39d7"),
(x"b913",x"3d5e",x"373a",x"3ae3",x"2b4f",x"380a",x"3bbc",x"39cf",x"b913",x"3d5c",x"373b",x"381d",x"3a67",x"34eb",x"3bbd",x"39cf",x"b91b",x"3d5c",x"3749",x"382b",x"a439",x"3ad3",x"3bbb",x"39cb"),
(x"b913",x"3d5e",x"373a",x"3b64",x"a9cf",x"3612",x"3beb",x"3979",x"b913",x"3d73",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"3978",x"b90f",x"3d73",x"3727",x"3bc1",x"a904",x"33bf",x"3bfb",x"3974"),
(x"b90f",x"3d73",x"3727",x"3bc1",x"a904",x"33bf",x"3bfb",x"3974",x"b90e",x"3d5d",x"370e",x"3bcb",x"a946",x"330f",x"3bea",x"3970",x"b913",x"3d5e",x"373a",x"3b64",x"a9cf",x"3612",x"3beb",x"3979"),
(x"b913",x"3d73",x"373e",x"3a92",x"a9a8",x"388c",x"3bfb",x"3978",x"b913",x"3d5e",x"373a",x"3b64",x"a9cf",x"3612",x"3beb",x"3979",x"b91b",x"3d5e",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"397d"),
(x"b91a",x"3d72",x"374d",x"36b8",x"aa9e",x"3b3f",x"3bfb",x"397c",x"b91b",x"3d5e",x"374a",x"38ae",x"aa28",x"3a79",x"3beb",x"397d",x"b924",x"3d5e",x"374d",x"af62",x"aa90",x"3bef",x"3beb",x"3980"),
(x"b928",x"3d72",x"374d",x"b867",x"a907",x"3aab",x"3bfb",x"3982",x"b922",x"3d72",x"3751",x"a11e",x"aa52",x"3bfd",x"3bfb",x"397f",x"b924",x"3d5e",x"374d",x"af62",x"aa90",x"3bef",x"3beb",x"3980"),
(x"b92f",x"3d72",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"3986",x"b928",x"3d72",x"374d",x"b867",x"a907",x"3aab",x"3bfb",x"3982",x"b92b",x"3d5e",x"3744",x"b96c",x"a921",x"39df",x"3beb",x"3984"),
(x"b935",x"3d73",x"3725",x"bb50",x"a638",x"3678",x"3bfb",x"398b",x"b92f",x"3d72",x"373f",x"baad",x"a687",x"3865",x"3bfb",x"3986",x"b930",x"3d5e",x"3738",x"bb36",x"a61e",x"36e8",x"3beb",x"3986"),
(x"b930",x"3d5e",x"3738",x"b75b",x"bae5",x"32d3",x"3bb7",x"39c3",x"b92a",x"3d5c",x"3733",x"b800",x"ba99",x"3437",x"3bba",x"39c3",x"b930",x"3d5c",x"3710",x"b6ff",x"bb23",x"2f0f",x"3bbd",x"39bd"),
(x"b913",x"3d5c",x"373b",x"3aa1",x"2559",x"3879",x"3a48",x"3369",x"b90c",x"3d45",x"3724",x"3af5",x"1a59",x"37e2",x"3a34",x"3352",x"b912",x"3d45",x"373c",x"3aea",x"2832",x"3802",x"3a34",x"336a"),
(x"b913",x"3d5c",x"373b",x"3aa1",x"2559",x"3879",x"3a48",x"3369",x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e",x"b90c",x"3d45",x"3724",x"3af5",x"1a59",x"37e2",x"3a34",x"3352"),
(x"b91b",x"3d5e",x"374a",x"3544",x"b37e",x"3b51",x"3bb9",x"39cc",x"b91b",x"3d5c",x"3749",x"382b",x"a439",x"3ad3",x"3bbb",x"39cb",x"b922",x"3d5c",x"3748",x"b511",x"b92e",x"398b",x"3bba",x"39c9"),
(x"b922",x"3d5c",x"3748",x"b511",x"b92e",x"398b",x"3bba",x"39c9",x"b92a",x"3d5c",x"3733",x"b800",x"ba99",x"3437",x"3bba",x"39c3",x"b92b",x"3d5e",x"3744",x"b778",x"ba1b",x"3724",x"3bb7",x"39c5"),
(x"b935",x"3d73",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3843",x"b93a",x"3d73",x"3710",x"b30f",x"3bcb",x"2938",x"3b20",x"383f",x"b931",x"3d74",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3842"),
(x"b92f",x"3d72",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3848",x"b935",x"3d73",x"3725",x"b551",x"3b77",x"3051",x"3b22",x"3843",x"b92a",x"3d74",x"3739",x"b604",x"3b4b",x"3149",x"3b22",x"3849"),
(x"b928",x"3d72",x"374d",x"b4d8",x"3aa2",x"3784",x"3b25",x"384c",x"b92f",x"3d72",x"373f",x"b66a",x"3af4",x"349e",x"3b24",x"3848",x"b925",x"3d74",x"3746",x"b589",x"3adc",x"3614",x"3b22",x"384d"),
(x"b91a",x"3d72",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3851",x"b922",x"3d72",x"3751",x"9a8d",x"39ac",x"39a3",x"3b24",x"384f",x"b920",x"3d74",x"374b",x"aa4f",x"39b7",x"3994",x"3b22",x"384f"),
(x"b913",x"3d73",x"373e",x"3a5b",x"3409",x"386a",x"3b1f",x"3854",x"b91a",x"3d72",x"374d",x"35fb",x"37c1",x"3a53",x"3b22",x"3851",x"b919",x"3d74",x"3749",x"3844",x"355f",x"3a35",x"3b21",x"3851"),
(x"b90f",x"3d73",x"3727",x"3b3e",x"b47e",x"3518",x"3b1b",x"3857",x"b913",x"3d73",x"373e",x"3a5b",x"3409",x"386a",x"3b1f",x"3854",x"b913",x"3d74",x"373e",x"3b0f",x"a04d",x"3786",x"3b1e",x"3853"),
(x"b90d",x"3d73",x"3711",x"b36e",x"a40b",x"3bc7",x"3a5b",x"3349",x"b906",x"3d73",x"3713",x"29ab",x"208e",x"3bfd",x"3a5b",x"333d",x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e"),
(x"b92f",x"3d8b",x"372b",x"bbac",x"a891",x"347c",x"3a6f",x"33b1",x"b92a",x"3d74",x"3739",x"bb13",x"a8dd",x"3771",x"3a5c",x"339e",x"b931",x"3d74",x"3710",x"bbea",x"a7ae",x"307d",x"3a5b",x"33c4"),
(x"b92a",x"3d74",x"3739",x"bb13",x"a8dd",x"3771",x"3a5c",x"339e",x"b92c",x"3d8b",x"373a",x"baa5",x"a5fd",x"3872",x"3a6f",x"33a3",x"b925",x"3d8a",x"3749",x"b926",x"a7c8",x"3a1d",x"3a6f",x"3391"),
(x"b920",x"3d74",x"374b",x"b451",x"a960",x"3bb2",x"3a5c",x"3385",x"b925",x"3d74",x"3746",x"b918",x"a84d",x"3a28",x"3a5c",x"338e",x"b925",x"3d8a",x"3749",x"b926",x"a7c8",x"3a1d",x"3a6f",x"3391"),
(x"b919",x"3d74",x"3749",x"3647",x"a97a",x"3b59",x"3a5c",x"3379",x"b920",x"3d74",x"374b",x"b451",x"a960",x"3bb2",x"3a5c",x"3385",x"b91f",x"3d8a",x"374f",x"a812",x"a959",x"3bfd",x"3a6f",x"3385"),
(x"b913",x"3d74",x"373e",x"3ac8",x"a7bb",x"383c",x"3a5c",x"336a",x"b919",x"3d74",x"3749",x"3647",x"a97a",x"3b59",x"3a5c",x"3379",x"b918",x"3d8a",x"374b",x"38ec",x"a7fc",x"3a4c",x"3a6f",x"3378"),
(x"b913",x"3d74",x"373e",x"3ac8",x"a7bb",x"383c",x"3a5c",x"336a",x"b911",x"3d8a",x"373c",x"3ac9",x"a6b5",x"383a",x"3a6f",x"3366",x"b90b",x"3d8a",x"3722",x"3b0f",x"a82c",x"3781",x"3a6f",x"334c"),
(x"b90b",x"3d74",x"371c",x"3aa9",x"a818",x"386b",x"3a5c",x"334a",x"b90b",x"3d8a",x"3722",x"3b0f",x"a82c",x"3781",x"3a6f",x"334c",x"b907",x"3d8a",x"3718",x"38f7",x"a86d",x"3a44",x"3a6f",x"3340"),
(x"b116",x"3d6c",x"3710",x"0000",x"8000",x"3c00",x"3a55",x"2451",x"b116",x"3d64",x"3710",x"0000",x"8000",x"3c00",x"3a4e",x"2451",x"b135",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"24c1"),
(x"b135",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"24c1",x"b135",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"24c1",x"b161",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"255f"),
(x"b161",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"255f",x"b1a1",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2643",x"b1a1",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2643"),
(x"b1a1",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2643",x"b1a1",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2643",x"b1c1",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"26b3"),
(x"b1c1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"26b3",x"b1c1",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"26b3",x"b1fd",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"278b"),
(x"b1fd",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"278b",x"b22d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"281a",x"b22d",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"281a"),
(x"b22d",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"281a",x"b22d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"281a",x"b261",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2878"),
(x"b261",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2878",x"b2aa",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"28fb",x"b2aa",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"28fb"),
(x"b2aa",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"28fb",x"b2aa",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"28fb",x"b2d6",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2949"),
(x"b2d6",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2949",x"b2d6",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2949",x"b326",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4b",x"29d7"),
(x"b326",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4b",x"29d7",x"b34f",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2a20",x"b34f",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2a20"),
(x"b451",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2c3f",x"b50c",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2d8d",x"b50c",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2d8d"),
(x"b451",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2c3f",x"b451",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2c3f",x"b441",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2c23"),
(x"b441",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2c23",x"b441",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"2c23",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b"),
(x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b",x"b34f",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2a20",x"b34f",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2a20"),
(x"b40b",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2b84",x"b3f4",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2b48",x"b413",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"2ba0"),
(x"b3f4",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2b48",x"b3d2",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2b0a",x"b409",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2b7d"),
(x"b3d2",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2b0a",x"b3a5",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2aba",x"b407",x"3d7d",x"3710",x"0000",x"8cea",x"3c00",x"3a63",x"2b76"),
(x"b40b",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2b84",x"b413",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2ba0",x"b413",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2ba0"),
(x"b3f4",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2b48",x"b413",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2ba0",x"b409",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2b7d"),
(x"b3d2",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2b0a",x"b409",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2b7d",x"b407",x"3d53",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2b76"),
(x"b3a5",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"2aba",x"b407",x"3d53",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2b76",x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b"),
(x"b3a5",x"3d85",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"2aba",x"b368",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a68",x"2a4d",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b"),
(x"b50c",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2d8d",x"b50c",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2d8d",x"b526",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2dbb"),
(x"b62a",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2f8b",x"b62a",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2f8b",x"b5ce",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2ee7"),
(x"b5ce",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2ee7",x"b5ce",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2ee7",x"b5bd",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ec9"),
(x"b5bd",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2ec9",x"b5bd",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ec9",x"b5a1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2e97"),
(x"b5a1",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2e97",x"b5a1",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2e97",x"b581",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2e5e"),
(x"b581",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"2e5e",x"b568",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2e30",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b50d",x"3d8e",x"3710",x"0000",x"8000",x"3c00",x"3a72",x"2d8e",x"b4f9",x"3d8c",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"2d6a",x"b4f5",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"2d63"),
(x"b52b",x"3d8d",x"3710",x"0000",x"8000",x"3c00",x"3a72",x"2dc4",x"b4f5",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"2d63",x"b4f2",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2d5e"),
(x"b4f5",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"2d63",x"b4f9",x"3d43",x"3710",x"0000",x"8000",x"3c00",x"3a32",x"2d6a",x"b50d",x"3d41",x"3710",x"0000",x"8000",x"3c00",x"3a30",x"2d8e"),
(x"b4f2",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2d5e",x"b4f5",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"2d63",x"b52b",x"3d42",x"3710",x"0000",x"8000",x"3c00",x"3a31",x"2dc4"),
(x"b568",x"3d46",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"2e32",x"b575",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2e49",x"b575",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2e47"),
(x"b558",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2e14",x"b575",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"2e47",x"b569",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"2e33"),
(x"b568",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"2e32",x"b558",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"2e14",x"b575",x"3d83",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"2e47"),
(x"b558",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"2e14",x"b544",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"2df0",x"b569",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"2e33"),
(x"b4e1",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2d40",x"b51a",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5f",x"2da6",x"b4da",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2d33"),
(x"b4e1",x"3d56",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2d40",x"b4d8",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2d2f",x"b4da",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2d33"),
(x"b51a",x"3d58",x"3710",x"0000",x"8000",x"3c00",x"3a44",x"2da6",x"b4da",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2d33",x"b4f2",x"3d4a",x"3710",x"0000",x"8000",x"3c00",x"3a38",x"2d5e"),
(x"b51a",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5f",x"2da6",x"b528",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2dbf",x"b4f2",x"3d86",x"3710",x"0000",x"8000",x"3c00",x"3a6b",x"2d5e"),
(x"b528",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2dbf",x"b569",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"2e33",x"b544",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"2df0"),
(x"b544",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"2df0",x"b569",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"2e33",x"b528",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2dbf"),
(x"b528",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"2dbf",x"b52c",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2dc5",x"b568",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"2e30"),
(x"b528",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a46",x"2dbf",x"b569",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"2e33",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b526",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"2dbb",x"b52c",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2dc5",x"b52c",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2dc5"),
(x"b52c",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2dc5",x"b52c",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2dc5",x"b568",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"2e30"),
(x"b62a",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2f8b",x"b62a",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2f8b",x"b63d",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2fac"),
(x"b669",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ffc",x"b63d",x"3d74",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"2fac",x"b63d",x"3d5c",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2fac"),
(x"b669",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2ffc",x"b669",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"2ffc",x"b721",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"30a2"),
(x"b72d",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"30ad",x"b721",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"30a2",x"b721",x"3d5e",x"3710",x"0000",x"8000",x"3c00",x"3a49",x"30a2"),
(x"b7c0",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"3130",x"b7c0",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"3130",x"b794",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"3109"),
(x"b794",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"3109",x"b77a",x"3d76",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"30f1",x"b77a",x"3d5a",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30f1"),
(x"b77a",x"3d76",x"3710",x"0000",x"8000",x"3c00",x"3a5d",x"30f1",x"b776",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"30ed",x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed"),
(x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed",x"b776",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"30ed",x"b72d",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"30ad"),
(x"b6fb",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"3080",x"b6ef",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"3075",x"b6f1",x"3d4b",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"3076"),
(x"b721",x"3d59",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30a2",x"b6fb",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"3080",x"b705",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a35",x"3088"),
(x"b6f1",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"3076",x"b6ef",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"3075",x"b6fb",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"3080"),
(x"b705",x"3d89",x"3710",x"0000",x"8000",x"3c00",x"3a6e",x"3088",x"b6fb",x"3d7b",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"3080",x"b721",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5e",x"30a2"),
(x"b73e",x"3d8c",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"30bc",x"b721",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5e",x"30a2",x"b72e",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"30ae"),
(x"b72e",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"30ae",x"b721",x"3d59",x"3710",x"0000",x"8000",x"3c00",x"3a45",x"30a2",x"b73e",x"3d44",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30bc"),
(x"b7c7",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"3135",x"b7c7",x"3d4d",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"3136",x"b7bd",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3d",x"312d"),
(x"b7c7",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"3135",x"b7a4",x"3d87",x"3710",x"0000",x"8000",x"3c00",x"3a6c",x"3117",x"b7bd",x"3d80",x"3710",x"0000",x"8000",x"3c00",x"3a66",x"312d"),
(x"b7a4",x"3d87",x"3710",x"0000",x"8000",x"3c00",x"3a6c",x"3117",x"b783",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"30f9",x"b7a8",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"311a"),
(x"b7a4",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3117",x"b7bd",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3d",x"312d",x"b7a8",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"311a"),
(x"b72e",x"3d5b",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"30ae",x"b77b",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"30f2",x"b776",x"3d57",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"30ed"),
(x"b72e",x"3d75",x"3710",x"0000",x"8000",x"3c00",x"3a5c",x"30ae",x"b72d",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"30ad",x"b776",x"3d78",x"3710",x"0000",x"8000",x"3c00",x"3a60",x"30ed"),
(x"b801",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"316b",x"b7c0",x"3d71",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"3130",x"b7c0",x"3d5f",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"3130"),
(x"b820",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"31a2",x"b801",x"3d73",x"3710",x"0000",x"8000",x"3c00",x"3a5b",x"316b",x"b801",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a48",x"316b"),
(x"b83a",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"31d0",x"b820",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"31a2",x"b820",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"31a2"),
(x"b84a",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"31ed",x"b83a",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"31d0",x"b83a",x"3d48",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"31d0"),
(x"b85e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3211",x"b84a",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a70",x"31ed",x"b84a",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"31ed"),
(x"b865",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"321d",x"b85e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3211",x"b85e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3211"),
(x"b867",x"3d81",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"3222",x"b865",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a6a",x"321d",x"b865",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a39",x"321d"),
(x"b867",x"3d81",x"3710",x"0000",x"8000",x"3c00",x"3a67",x"3222",x"b867",x"3d4f",x"3710",x"0000",x"8000",x"3c00",x"3a3c",x"3222",x"b86e",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"322d"),
(x"b87d",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"3248",x"b86e",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"322d",x"b86e",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"322d"),
(x"b88f",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"3269",x"b87d",x"3d7f",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"3248",x"b87d",x"3d50",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"3248"),
(x"b89e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3284",x"b88f",x"3d84",x"3710",x"0000",x"8000",x"3c00",x"3a69",x"3269",x"b88f",x"3d4c",x"3710",x"0000",x"8000",x"3c00",x"3a3a",x"3269"),
(x"b8a3",x"3d89",x"3710",x"2160",x"1cd0",x"3bff",x"3a6e",x"328d",x"b89e",x"3d88",x"3710",x"0000",x"8000",x"3c00",x"3a6d",x"3284",x"b89e",x"3d47",x"3710",x"0000",x"8000",x"3c00",x"3a36",x"3284"),
(x"b8a3",x"3d89",x"3710",x"2160",x"1cd0",x"3bff",x"3a6e",x"328d",x"b8a3",x"3d47",x"3710",x"2081",x"9ea7",x"3bff",x"3a35",x"328d",x"b907",x"3d5d",x"3713",x"2c13",x"9f5f",x"3bfb",x"3a48",x"333e"),
(x"b8ff",x"3d8a",x"3710",x"2904",x"26d5",x"3bfd",x"3a6f",x"3331",x"b8a3",x"3d89",x"3710",x"2160",x"1cd0",x"3bff",x"3a6e",x"328d",x"b906",x"3d73",x"3713",x"29ab",x"208e",x"3bfd",x"3a5b",x"333d"),
(x"b918",x"3d8a",x"374b",x"270a",x"3bfd",x"287a",x"3bc0",x"3a1e",x"b91f",x"3d8a",x"374f",x"28f4",x"3bfa",x"ac27",x"3bbf",x"3a20",x"b925",x"3d8a",x"3749",x"257a",x"3bfd",x"28f4",x"3bc0",x"3a23"),
(x"b911",x"3d8a",x"373c",x"2504",x"3bff",x"2111",x"3bc3",x"3a1b",x"b925",x"3d8a",x"3749",x"257a",x"3bfd",x"28f4",x"3bc0",x"3a23",x"b92c",x"3d8b",x"373a",x"25e9",x"3bff",x"17c8",x"3bc3",x"3a25"),
(x"b90b",x"3d8a",x"3722",x"2773",x"3bfe",x"22dc",x"3bc8",x"3a19",x"b92c",x"3d8b",x"373a",x"25e9",x"3bff",x"17c8",x"3bc3",x"3a25",x"b92f",x"3d8b",x"372b",x"26c2",x"3bfe",x"24a2",x"3bc6",x"3a27"),
(x"b907",x"3d8a",x"3718",x"25bc",x"3bfe",x"2680",x"3bc9",x"3a17",x"b92f",x"3d8b",x"372b",x"26c2",x"3bfe",x"24a2",x"3bc6",x"3a27",x"b931",x"3d8b",x"3710",x"2418",x"3bff",x"1a24",x"3bcb",x"3a28"),
(x"b924",x"3d45",x"3749",x"1ef6",x"bbff",x"23ef",x"3a5a",x"3a5e",x"b91f",x"3d45",x"374e",x"281b",x"bbe6",x"b0f3",x"3a5b",x"3a5c",x"b918",x"3d45",x"374b",x"2511",x"bbff",x"2259",x"3a5a",x"3a5a"),
(x"b92b",x"3d45",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a55",x"3a61",x"b924",x"3d45",x"3749",x"1ef6",x"bbff",x"23ef",x"3a5a",x"3a5e",x"b912",x"3d45",x"373c",x"184d",x"bbff",x"26c2",x"3a57",x"3a57"),
(x"b931",x"3d45",x"3710",x"9edc",x"bc00",x"9da1",x"3a4f",x"3a63",x"b92b",x"3d45",x"3732",x"9cd0",x"bc00",x"1bfc",x"3a55",x"3a61",x"b90c",x"3d45",x"3724",x"9e3f",x"bbff",x"a00b",x"3a53",x"3a55"),
(x"b1fd",x"3d56",x"36da",x"35da",x"bb72",x"8000",x"3a5f",x"3b8f",x"b22d",x"3d55",x"36da",x"ae8a",x"bbf5",x"8000",x"3a5f",x"3b94",x"b22d",x"3d55",x"3710",x"2c28",x"bbfb",x"0000",x"3a6a",x"3b94"),
(x"b6fb",x"3d54",x"36da",x"38e1",x"3a57",x"0000",x"3a33",x"39d2",x"b6ef",x"3d51",x"36da",x"3be9",x"30b7",x"068d",x"3a33",x"39d5",x"b6ef",x"3d51",x"3710",x"3b57",x"3658",x"868d",x"3a3e",x"39d5"),
(x"b63d",x"3d74",x"36da",x"ab45",x"3bfc",x"0000",x"3a3d",x"3b80",x"b62a",x"3d74",x"36da",x"303b",x"3bed",x"8000",x"3a3d",x"3b7d",x"b62a",x"3d74",x"3710",x"2fbb",x"3bf1",x"0000",x"3a32",x"3b7d"),
(x"b1c1",x"3d5b",x"36da",x"37bd",x"bb00",x"0000",x"3a5f",x"3b88",x"b1fd",x"3d56",x"36da",x"35da",x"bb72",x"8000",x"3a5f",x"3b8f",x"b1fd",x"3d56",x"3710",x"375d",x"bb1a",x"0000",x"3a6a",x"3b8f"),
(x"b906",x"3d45",x"36da",x"224c",x"bbff",x"0000",x"3a44",x"3a53",x"b931",x"3d45",x"36da",x"9e3f",x"bc00",x"0000",x"3a44",x"3a63",x"b931",x"3d45",x"3710",x"9edc",x"bc00",x"9da1",x"3a4f",x"3a63"),
(x"b721",x"3d59",x"36da",x"3711",x"3b2d",x"0000",x"3a33",x"39ca",x"b6fb",x"3d54",x"36da",x"38e1",x"3a57",x"0000",x"3a33",x"39d2",x"b6fb",x"3d54",x"3710",x"37ed",x"3af2",x"0000",x"3a3e",x"39d2"),
(x"b575",x"3d83",x"36da",x"bb59",x"b650",x"8000",x"3a3d",x"3b4e",x"b575",x"3d86",x"36da",x"bab5",x"385c",x"068d",x"3a3d",x"3b4c",x"b575",x"3d86",x"3710",x"bb97",x"350d",x"8000",x"3a32",x"3b4c"),
(x"b1a1",x"3d5c",x"36da",x"314f",x"bbe3",x"0000",x"3a5f",x"3b85",x"b1c1",x"3d5b",x"36da",x"37bd",x"bb00",x"0000",x"3a5f",x"3b88",x"b1c1",x"3d5b",x"3710",x"3680",x"bb4f",x"8000",x"3a6a",x"3b88"),
(x"b72e",x"3d5b",x"36da",x"39a7",x"39a9",x"0000",x"3a33",x"39c7",x"b721",x"3d59",x"36da",x"3711",x"3b2d",x"0000",x"3a33",x"39ca",x"b721",x"3d59",x"3710",x"37a6",x"3b06",x"8000",x"3a3e",x"39ca"),
(x"b62a",x"3d74",x"36da",x"303b",x"3bed",x"8000",x"3a3d",x"3b7d",x"b5ce",x"3d71",x"36da",x"2ae9",x"3bfc",x"8000",x"3a3d",x"3b6a",x"b5ce",x"3d71",x"3710",x"2f26",x"3bf3",x"0000",x"3a32",x"3b6a"),
(x"b161",x"3d5d",x"36da",x"30d8",x"bbe8",x"8000",x"3a5f",x"3b7f",x"b1a1",x"3d5c",x"36da",x"314f",x"bbe3",x"0000",x"3a5f",x"3b85",x"b1a1",x"3d5c",x"3710",x"2ede",x"bbf4",x"0000",x"3a6a",x"3b85"),
(x"b72d",x"3d5d",x"36da",x"3a45",x"b8f8",x"0000",x"3a33",x"39c5",x"b72e",x"3d5b",x"36da",x"39a7",x"39a9",x"0000",x"3a33",x"39c7",x"b72e",x"3d5b",x"3710",x"3b4f",x"367e",x"0000",x"3a3e",x"39c7"),
(x"b5ce",x"3d71",x"36da",x"2ae9",x"3bfc",x"8000",x"3a3d",x"3b6a",x"b5bd",x"3d71",x"36da",x"b6e1",x"3b38",x"0000",x"3a3d",x"3b67",x"b5bd",x"3d71",x"3710",x"b559",x"3b8a",x"0000",x"3a32",x"3b67"),
(x"b135",x"3d5f",x"36da",x"3822",x"bad9",x"8000",x"3a5f",x"3b7b",x"b161",x"3d5d",x"36da",x"30d8",x"bbe8",x"8000",x"3a5f",x"3b7f",x"b161",x"3d5d",x"3710",x"3407",x"bbbd",x"8000",x"3a6a",x"3b7f"),
(x"b721",x"3d5e",x"36da",x"2560",x"bbff",x"8000",x"3a0c",x"3b9a",x"b72d",x"3d5d",x"36da",x"3a45",x"b8f8",x"0000",x"3a0c",x"3b9c",x"b72d",x"3d5d",x"3710",x"3778",x"bb13",x"0000",x"3a17",x"3b9c"),
(x"b5bd",x"3d71",x"36da",x"b6e1",x"3b38",x"0000",x"3a3d",x"3b67",x"b5a1",x"3d75",x"36da",x"b67b",x"3b50",x"0000",x"3a3d",x"3b60",x"b5a1",x"3d75",x"3710",x"b72c",x"3b26",x"8000",x"3a32",x"3b60"),
(x"b93a",x"3d73",x"36da",x"b311",x"3bcd",x"0000",x"3b18",x"3838",x"b931",x"3d74",x"36da",x"b311",x"3bcd",x"0000",x"3b16",x"383b",x"b931",x"3d74",x"3710",x"b3e2",x"3bbf",x"28c2",x"3b1e",x"3842"),
(x"b116",x"3d64",x"36da",x"3b51",x"b675",x"8000",x"3a5f",x"3b76",x"b135",x"3d5f",x"36da",x"3822",x"bad9",x"8000",x"3a5f",x"3b7b",x"b135",x"3d5f",x"3710",x"3934",x"ba13",x"0000",x"3a6a",x"3b7b"),
(x"b568",x"3d46",x"36da",x"b919",x"ba29",x"0000",x"3a0c",x"3b39",x"b575",x"3d4a",x"36da",x"bb97",x"b50d",x"8000",x"3a0c",x"3b3c",x"b575",x"3d4a",x"3710",x"bab5",x"b85c",x"0000",x"3a17",x"3b3c"),
(x"b5a1",x"3d75",x"36da",x"b67b",x"3b50",x"0000",x"3a3d",x"3b60",x"b581",x"3d78",x"36da",x"b89f",x"3a87",x"0000",x"3a3d",x"3b5a",x"b581",x"3d78",x"3710",x"b794",x"3b0b",x"0000",x"3a32",x"3b5a"),
(x"b669",x"3d5d",x"36da",x"a65f",x"bbff",x"0000",x"3a0c",x"3b77",x"b721",x"3d5e",x"36da",x"2560",x"bbff",x"8000",x"3a0c",x"3b9a",x"b721",x"3d5e",x"3710",x"0cea",x"bc00",x"0000",x"3a17",x"3b9a"),
(x"b581",x"3d78",x"36da",x"b89f",x"3a87",x"0000",x"3a3d",x"3b5a",x"b568",x"3d7e",x"36da",x"bb03",x"37b2",x"868d",x"3a3d",x"3b53",x"b568",x"3d7e",x"3710",x"b9f3",x"3958",x"0000",x"3a32",x"3b53"),
(x"b8a3",x"3d47",x"36da",x"2850",x"bbfe",x"8000",x"3a44",x"3a2e",x"b906",x"3d45",x"36da",x"224c",x"bbff",x"0000",x"3a44",x"3a53",x"b906",x"3d45",x"3710",x"2546",x"bbff",x"9624",x"3a4f",x"3a53"),
(x"b63d",x"3d5c",x"36da",x"affc",x"bbf0",x"8000",x"3a0c",x"3b6e",x"b669",x"3d5d",x"36da",x"a65f",x"bbff",x"0000",x"3a0c",x"3b77",x"b669",x"3d5d",x"3710",x"abaa",x"bbfc",x"0000",x"3a17",x"3b77"),
(x"b568",x"3d89",x"36da",x"b810",x"3ae4",x"8000",x"3a3d",x"3b48",x"b558",x"3d8b",x"36da",x"b02d",x"3bee",x"0000",x"3a3d",x"3b44",x"b558",x"3d8b",x"3710",x"b3cc",x"3bc2",x"8000",x"3a32",x"3b44"),
(x"b62a",x"3d5c",x"36da",x"2fb9",x"bbf1",x"0000",x"3a0c",x"3b6b",x"b63d",x"3d5c",x"36da",x"affc",x"bbf0",x"8000",x"3a0c",x"3b6e",x"b63d",x"3d5c",x"3710",x"ab45",x"bbfc",x"0000",x"3a17",x"3b6e"),
(x"b558",x"3d8b",x"36da",x"b02d",x"3bee",x"0000",x"3a3d",x"3b44",x"b544",x"3d8b",x"36da",x"b46b",x"3bb0",x"0000",x"3a3d",x"3b40",x"b544",x"3d8b",x"3710",x"b138",x"3be4",x"0000",x"3a32",x"3b40"),
(x"b575",x"3d4a",x"36da",x"bb97",x"b50d",x"8000",x"3a0c",x"3b3c",x"b575",x"3d4c",x"36da",x"ba67",x"38cb",x"068d",x"3a0c",x"3b3e",x"b575",x"3d4c",x"3710",x"bb59",x"3650",x"8000",x"3a17",x"3b3e"),
(x"b544",x"3d8b",x"36da",x"b46b",x"3bb0",x"0000",x"3a3d",x"3b40",x"b52b",x"3d8d",x"36da",x"b238",x"3bd8",x"8000",x"3a3d",x"3b3b",x"b52b",x"3d8d",x"3710",x"b472",x"3baf",x"0000",x"3a32",x"3b3b"),
(x"b5ce",x"3d5f",x"36da",x"2f26",x"bbf3",x"0000",x"3a0c",x"3b59",x"b62a",x"3d5c",x"36da",x"2fb9",x"bbf1",x"0000",x"3a0c",x"3b6b",x"b62a",x"3d5c",x"3710",x"303b",x"bbed",x"0000",x"3a17",x"3b6b"),
(x"b52b",x"3d8d",x"36da",x"b238",x"3bd8",x"8000",x"3a3d",x"3b3b",x"b50d",x"3d8e",x"36da",x"324a",x"3bd8",x"8000",x"3a3d",x"3b35",x"b50d",x"3d8e",x"3710",x"253f",x"3bff",x"0000",x"3a32",x"3b35"),
(x"b5bd",x"3d5e",x"36da",x"b559",x"bb8a",x"0000",x"3a0c",x"3b56",x"b5ce",x"3d5f",x"36da",x"2f26",x"bbf3",x"0000",x"3a0c",x"3b59",x"b5ce",x"3d5f",x"3710",x"2ae9",x"bbfc",x"0000",x"3a17",x"3b59"),
(x"b50d",x"3d8e",x"36da",x"324a",x"3bd8",x"8000",x"3a3d",x"3b35",x"b4f9",x"3d8c",x"36da",x"3a57",x"38e0",x"8000",x"3a3d",x"3b31",x"b4f9",x"3d8c",x"3710",x"38a5",x"3a82",x"0000",x"3a32",x"3b31"),
(x"b5a1",x"3d5a",x"36da",x"b72c",x"bb26",x"8000",x"3a0c",x"3b50",x"b5bd",x"3d5e",x"36da",x"b559",x"bb8a",x"0000",x"3a0c",x"3b56",x"b5bd",x"3d5e",x"3710",x"b6e1",x"bb38",x"0000",x"3a17",x"3b56"),
(x"b4f9",x"3d8c",x"36da",x"3a57",x"38e0",x"8000",x"3a3d",x"3b31",x"b4f5",x"3d89",x"36da",x"3bc4",x"33a2",x"0000",x"3a3d",x"3b2e",x"b4f5",x"3d89",x"3710",x"3bbb",x"341b",x"8000",x"3a32",x"3b2e"),
(x"b581",x"3d57",x"36da",x"b794",x"bb0b",x"0000",x"3a0c",x"3b4a",x"b5a1",x"3d5a",x"36da",x"b72c",x"bb26",x"8000",x"3a0c",x"3b50",x"b5a1",x"3d5a",x"3710",x"b67b",x"bb50",x"8000",x"3a17",x"3b50"),
(x"b4f5",x"3d89",x"36da",x"3bc4",x"33a2",x"0000",x"3a3d",x"3b2e",x"b4f2",x"3d86",x"36da",x"3a46",x"38f6",x"0000",x"3a3d",x"3b2c",x"b4f2",x"3d86",x"3710",x"3aea",x"3805",x"8000",x"3a32",x"3b2c"),
(x"b931",x"3d74",x"36da",x"bbff",x"a4d0",x"0000",x"3a5a",x"33f3",x"b931",x"3d8b",x"36da",x"bbff",x"a4d0",x"0000",x"3a6e",x"33f9",x"b931",x"3d8b",x"3710",x"bbfe",x"a4d0",x"28c6",x"3a6f",x"33c9"),
(x"b8ff",x"3d8a",x"36da",x"26a7",x"3bff",x"8000",x"3bd5",x"3a14",x"b8a3",x"3d89",x"36da",x"2a59",x"3bfd",x"0000",x"3bd5",x"39f0",x"b8a3",x"3d89",x"3710",x"286a",x"3bfe",x"8000",x"3bcb",x"39f0"),
(x"b568",x"3d51",x"36da",x"b9f3",x"b958",x"0000",x"3a0c",x"3b43",x"b581",x"3d57",x"36da",x"b794",x"bb0b",x"0000",x"3a0c",x"3b4a",x"b581",x"3d57",x"3710",x"b89f",x"ba87",x"0000",x"3a17",x"3b4a"),
(x"b4f2",x"3d86",x"36da",x"3a46",x"38f6",x"0000",x"3a3d",x"3b2c",x"b4da",x"3d7f",x"36da",x"3afc",x"37cc",x"0000",x"3a3d",x"3b25",x"b4da",x"3d7f",x"3710",x"3a4b",x"38ef",x"068d",x"3a32",x"3b25"),
(x"b8a3",x"3d89",x"36da",x"2a59",x"3bfd",x"0000",x"3bd5",x"39f0",x"b89e",x"3d88",x"36da",x"380f",x"3ae4",x"0000",x"3bd5",x"39ee",x"b89e",x"3d88",x"3710",x"36f0",x"3b35",x"0000",x"3bcb",x"39ee"),
(x"b558",x"3d45",x"36da",x"b3cc",x"bbc2",x"8000",x"3a0c",x"3b35",x"b568",x"3d46",x"36da",x"b919",x"ba29",x"0000",x"3a0c",x"3b39",x"b568",x"3d46",x"3710",x"b810",x"bae4",x"0000",x"3a17",x"3b39"),
(x"b4da",x"3d7f",x"36da",x"3afc",x"37cc",x"0000",x"3a3d",x"3b25",x"b4d8",x"3d7c",x"36da",x"3af9",x"b7d7",x"068d",x"3a3d",x"3b22",x"b4d8",x"3d7c",x"3710",x"3be5",x"b11d",x"068d",x"3a32",x"3b22"),
(x"b89e",x"3d88",x"36da",x"380f",x"3ae4",x"0000",x"3bd5",x"39ee",x"b88f",x"3d84",x"36da",x"377a",x"3b12",x"0000",x"3bd5",x"39e7",x"b88f",x"3d84",x"3710",x"380a",x"3ae7",x"0000",x"3bcb",x"39e7"),
(x"b544",x"3d45",x"36da",x"b138",x"bbe4",x"0000",x"3a0c",x"3b31",x"b558",x"3d45",x"36da",x"b3cc",x"bbc2",x"8000",x"3a0c",x"3b35",x"b558",x"3d45",x"3710",x"b02d",x"bbee",x"0000",x"3a17",x"3b35"),
(x"b4d8",x"3d7c",x"36da",x"3af9",x"b7d7",x"068d",x"3a3d",x"3b22",x"b4e1",x"3d7a",x"36da",x"33d2",x"bbc1",x"8000",x"3a3d",x"3b20",x"b4e1",x"3d7a",x"3710",x"3599",x"bb7e",x"0000",x"3a32",x"3b20"),
(x"b88f",x"3d84",x"36da",x"377a",x"3b12",x"0000",x"3bd5",x"39e7",x"b87d",x"3d7f",x"36da",x"3244",x"3bd8",x"0000",x"3bd5",x"39df",x"b87d",x"3d7f",x"3710",x"3541",x"3b8e",x"0000",x"3bcb",x"39df"),
(x"b52b",x"3d42",x"36da",x"b472",x"bbaf",x"0000",x"3a0c",x"3b2c",x"b544",x"3d45",x"36da",x"b138",x"bbe4",x"0000",x"3a0c",x"3b31",x"b544",x"3d45",x"3710",x"b46b",x"bbb0",x"0000",x"3a17",x"3b31"),
(x"b4e1",x"3d7a",x"36da",x"33d2",x"bbc1",x"8000",x"3a3d",x"3b20",x"b51a",x"3d77",x"36da",x"347c",x"bbad",x"0000",x"3a3d",x"3b14",x"b51a",x"3d77",x"3710",x"332b",x"bbcb",x"8000",x"3a32",x"3b14"),
(x"b87d",x"3d7f",x"36da",x"3244",x"3bd8",x"0000",x"3bd5",x"39df",x"b86e",x"3d7f",x"36da",x"b406",x"3bbe",x"0000",x"3bd5",x"39d8",x"b86e",x"3d7f",x"3710",x"ad01",x"3bf9",x"0000",x"3bcb",x"39d8"),
(x"b50d",x"3d41",x"36da",x"253f",x"bbff",x"068d",x"3a0c",x"3b27",x"b52b",x"3d42",x"36da",x"b472",x"bbaf",x"0000",x"3a0c",x"3b2c",x"b52b",x"3d42",x"3710",x"b238",x"bbd8",x"8000",x"3a17",x"3b2c"),
(x"b51a",x"3d77",x"36da",x"347c",x"bbad",x"0000",x"3a3d",x"3b14",x"b528",x"3d75",x"36da",x"38ed",x"ba4d",x"8000",x"3a3d",x"3b11",x"b528",x"3d75",x"3710",x"37fe",x"baed",x"0000",x"3a32",x"3b11"),
(x"b86e",x"3d7f",x"36da",x"b406",x"3bbe",x"0000",x"3bd5",x"39d8",x"b867",x"3d81",x"36da",x"baa2",x"3877",x"0000",x"3bd5",x"39d5",x"b867",x"3d81",x"3710",x"b975",x"39d9",x"0000",x"3bcb",x"39d5"),
(x"b4f9",x"3d43",x"36da",x"38a5",x"ba82",x"8000",x"3a0c",x"3b22",x"b50d",x"3d41",x"36da",x"253f",x"bbff",x"068d",x"3a0c",x"3b27",x"b50d",x"3d41",x"3710",x"324a",x"bbd8",x"8000",x"3a17",x"3b27"),
(x"b528",x"3d75",x"36da",x"38ed",x"ba4d",x"8000",x"3a3d",x"3b11",x"b52c",x"3d74",x"36da",x"3b0d",x"378c",x"0000",x"3a3d",x"3b10",x"b52c",x"3d74",x"3710",x"3bfc",x"ab6c",x"0000",x"3a32",x"3b10"),
(x"b867",x"3d81",x"36da",x"baa2",x"3877",x"0000",x"3bd5",x"39d5",x"b865",x"3d84",x"36da",x"baaf",x"3865",x"8000",x"3bd5",x"39d3",x"b865",x"3d84",x"3710",x"bb0e",x"378a",x"8000",x"3bcb",x"39d3"),
(x"b4f5",x"3d47",x"36da",x"3bbb",x"b41b",x"8000",x"3a0c",x"3b20",x"b4f9",x"3d43",x"36da",x"38a5",x"ba82",x"8000",x"3a0c",x"3b22",x"b4f9",x"3d43",x"3710",x"3a57",x"b8e0",x"0000",x"3a17",x"3b22"),
(x"b52c",x"3d74",x"36da",x"3b0d",x"378c",x"0000",x"3b06",x"39ae",x"b526",x"3d73",x"36da",x"33bb",x"3bc3",x"0000",x"3b06",x"39af",x"b526",x"3d73",x"3710",x"35f8",x"3b6b",x"0000",x"3b11",x"39af"),
(x"b865",x"3d84",x"36da",x"baaf",x"3865",x"8000",x"3bd5",x"39d3",x"b85e",x"3d88",x"36da",x"b5f3",x"3b6d",x"068d",x"3bd5",x"39ce",x"b85e",x"3d88",x"3710",x"b878",x"3aa2",x"0000",x"3bcb",x"39ce"),
(x"b4f2",x"3d4a",x"36da",x"3aea",x"b805",x"8000",x"3a0c",x"3b1d",x"b4f5",x"3d47",x"36da",x"3bbb",x"b41b",x"8000",x"3a0c",x"3b20",x"b4f5",x"3d47",x"3710",x"3bc4",x"b3a2",x"8000",x"3a17",x"3b20"),
(x"b526",x"3d73",x"36da",x"33bb",x"3bc3",x"0000",x"3b06",x"39af",x"b50c",x"3d72",x"36da",x"236c",x"3bff",x"0000",x"3b06",x"39b4",x"b50c",x"3d72",x"3710",x"292b",x"3bfe",x"8000",x"3b11",x"39b4"),
(x"b116",x"3d6c",x"36da",x"3bdf",x"31b0",x"868d",x"3a5f",x"3b70",x"b116",x"3d64",x"36da",x"3b51",x"b675",x"8000",x"3a5f",x"3b76",x"b116",x"3d64",x"3710",x"3bdf",x"b1b0",x"068d",x"3a6a",x"3b76"),
(x"b85e",x"3d88",x"36da",x"b5f3",x"3b6d",x"068d",x"3bd5",x"39ce",x"b84a",x"3d8b",x"36da",x"30e0",x"3be8",x"8000",x"3bd5",x"39c6",x"b84a",x"3d8b",x"3710",x"ac15",x"3bfb",x"8000",x"3bcb",x"39c6"),
(x"b4da",x"3d51",x"36da",x"3a4b",x"b8ef",x"8000",x"3a0c",x"3b17",x"b4f2",x"3d4a",x"36da",x"3aea",x"b805",x"8000",x"3a0c",x"3b1d",x"b4f2",x"3d4a",x"3710",x"3a46",x"b8f6",x"0000",x"3a17",x"3b1d"),
(x"b451",x"3d72",x"36da",x"a987",x"3bfe",x"8000",x"3b06",x"39d8",x"b441",x"3d73",x"36da",x"b7a3",x"3b07",x"0000",x"3b06",x"39db",x"b441",x"3d73",x"3710",x"b6f3",x"3b34",x"0000",x"3b11",x"39db"),
(x"b89e",x"3d47",x"36da",x"36f0",x"bb35",x"0000",x"3a44",x"3a2c",x"b8a3",x"3d47",x"36da",x"2850",x"bbfe",x"8000",x"3a44",x"3a2e",x"b8a3",x"3d47",x"3710",x"2a1e",x"bbfd",x"0000",x"3a4f",x"3a2e"),
(x"b84a",x"3d8b",x"36da",x"30e0",x"3be8",x"8000",x"3bd5",x"39c6",x"b83a",x"3d88",x"36da",x"3953",x"39f7",x"8000",x"3bd5",x"39bf",x"b83a",x"3d88",x"3710",x"3890",x"3a92",x"0000",x"3bcb",x"39bf"),
(x"b4d8",x"3d54",x"36da",x"3be5",x"311d",x"068d",x"3a0c",x"3b14",x"b4da",x"3d51",x"36da",x"3a4b",x"b8ef",x"8000",x"3a0c",x"3b17",x"b4da",x"3d51",x"3710",x"3afc",x"b7cc",x"8000",x"3a17",x"3b17"),
(x"b50c",x"3d72",x"36da",x"236c",x"3bff",x"0000",x"3b06",x"39b4",x"b451",x"3d72",x"36da",x"a987",x"3bfe",x"8000",x"3b06",x"39d8",x"b451",x"3d72",x"3710",x"a0ea",x"3c00",x"0000",x"3b11",x"39d8"),
(x"b88f",x"3d4c",x"36da",x"380a",x"bae7",x"0000",x"3a44",x"3a25",x"b89e",x"3d47",x"36da",x"36f0",x"bb35",x"0000",x"3a44",x"3a2c",x"b89e",x"3d47",x"3710",x"380f",x"bae4",x"0000",x"3a4f",x"3a2c"),
(x"b568",x"3d7e",x"36da",x"bb03",x"37b2",x"868d",x"3a3d",x"3b53",x"b569",x"3d80",x"36da",x"ba4b",x"b8f0",x"0000",x"3a3d",x"3b51",x"b569",x"3d80",x"3710",x"bb2d",x"b70f",x"0000",x"3a32",x"3b51"),
(x"b4e1",x"3d56",x"36da",x"3599",x"3b7e",x"0000",x"3a0c",x"3b12",x"b4d8",x"3d54",x"36da",x"3be5",x"311d",x"068d",x"3a0c",x"3b14",x"b4d8",x"3d54",x"3710",x"3af9",x"37d7",x"868d",x"3a17",x"3b14"),
(x"b441",x"3d73",x"36da",x"b7a3",x"3b07",x"0000",x"3b06",x"39db",x"b40d",x"3d7a",x"36da",x"b8bf",x"3a70",x"068d",x"3b06",x"39e6",x"b40d",x"3d7a",x"3710",x"b83a",x"3aca",x"0000",x"3b11",x"39e6"),
(x"b87d",x"3d50",x"36da",x"3541",x"bb8e",x"0000",x"3a44",x"3a1d",x"b88f",x"3d4c",x"36da",x"380a",x"bae7",x"0000",x"3a44",x"3a25",x"b88f",x"3d4c",x"3710",x"377a",x"bb12",x"8000",x"3a4f",x"3a25"),
(x"b83a",x"3d88",x"36da",x"3953",x"39f7",x"8000",x"3bd5",x"39bf",x"b820",x"3d7a",x"36da",x"385c",x"3ab4",x"0000",x"3bd5",x"39b0",x"b820",x"3d7a",x"3710",x"391f",x"3a25",x"0000",x"3bcb",x"39b0"),
(x"b51a",x"3d58",x"36da",x"332b",x"3bcb",x"0000",x"3a0c",x"3b07",x"b4e1",x"3d56",x"36da",x"3599",x"3b7e",x"0000",x"3a0c",x"3b12",x"b4e1",x"3d56",x"3710",x"33d2",x"3bc1",x"868d",x"3a17",x"3b12"),
(x"b40d",x"3d7a",x"36da",x"b8bf",x"3a70",x"068d",x"3b06",x"39e6",x"b407",x"3d7d",x"36da",x"bbf7",x"2ddb",x"0000",x"3b06",x"39e8",x"b407",x"3d7d",x"3710",x"bb61",x"3629",x"0000",x"3b11",x"39e8"),
(x"b86e",x"3d51",x"36da",x"ad01",x"bbf9",x"0000",x"3a44",x"3a17",x"b87d",x"3d50",x"36da",x"3541",x"bb8e",x"0000",x"3a44",x"3a1d",x"b87d",x"3d50",x"3710",x"3244",x"bbd8",x"0000",x"3a4f",x"3a1d"),
(x"b569",x"3d80",x"36da",x"ba4b",x"b8f0",x"0000",x"3a3d",x"3b51",x"b575",x"3d83",x"36da",x"bb59",x"b650",x"8000",x"3a3d",x"3b4e",x"b575",x"3d83",x"3710",x"ba67",x"b8cb",x"868d",x"3a32",x"3b4e"),
(x"b528",x"3d5a",x"36da",x"37fe",x"3aed",x"0000",x"3a0c",x"3b04",x"b51a",x"3d58",x"36da",x"332b",x"3bcb",x"0000",x"3a0c",x"3b07",x"b51a",x"3d58",x"3710",x"347c",x"3bad",x"8000",x"3a17",x"3b07"),
(x"b407",x"3d7d",x"36da",x"bbf7",x"2ddb",x"0000",x"3b06",x"39e8",x"b409",x"3d7e",x"36da",x"bab5",x"b85b",x"0000",x"3b06",x"39e9",x"b409",x"3d7e",x"3710",x"bb1a",x"b75c",x"8000",x"3b11",x"39e9"),
(x"b867",x"3d4f",x"36da",x"b975",x"b9d8",x"0000",x"3a44",x"3a15",x"b86e",x"3d51",x"36da",x"ad01",x"bbf9",x"0000",x"3a44",x"3a17",x"b86e",x"3d51",x"3710",x"b406",x"bbbe",x"0000",x"3a4f",x"3a17"),
(x"b820",x"3d7a",x"36da",x"385c",x"3ab4",x"0000",x"3bd5",x"39b0",x"b801",x"3d73",x"36da",x"3346",x"3bca",x"0000",x"3bd5",x"39a3",x"b801",x"3d73",x"3710",x"3561",x"3b88",x"0000",x"3bcb",x"39a3"),
(x"b52c",x"3d5b",x"36da",x"3bfc",x"2b6c",x"0000",x"3a0c",x"3b03",x"b528",x"3d5a",x"36da",x"37fe",x"3aed",x"0000",x"3a0c",x"3b04",x"b528",x"3d5a",x"3710",x"38ed",x"3a4d",x"0000",x"3a17",x"3b04"),
(x"b409",x"3d7e",x"36da",x"bab5",x"b85b",x"0000",x"3b06",x"39e9",x"b413",x"3d82",x"36da",x"bba9",x"b499",x"0000",x"3b06",x"39ed",x"b413",x"3d82",x"3710",x"bb08",x"b7a0",x"0000",x"3b11",x"39ed"),
(x"b865",x"3d4c",x"36da",x"bb0e",x"b78a",x"8000",x"3a44",x"3a12",x"b867",x"3d4f",x"36da",x"b975",x"b9d8",x"0000",x"3a44",x"3a15",x"b867",x"3d4f",x"3710",x"baa2",x"b877",x"0000",x"3a4f",x"3a15"),
(x"b801",x"3d73",x"36da",x"3346",x"3bca",x"0000",x"3bd5",x"39a3",x"b7c0",x"3d71",x"36da",x"a984",x"3bfe",x"8000",x"3bd5",x"3996",x"b7c0",x"3d71",x"3710",x"29e3",x"3bfd",x"0000",x"3bcb",x"3996"),
(x"b526",x"3d5d",x"36da",x"35f9",x"bb6b",x"0000",x"3a18",x"3a1a",x"b52c",x"3d5b",x"36da",x"3bfc",x"2b6c",x"0000",x"3a18",x"3a1b",x"b52c",x"3d5b",x"3710",x"3b0d",x"b78c",x"0000",x"3a23",x"3a1b"),
(x"b413",x"3d82",x"36da",x"bba9",x"b499",x"0000",x"3b06",x"39ed",x"b413",x"3d84",x"36da",x"ba12",x"3935",x"868d",x"3b06",x"39ee",x"b413",x"3d84",x"3710",x"bb8c",x"354a",x"8000",x"3b11",x"39ee"),
(x"b85e",x"3d47",x"36da",x"b878",x"baa2",x"0000",x"3a44",x"3a0e",x"b865",x"3d4c",x"36da",x"bb0e",x"b78a",x"8000",x"3a44",x"3a12",x"b865",x"3d4c",x"3710",x"baaf",x"b865",x"8000",x"3a4f",x"3a12"),
(x"b7c0",x"3d71",x"36da",x"a984",x"3bfe",x"8000",x"3bd5",x"3996",x"b794",x"3d73",x"36da",x"b51c",x"3b94",x"0000",x"3bd5",x"398d",x"b794",x"3d73",x"3710",x"b358",x"3bc9",x"0000",x"3bcb",x"398d"),
(x"b50c",x"3d5e",x"36da",x"292b",x"bbfe",x"8000",x"3a18",x"3a15",x"b526",x"3d5d",x"36da",x"35f9",x"bb6b",x"0000",x"3a18",x"3a1a",x"b526",x"3d5d",x"3710",x"33bc",x"bbc3",x"0000",x"3a23",x"3a1a"),
(x"b413",x"3d84",x"36da",x"ba12",x"3935",x"868d",x"3b06",x"39ee",x"b40b",x"3d85",x"36da",x"aabe",x"3bfd",x"868d",x"3b06",x"39f0",x"b40b",x"3d85",x"3710",x"b3aa",x"3bc4",x"8000",x"3b11",x"39f0"),
(x"b84a",x"3d45",x"36da",x"ac15",x"bbfb",x"868d",x"3a44",x"3a06",x"b85e",x"3d47",x"36da",x"b878",x"baa2",x"0000",x"3a44",x"3a0e",x"b85e",x"3d47",x"3710",x"b5f3",x"bb6d",x"8000",x"3a4f",x"3a0e"),
(x"b794",x"3d73",x"36da",x"b51c",x"3b94",x"0000",x"3bd5",x"398d",x"b77a",x"3d76",x"36da",x"b97c",x"39d2",x"0000",x"3bd5",x"3987",x"b77a",x"3d76",x"3710",x"b83f",x"3ac7",x"0000",x"3bcb",x"3987"),
(x"b441",x"3d5d",x"36da",x"b6f3",x"bb34",x"0000",x"3a18",x"39ee",x"b451",x"3d5e",x"36da",x"a0ea",x"bc00",x"0000",x"3a18",x"39f1",x"b451",x"3d5e",x"3710",x"a987",x"bbfe",x"8000",x"3a23",x"39f1"),
(x"b40b",x"3d85",x"36da",x"aabe",x"3bfd",x"868d",x"3b06",x"39f0",x"b3f4",x"3d85",x"36da",x"3408",x"3bbd",x"0000",x"3b06",x"39f3",x"b3f4",x"3d85",x"3710",x"3149",x"3be3",x"0000",x"3b11",x"39f3"),
(x"b83a",x"3d48",x"36da",x"3890",x"ba92",x"0000",x"3a44",x"39ff",x"b84a",x"3d45",x"36da",x"ac15",x"bbfb",x"868d",x"3a44",x"3a06",x"b84a",x"3d45",x"3710",x"30e0",x"bbe8",x"8000",x"3a4f",x"3a06"),
(x"b77a",x"3d76",x"36da",x"b97c",x"39d2",x"0000",x"3bd5",x"3987",x"b776",x"3d78",x"36da",x"bbce",x"b2fb",x"0000",x"3bd5",x"3985",x"b776",x"3d78",x"3710",x"bbee",x"3037",x"0000",x"3bcb",x"3985"),
(x"b451",x"3d5e",x"36da",x"a0ea",x"bc00",x"0000",x"3a18",x"39f1",x"b50c",x"3d5e",x"36da",x"292b",x"bbfe",x"8000",x"3a18",x"3a15",x"b50c",x"3d5e",x"3710",x"236c",x"bbff",x"0000",x"3a23",x"3a15"),
(x"b3f4",x"3d85",x"36da",x"3408",x"3bbd",x"0000",x"3b06",x"39f3",x"b3d2",x"3d83",x"36da",x"abf9",x"3bfc",x"0000",x"3b06",x"39f7",x"b3d2",x"3d83",x"3710",x"2ffb",x"3bf0",x"0000",x"3b11",x"39f7"),
(x"b569",x"3d4f",x"36da",x"bb2d",x"370f",x"0000",x"3a0c",x"3b41",x"b568",x"3d51",x"36da",x"b9f3",x"b958",x"0000",x"3a0c",x"3b43",x"b568",x"3d51",x"3710",x"bb03",x"b7b2",x"0000",x"3a17",x"3b43"),
(x"b776",x"3d78",x"36da",x"bbce",x"b2fb",x"0000",x"3bd5",x"3985",x"b77b",x"3d7a",x"36da",x"b853",x"baba",x"0000",x"3bd5",x"3983",x"b77b",x"3d7a",x"3710",x"b937",x"ba10",x"0000",x"3bcb",x"3983"),
(x"b40d",x"3d55",x"36da",x"b83a",x"baca",x"0000",x"3a18",x"39e3",x"b441",x"3d5d",x"36da",x"b6f3",x"bb34",x"0000",x"3a18",x"39ee",x"b441",x"3d5d",x"3710",x"b7a3",x"bb07",x"0000",x"3a23",x"39ee"),
(x"b3d2",x"3d83",x"36da",x"abf9",x"3bfc",x"0000",x"3b06",x"39f7",x"b3a5",x"3d85",x"36da",x"32b6",x"3bd2",x"0000",x"3b06",x"39fb",x"b3a5",x"3d85",x"3710",x"24fd",x"3bff",x"0000",x"3b11",x"39fb"),
(x"b820",x"3d55",x"36da",x"391f",x"ba25",x"0000",x"3a44",x"39f1",x"b83a",x"3d48",x"36da",x"3890",x"ba92",x"0000",x"3a44",x"39ff",x"b83a",x"3d48",x"3710",x"3953",x"b9f7",x"8000",x"3a4f",x"39ff"),
(x"b77b",x"3d7a",x"36da",x"b853",x"baba",x"0000",x"3a93",x"3ac5",x"b790",x"3d7d",x"36da",x"b461",x"bbb1",x"0000",x"3a93",x"3ac9",x"b790",x"3d7d",x"3710",x"b606",x"bb69",x"0000",x"3a9e",x"3ac9"),
(x"b407",x"3d53",x"36da",x"bb61",x"b629",x"0000",x"3a18",x"39e1",x"b40d",x"3d55",x"36da",x"b83a",x"baca",x"0000",x"3a18",x"39e3",x"b40d",x"3d55",x"3710",x"b8bf",x"ba70",x"8000",x"3a23",x"39e3"),
(x"b3a5",x"3d85",x"36da",x"32b6",x"3bd2",x"0000",x"3b06",x"39fb",x"b368",x"3d82",x"36da",x"3912",x"3a2f",x"8000",x"3b06",x"3a01",x"b368",x"3d82",x"3710",x"37ea",x"3af3",x"8000",x"3b11",x"3a01"),
(x"b575",x"3d4c",x"36da",x"ba67",x"38cb",x"068d",x"3a0c",x"3b3e",x"b569",x"3d4f",x"36da",x"bb2d",x"370f",x"0000",x"3a0c",x"3b41",x"b569",x"3d4f",x"3710",x"ba4b",x"38f0",x"0000",x"3a17",x"3b41"),
(x"b790",x"3d7d",x"36da",x"b461",x"bbb1",x"0000",x"3a93",x"3ac9",x"b7a8",x"3d7e",x"36da",x"b4b8",x"bba4",x"8000",x"3a93",x"3ace",x"b7a8",x"3d7e",x"3710",x"b360",x"bbc8",x"0000",x"3a9e",x"3ace"),
(x"b409",x"3d51",x"36da",x"bb1a",x"375d",x"0000",x"3a18",x"39e0",x"b407",x"3d53",x"36da",x"bb61",x"b629",x"0000",x"3a18",x"39e1",x"b407",x"3d53",x"3710",x"bbf7",x"addb",x"0000",x"3a23",x"39e1"),
(x"b368",x"3d82",x"36da",x"3912",x"3a2f",x"8000",x"3b06",x"3a01",x"b340",x"3d7c",x"36da",x"3b6b",x"35fb",x"8000",x"3b06",x"3a07",x"b340",x"3d7c",x"3710",x"3aba",x"3853",x"0000",x"3b11",x"3a07"),
(x"b801",x"3d5d",x"36da",x"3561",x"bb88",x"0000",x"3a44",x"39e4",x"b820",x"3d55",x"36da",x"391f",x"ba25",x"0000",x"3a44",x"39f1",x"b820",x"3d55",x"3710",x"385c",x"bab4",x"8000",x"3a4f",x"39f1"),
(x"b7a8",x"3d7e",x"36da",x"b4b8",x"bba4",x"8000",x"3a93",x"3ace",x"b7bd",x"3d80",x"36da",x"b821",x"bada",x"8000",x"3a93",x"3ad2",x"b7bd",x"3d80",x"3710",x"b6d2",x"bb3c",x"0000",x"3a9e",x"3ad2"),
(x"b413",x"3d4e",x"36da",x"bb08",x"37a1",x"068d",x"3a18",x"39dc",x"b409",x"3d51",x"36da",x"bb1a",x"375d",x"0000",x"3a18",x"39e0",x"b409",x"3d51",x"3710",x"bab5",x"385b",x"0000",x"3a23",x"39e0"),
(x"b340",x"3d7c",x"36da",x"3b6b",x"35fb",x"8000",x"3b06",x"3a07",x"b33a",x"3d77",x"36da",x"3b88",x"b564",x"8000",x"3b06",x"3a0b",x"b33a",x"3d77",x"3710",x"3bf6",x"ae02",x"868d",x"3b11",x"3a0b"),
(x"b7c0",x"3d5f",x"36da",x"29e3",x"bbfd",x"0000",x"3a44",x"39d8",x"b801",x"3d5d",x"36da",x"3561",x"bb88",x"0000",x"3a44",x"39e4",x"b801",x"3d5d",x"3710",x"3346",x"bbca",x"0000",x"3a4f",x"39e4"),
(x"b7bd",x"3d80",x"36da",x"b821",x"bada",x"8000",x"3a93",x"3ad2",x"b7c7",x"3d82",x"36da",x"bb43",x"b6b4",x"0000",x"3a93",x"3ad5",x"b7c7",x"3d82",x"3710",x"ba01",x"b948",x"8a8d",x"3a9e",x"3ad5"),
(x"b931",x"3d45",x"36da",x"bbff",x"26b5",x"0000",x"3a38",x"33fa",x"b930",x"3d5c",x"36da",x"bbff",x"26b5",x"0000",x"3a4b",x"33f0",x"b930",x"3d5c",x"3710",x"bbeb",x"2604",x"3075",x"3a49",x"33c0"),
(x"b413",x"3d4c",x"36da",x"bb8c",x"b54a",x"8000",x"3a18",x"39db",x"b413",x"3d4e",x"36da",x"bb08",x"37a1",x"068d",x"3a18",x"39dc",x"b413",x"3d4e",x"3710",x"bba9",x"3498",x"0000",x"3a23",x"39dc"),
(x"b33a",x"3d77",x"36da",x"3b88",x"b564",x"8000",x"3b06",x"3a0b",x"b351",x"3d72",x"36da",x"3bb2",x"b458",x"0000",x"3b06",x"3a0f",x"b351",x"3d72",x"3710",x"3b23",x"b738",x"0000",x"3b11",x"3a0f"),
(x"b794",x"3d5d",x"36da",x"b358",x"bbc9",x"0000",x"3a44",x"39cf",x"b7c0",x"3d5f",x"36da",x"29e3",x"bbfd",x"0000",x"3a44",x"39d8",x"b7c0",x"3d5f",x"3710",x"a984",x"bbfe",x"0000",x"3a4f",x"39d8"),
(x"b7c7",x"3d82",x"36da",x"bb43",x"b6b4",x"0000",x"3a93",x"3ad5",x"b7c7",x"3d84",x"36da",x"b744",x"3b20",x"8a8d",x"3a93",x"3ad6",x"b7c7",x"3d84",x"3710",x"b8b7",x"3a76",x"0000",x"3a9e",x"3ad6"),
(x"b40b",x"3d4b",x"36da",x"b3aa",x"bbc4",x"0000",x"3a18",x"39d9",x"b413",x"3d4c",x"36da",x"bb8c",x"b54a",x"8000",x"3a18",x"39db",x"b413",x"3d4c",x"3710",x"ba12",x"b935",x"868d",x"3a23",x"39db"),
(x"b351",x"3d72",x"36da",x"3bb2",x"b458",x"0000",x"3b06",x"3a0f",x"b34f",x"3d70",x"36da",x"3448",x"3bb5",x"0000",x"3b06",x"3a11",x"b34f",x"3d70",x"3710",x"3913",x"3a2f",x"0000",x"3b11",x"3a11"),
(x"b77a",x"3d5a",x"36da",x"b83f",x"bac7",x"0000",x"3a44",x"39ca",x"b794",x"3d5d",x"36da",x"b358",x"bbc9",x"0000",x"3a44",x"39cf",x"b794",x"3d5d",x"3710",x"b51c",x"bb94",x"0000",x"3a4f",x"39cf"),
(x"b7c7",x"3d84",x"36da",x"b744",x"3b20",x"8a8d",x"3a93",x"3ad6",x"b7a4",x"3d87",x"36da",x"b64a",x"3b5a",x"8000",x"3a93",x"3add",x"b7a4",x"3d87",x"3710",x"b654",x"3b58",x"0000",x"3a9e",x"3add"),
(x"b3f4",x"3d4b",x"36da",x"3149",x"bbe3",x"0000",x"3a18",x"39d6",x"b40b",x"3d4b",x"36da",x"b3aa",x"bbc4",x"0000",x"3a18",x"39d9",x"b40b",x"3d4b",x"3710",x"aabe",x"bbfd",x"068d",x"3a23",x"39d9"),
(x"b34f",x"3d70",x"36da",x"3448",x"3bb5",x"0000",x"3a5f",x"3b35",x"b326",x"3d70",x"36da",x"ad8e",x"3bf8",x"0000",x"3a5f",x"3b39",x"b326",x"3d70",x"3710",x"a5e3",x"3bff",x"0000",x"3a6a",x"3b39"),
(x"b776",x"3d57",x"36da",x"bbee",x"b037",x"0000",x"3a33",x"3a17",x"b77a",x"3d5a",x"36da",x"b83f",x"bac7",x"0000",x"3a33",x"3a19",x"b77a",x"3d5a",x"3710",x"b97c",x"b9d2",x"0000",x"3a3e",x"3a19"),
(x"b7a4",x"3d87",x"36da",x"b64a",x"3b5a",x"8000",x"3a93",x"3add",x"b783",x"3d8b",x"36da",x"afa0",x"3bf1",x"0000",x"3a93",x"3ae4",x"b783",x"3d8b",x"3710",x"b33d",x"3bca",x"0000",x"3a9e",x"3ae4"),
(x"b3d2",x"3d4c",x"36da",x"2ffb",x"bbf0",x"0000",x"3a18",x"39d2",x"b3f4",x"3d4b",x"36da",x"3149",x"bbe3",x"0000",x"3a18",x"39d6",x"b3f4",x"3d4b",x"3710",x"3408",x"bbbd",x"0000",x"3a23",x"39d6"),
(x"b326",x"3d70",x"36da",x"ad8e",x"3bf8",x"0000",x"3a5f",x"3b39",x"b2d6",x"3d71",x"36da",x"b4dc",x"3b9f",x"0000",x"3a5f",x"3b40",x"b2d6",x"3d71",x"3710",x"b287",x"3bd4",x"0000",x"3a6a",x"3b40"),
(x"b77b",x"3d55",x"36da",x"b937",x"3a10",x"8000",x"3a33",x"3a15",x"b776",x"3d57",x"36da",x"bbee",x"b037",x"0000",x"3a33",x"3a17",x"b776",x"3d57",x"3710",x"bbce",x"32fb",x"0000",x"3a3e",x"3a17"),
(x"b783",x"3d8b",x"36da",x"afa0",x"3bf1",x"0000",x"3a93",x"3ae4",x"b73e",x"3d8c",x"36da",x"2f57",x"3bf2",x"8000",x"3a93",x"3af1",x"b73e",x"3d8c",x"3710",x"27ae",x"3bfe",x"0000",x"3a9e",x"3af1"),
(x"b3a5",x"3d4b",x"36da",x"2504",x"bbff",x"0000",x"3a18",x"39ce",x"b3d2",x"3d4c",x"36da",x"2ffb",x"bbf0",x"0000",x"3a18",x"39d2",x"b3d2",x"3d4c",x"3710",x"abf9",x"bbfc",x"8000",x"3a23",x"39d2"),
(x"b2d6",x"3d71",x"36da",x"b4dc",x"3b9f",x"0000",x"3a5f",x"3b40",x"b2aa",x"3d74",x"36da",x"b7e2",x"3af5",x"0000",x"3a5f",x"3b45",x"b2aa",x"3d74",x"3710",x"b78b",x"3b0e",x"0000",x"3a6a",x"3b45"),
(x"b790",x"3d52",x"36da",x"b606",x"3b69",x"0000",x"3a33",x"3a11",x"b77b",x"3d55",x"36da",x"b937",x"3a10",x"8000",x"3a33",x"3a15",x"b77b",x"3d55",x"3710",x"b853",x"3aba",x"0000",x"3a3e",x"3a15"),
(x"b73e",x"3d8c",x"36da",x"2f57",x"3bf2",x"8000",x"3a93",x"3af1",x"b705",x"3d89",x"36da",x"36ee",x"3b35",x"0000",x"3a93",x"3afc",x"b705",x"3d89",x"3710",x"34b8",x"3ba4",x"0000",x"3a9e",x"3afc"),
(x"b368",x"3d4e",x"36da",x"37ea",x"baf3",x"8000",x"3a18",x"39c8",x"b3a5",x"3d4b",x"36da",x"2504",x"bbff",x"0000",x"3a18",x"39ce",x"b3a5",x"3d4b",x"3710",x"32b6",x"bbd2",x"868d",x"3a23",x"39ce"),
(x"b2aa",x"3d74",x"36da",x"b7e2",x"3af5",x"0000",x"3a5f",x"3b45",x"b261",x"3d79",x"36da",x"b5e0",x"3b70",x"8000",x"3a5f",x"3b4d",x"b261",x"3d79",x"3710",x"b72e",x"3b26",x"8000",x"3a6a",x"3b4d"),
(x"b7a8",x"3d51",x"36da",x"b360",x"3bc8",x"8000",x"3a33",x"3a0c",x"b790",x"3d52",x"36da",x"b606",x"3b69",x"0000",x"3a33",x"3a11",x"b790",x"3d52",x"3710",x"b461",x"3bb1",x"0000",x"3a3e",x"3a11"),
(x"b705",x"3d89",x"36da",x"36ee",x"3b35",x"0000",x"3a93",x"3afc",x"b6f1",x"3d84",x"36da",x"3b73",x"35d3",x"8000",x"3a93",x"3b01",x"b6f1",x"3d84",x"3710",x"3a69",x"38c9",x"068d",x"3a9e",x"3b01"),
(x"b340",x"3d54",x"36da",x"3aba",x"b853",x"8000",x"3a18",x"39c2",x"b368",x"3d4e",x"36da",x"37ea",x"baf3",x"8000",x"3a18",x"39c8",x"b368",x"3d4e",x"3710",x"3912",x"ba2f",x"8000",x"3a23",x"39c8"),
(x"b261",x"3d79",x"36da",x"b5e0",x"3b70",x"8000",x"3a5f",x"3b4d",x"b22d",x"3d7b",x"36da",x"2c28",x"3bfb",x"0000",x"3a5f",x"3b52",x"b22d",x"3d7b",x"3710",x"ae88",x"3bf5",x"0000",x"3a6a",x"3b52"),
(x"b7bd",x"3d4f",x"36da",x"b6d2",x"3b3c",x"0000",x"3a33",x"3a08",x"b7a8",x"3d51",x"36da",x"b360",x"3bc8",x"8000",x"3a33",x"3a0c",x"b7a8",x"3d51",x"3710",x"b4b8",x"3ba4",x"8000",x"3a3e",x"3a0c"),
(x"b6f1",x"3d84",x"36da",x"3b73",x"35d3",x"8000",x"3a93",x"3b01",x"b6ef",x"3d7f",x"36da",x"3b57",x"b658",x"8000",x"3a93",x"3b05",x"b6ef",x"3d7f",x"3710",x"3be9",x"b0b7",x"0000",x"3a9e",x"3b05"),
(x"b33a",x"3d59",x"36da",x"3bf6",x"2e02",x"8000",x"3a18",x"39be",x"b340",x"3d54",x"36da",x"3aba",x"b853",x"8000",x"3a18",x"39c2",x"b340",x"3d54",x"3710",x"3b6b",x"b5fb",x"0000",x"3a23",x"39c2"),
(x"b22d",x"3d7b",x"36da",x"2c28",x"3bfb",x"0000",x"3a5f",x"3b52",x"b1fd",x"3d79",x"36da",x"375d",x"3b1a",x"8000",x"3a5f",x"3b57",x"b1fd",x"3d79",x"3710",x"35da",x"3b72",x"0000",x"3a6a",x"3b57"),
(x"b7c7",x"3d4d",x"36da",x"ba01",x"3948",x"8000",x"3a33",x"3a06",x"b7bd",x"3d4f",x"36da",x"b6d2",x"3b3c",x"0000",x"3a33",x"3a08",x"b7bd",x"3d4f",x"3710",x"b821",x"3ad9",x"0000",x"3a3e",x"3a08"),
(x"b6ef",x"3d7f",x"36da",x"3b57",x"b658",x"8000",x"3a93",x"3b05",x"b6fb",x"3d7b",x"36da",x"37ed",x"baf2",x"868d",x"3a93",x"3b08",x"b6fb",x"3d7b",x"3710",x"38e1",x"ba57",x"0000",x"3a9e",x"3b08"),
(x"b351",x"3d5d",x"36da",x"3b23",x"3738",x"0000",x"3a18",x"39ba",x"b33a",x"3d59",x"36da",x"3bf6",x"2e02",x"8000",x"3a18",x"39be",x"b33a",x"3d59",x"3710",x"3b88",x"3564",x"868d",x"3a23",x"39be"),
(x"b1fd",x"3d79",x"36da",x"375d",x"3b1a",x"8000",x"3a5f",x"3b57",x"b1c1",x"3d75",x"36da",x"367f",x"3b4f",x"8000",x"3a5f",x"3b5d",x"b1c1",x"3d75",x"3710",x"37bc",x"3b00",x"0000",x"3a6a",x"3b5d"),
(x"b7c7",x"3d4c",x"36da",x"b8b7",x"ba76",x"0000",x"3a33",x"3a05",x"b7c7",x"3d4d",x"36da",x"ba01",x"3948",x"8000",x"3a33",x"3a06",x"b7c7",x"3d4d",x"3710",x"bb43",x"36b4",x"0000",x"3a3e",x"3a06"),
(x"b6fb",x"3d7b",x"36da",x"37ed",x"baf2",x"868d",x"3a93",x"3b08",x"b721",x"3d77",x"36da",x"37a6",x"bb06",x"0000",x"3a93",x"3b10",x"b721",x"3d77",x"3710",x"3711",x"bb2d",x"0000",x"3a9e",x"3b10"),
(x"b34f",x"3d60",x"36da",x"3913",x"ba2f",x"0000",x"3a18",x"39b8",x"b351",x"3d5d",x"36da",x"3b23",x"3738",x"0000",x"3a18",x"39ba",x"b351",x"3d5d",x"3710",x"3bb2",x"3458",x"8000",x"3a23",x"39ba"),
(x"b1c1",x"3d75",x"36da",x"367f",x"3b4f",x"8000",x"3a5f",x"3b5d",x"b1a1",x"3d73",x"36da",x"2ede",x"3bf4",x"0000",x"3a5f",x"3b60",x"b1a1",x"3d73",x"3710",x"314f",x"3be3",x"8000",x"3a6a",x"3b60"),
(x"b7a4",x"3d48",x"36da",x"b654",x"bb58",x"8000",x"3a33",x"39fd",x"b7c7",x"3d4c",x"36da",x"b8b7",x"ba76",x"0000",x"3a33",x"3a05",x"b7c7",x"3d4c",x"3710",x"b744",x"bb20",x"0000",x"3a3e",x"3a05"),
(x"b721",x"3d77",x"36da",x"37a6",x"bb06",x"0000",x"3a93",x"3b10",x"b72e",x"3d75",x"36da",x"3b4f",x"b67e",x"8000",x"3a93",x"3b13",x"b72e",x"3d75",x"3710",x"39a7",x"b9a8",x"0000",x"3a9e",x"3b13"),
(x"b326",x"3d60",x"36da",x"a5e3",x"bbff",x"0000",x"3a5f",x"3bad",x"b34f",x"3d60",x"36da",x"3913",x"ba2f",x"0000",x"3a5f",x"3bb1",x"b34f",x"3d60",x"3710",x"3448",x"bbb5",x"0000",x"3a6a",x"3bb1"),
(x"b1a1",x"3d73",x"36da",x"2ede",x"3bf4",x"0000",x"3a5f",x"3b60",x"b161",x"3d73",x"36da",x"3408",x"3bbd",x"0000",x"3a5f",x"3b66",x"b161",x"3d73",x"3710",x"30d8",x"3be8",x"8000",x"3a6a",x"3b66"),
(x"b783",x"3d45",x"36da",x"b33d",x"bbca",x"8000",x"3a33",x"39f7",x"b7a4",x"3d48",x"36da",x"b654",x"bb58",x"8000",x"3a33",x"39fd",x"b7a4",x"3d48",x"3710",x"b64a",x"bb5a",x"0000",x"3a3e",x"39fd"),
(x"b72e",x"3d75",x"36da",x"3b4f",x"b67e",x"8000",x"3a3d",x"3bb1",x"b72d",x"3d73",x"36da",x"3778",x"3b13",x"0000",x"3a3d",x"3bb0",x"b72d",x"3d73",x"3710",x"3a45",x"38f8",x"0000",x"3a32",x"3bb0"),
(x"b2d6",x"3d5f",x"36da",x"b287",x"bbd4",x"0000",x"3a5f",x"3ba5",x"b326",x"3d60",x"36da",x"a5e3",x"bbff",x"0000",x"3a5f",x"3bad",x"b326",x"3d60",x"3710",x"ad8e",x"bbf8",x"0000",x"3a6a",x"3bad"),
(x"b161",x"3d73",x"36da",x"3408",x"3bbd",x"0000",x"3a5f",x"3b66",x"b135",x"3d71",x"36da",x"3934",x"3a13",x"8000",x"3a5f",x"3b6b",x"b135",x"3d71",x"3710",x"3822",x"3ad9",x"0000",x"3a6a",x"3b6b"),
(x"b73e",x"3d44",x"36da",x"27ae",x"bbff",x"0000",x"3a33",x"39ea",x"b783",x"3d45",x"36da",x"b33d",x"bbca",x"8000",x"3a33",x"39f7",x"b783",x"3d45",x"3710",x"afa0",x"bbf1",x"0000",x"3a3e",x"39f7"),
(x"b72d",x"3d73",x"36da",x"3778",x"3b13",x"0000",x"3a3d",x"3bb0",x"b721",x"3d72",x"36da",x"0cea",x"3c00",x"0000",x"3a3d",x"3bad",x"b721",x"3d72",x"3710",x"2560",x"3bff",x"0000",x"3a32",x"3bad"),
(x"b2aa",x"3d5c",x"36da",x"b78b",x"bb0e",x"0000",x"3a5f",x"3ba1",x"b2d6",x"3d5f",x"36da",x"b287",x"bbd4",x"0000",x"3a5f",x"3ba5",x"b2d6",x"3d5f",x"3710",x"b4dc",x"bb9f",x"0000",x"3a6a",x"3ba5"),
(x"b135",x"3d71",x"36da",x"3934",x"3a13",x"8000",x"3a5f",x"3b6b",x"b116",x"3d6c",x"36da",x"3bdf",x"31b0",x"868d",x"3a5f",x"3b70",x"b116",x"3d6c",x"3710",x"3b51",x"3675",x"0000",x"3a6a",x"3b70"),
(x"b705",x"3d47",x"36da",x"34b8",x"bba4",x"868d",x"3a33",x"39de",x"b73e",x"3d44",x"36da",x"27ae",x"bbff",x"0000",x"3a33",x"39ea",x"b73e",x"3d44",x"3710",x"2f57",x"bbf2",x"0000",x"3a3e",x"39ea"),
(x"b575",x"3d86",x"36da",x"bab5",x"385c",x"068d",x"3a3d",x"3b4c",x"b568",x"3d89",x"36da",x"b810",x"3ae4",x"8000",x"3a3d",x"3b48",x"b568",x"3d89",x"3710",x"b919",x"3a29",x"0000",x"3a32",x"3b48"),
(x"b938",x"3d5e",x"36da",x"bbfe",x"a8f0",x"0000",x"3bea",x"3999",x"b93a",x"3d73",x"36da",x"bbfe",x"a8f0",x"0000",x"3bfb",x"3999",x"b93a",x"3d73",x"3710",x"bbf8",x"a8ed",x"2cf7",x"3bfb",x"398f"),
(x"b261",x"3d57",x"36da",x"b72e",x"bb26",x"0000",x"3a5f",x"3b99",x"b2aa",x"3d5c",x"36da",x"b78b",x"bb0e",x"0000",x"3a5f",x"3ba1",x"b2aa",x"3d5c",x"3710",x"b7e2",x"baf5",x"0000",x"3a6a",x"3ba1"),
(x"b931",x"3d8b",x"36da",x"23ae",x"3bff",x"0000",x"3bd5",x"3a28",x"b8ff",x"3d8a",x"36da",x"26a7",x"3bff",x"8000",x"3bd5",x"3a14",x"b8ff",x"3d8a",x"3710",x"257a",x"3bff",x"15bc",x"3bcb",x"3a14"),
(x"b6f1",x"3d4b",x"36da",x"3a69",x"b8c9",x"8000",x"3a33",x"39d9",x"b705",x"3d47",x"36da",x"34b8",x"bba4",x"868d",x"3a33",x"39de",x"b705",x"3d47",x"3710",x"36ee",x"bb35",x"0000",x"3a3e",x"39de"),
(x"b721",x"3d72",x"36da",x"0cea",x"3c00",x"0000",x"3a3d",x"3bad",x"b669",x"3d72",x"36da",x"abae",x"3bfc",x"8000",x"3a3d",x"3b89",x"b669",x"3d72",x"3710",x"a666",x"3bff",x"0000",x"3a32",x"3b89"),
(x"b22d",x"3d55",x"36da",x"ae8a",x"bbf5",x"8000",x"3a5f",x"3b94",x"b261",x"3d57",x"36da",x"b72e",x"bb26",x"0000",x"3a5f",x"3b99",x"b261",x"3d57",x"3710",x"b5e0",x"bb70",x"8000",x"3a6a",x"3b99"),
(x"b6ef",x"3d51",x"36da",x"3be9",x"30b7",x"068d",x"3a33",x"39d5",x"b6f1",x"3d4b",x"36da",x"3a69",x"b8c9",x"8000",x"3a33",x"39d9",x"b6f1",x"3d4b",x"3710",x"3b73",x"b5d3",x"0000",x"3a3e",x"39d9"),
(x"b669",x"3d72",x"36da",x"abae",x"3bfc",x"8000",x"3a3d",x"3b89",x"b63d",x"3d74",x"36da",x"ab45",x"3bfc",x"0000",x"3a3d",x"3b80",x"b63d",x"3d74",x"3710",x"affc",x"3bf0",x"0000",x"3a32",x"3b80"),
(x"b930",x"3d5c",x"36da",x"b67a",x"bb50",x"0000",x"3bc3",x"39b4",x"b938",x"3d5e",x"36da",x"b67a",x"bb50",x"0000",x"3bc0",x"39b2",x"b938",x"3d5e",x"3710",x"b678",x"bb4d",x"2af3",x"3bba",x"39ba"),
(x"b40d",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"2b8b",x"b368",x"4054",x"3710",x"0000",x"8000",x"3c00",x"39e3",x"2a4d",x"b351",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2a24"),
(x"b34f",x"4043",x"3710",x"0000",x"8000",x"3c00",x"39c6",x"2a20",x"b351",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2a27",x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b"),
(x"b34f",x"3d70",x"3710",x"0000",x"8000",x"3c00",x"3a59",x"2a20",x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b",x"b351",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2a22"),
(x"b368",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2a4d",x"b351",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2a27",x"b340",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2a0e"),
(x"b34f",x"3d60",x"3710",x"0000",x"8000",x"3c00",x"3a4a",x"2a20",x"b351",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2a27",x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b"),
(x"b77b",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"30f2",x"b790",x"3d7d",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"3107",x"b783",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"30f9"),
(x"b77b",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"30f2",x"b783",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30f9",x"b790",x"3d52",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"3107"),
(x"b351",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2a27",x"b33a",x"4040",x"3710",x"0000",x"8000",x"3c00",x"39bf",x"2a03",x"b340",x"403d",x"3710",x"0000",x"8000",x"3c00",x"39bb",x"2a0d"),
(x"b783",x"4036",x"3710",x"0000",x"8000",x"3c00",x"39af",x"30f9",x"b7a8",x"403c",x"3710",x"0000",x"8000",x"3c00",x"39ba",x"311a",x"b790",x"403d",x"3710",x"0000",x"8000",x"3c00",x"39bc",x"3107"),
(x"b783",x"4059",x"3710",x"0000",x"8000",x"3c00",x"39eb",x"30f9",x"b77b",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39dd",x"30f2",x"b790",x"4052",x"3710",x"0000",x"8000",x"3c00",x"39de",x"3107"),
(x"b340",x"3d7c",x"3710",x"0000",x"8000",x"3c00",x"3a63",x"2a04",x"b33a",x"3d77",x"3710",x"0000",x"8000",x"3c00",x"3a5e",x"29f9",x"b351",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2a22"),
(x"b340",x"4051",x"3710",x"0000",x"8000",x"3c00",x"39de",x"2a05",x"b33a",x"404f",x"3710",x"0000",x"8000",x"3c00",x"39da",x"29fa",x"b351",x"404d",x"3710",x"0000",x"8000",x"3c00",x"39d6",x"2a24"),
(x"b351",x"4042",x"3710",x"0000",x"8000",x"3c00",x"39c2",x"2a27",x"b368",x"403a",x"3710",x"0000",x"8000",x"3c00",x"39b7",x"2a4d",x"b40d",x"403e",x"3710",x"0000",x"8000",x"3c00",x"39bd",x"2b8b"),
(x"b40d",x"3d7a",x"3710",x"0000",x"8000",x"3c00",x"3a61",x"2b8b",x"b368",x"3d82",x"3710",x"0000",x"8000",x"3c00",x"3a68",x"2a4d",x"b351",x"3d72",x"3710",x"0000",x"8000",x"3c00",x"3a5a",x"2a22"),
(x"b351",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2a27",x"b33a",x"3d59",x"3710",x"0000",x"8000",x"3c00",x"3a43",x"2a04",x"b340",x"3d54",x"3710",x"0000",x"8000",x"3c00",x"3a40",x"2a0e"),
(x"b351",x"3d5d",x"3710",x"0000",x"8000",x"3c00",x"3a47",x"2a27",x"b368",x"3d4e",x"3710",x"0000",x"8000",x"3c00",x"3a3b",x"2a4d",x"b40d",x"3d55",x"3710",x"0000",x"8000",x"3c00",x"3a42",x"2b8b"),
(x"b790",x"3d7d",x"3710",x"0000",x"8000",x"3c00",x"3a62",x"3107",x"b7a8",x"3d7e",x"3710",x"0000",x"8000",x"3c00",x"3a65",x"311a",x"b783",x"3d8b",x"3710",x"0000",x"8000",x"3c00",x"3a6f",x"30f9"),
(x"b783",x"3d45",x"3710",x"0000",x"8000",x"3c00",x"3a33",x"30f9",x"b7a8",x"3d51",x"3710",x"0000",x"8000",x"3c00",x"3a3e",x"311a",x"b790",x"3d52",x"3710",x"0000",x"8000",x"3c00",x"3a41",x"3107"),
others => empty_m_tri);

end model_presets;

package body model_presets is

end model_presets;
