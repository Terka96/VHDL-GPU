----------------------------------------------------------------------------------
-- Copyright 2020 Piotr Terczyński
--
-- Permission is hereby granted, free of charge, to any person
-- obtaining a copy of this software and associated           
-- documentation files (the "Software"), to deal in the       
-- Software without restriction, including without limitation 
-- the rights to use, copy, modify, merge, publish,           
-- distribute, sublicense, and/or sell copies of the Software,
-- and to permit persons to whom the Software is furnished to
-- do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice 
-- shall be included in all copies or substantial portions of
-- the Software.
--
-- 		THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF 
-- ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO 
-- THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR
-- PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS 
-- OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR   
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR 
-- OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE 
-- SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.definitions.all;

package texture is

constant TEX_SIZE_F : FLOAT16 := x"6000";
constant TEX_SIZE	: integer := 512;
constant TEX_MODULO : std_logic_vector(12 downto 0) := "0000111111111";
type TEXTURE_MEM_LINE is array (0 to (TEX_SIZE-1)) of COLOR24;
type TEXTURE_MEM is array (0 to (TEX_SIZE-1)) of TEXTURE_MEM_LINE;

constant texture_memory_const : TEXTURE_MEM := (
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"685646",x"685646",x"5c4e41",x"5e5043",x"564a3d",x"54483e",x"554a3f",x"584c40",x"574b40",x"584c41",x"574b3f",x"574c40",x"53483d",x"4e4338",x"4d4137",x"463c32",x"463b31",x"45392f",x"473c31",x"493d32",x"4a3d33",x"463a2f",x"4a3f35",x"4b3f34",x"4d4136",x"4f4338",x"4f4338",x"4b3e33",x"4c3f34",x"4d4136",x"4d4034",x"4a3e33",x"4a3e34",x"4a3f34",x"514439",x"574a3e",x"55483c",x"54473b",x"56493d",x"53463b",x"4e4237",x"4d4035",x"4b3e32",x"493d32",x"4d4136",x"4f4439",x"52463a",x"514539",x"54483d",x"524539",x"55493d",x"574a3e",x"54483c",x"574b3f",x"594d41",x"584c3f",x"5c4f43",x"5c5044",x"5d5145",x"5b4f43",x"5c5044",x"5c4f43",x"54473b",x"5a4e42",x"5b4f44",x"594c3f",x"584b3e",x"524538",x"4f4135",x"514336",x"4d4034",x"4e4034",x"514539",x"55493d",x"584c40",x"584d42",x"554a3f",x"4f4339",x"51463c",x"54473b",x"56483c",x"56483c",x"604e3d",x"000000",x"2d1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a140d",x"271e16",x"241d17",x"251f18",x"231c16",x"1f1912",x"1b150d",x"161009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a140d",x"3a2b1e",x"211b14",x"221c15",x"211b14",x"1f1811",x"19130c",x"160f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17100a",x"18120b",x"19130c",x"1b140e",x"1b140e",x"1b140e",x"1b150e",x"1d1710",x"1d1710",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1a0f",x"2a1a0f",x"412411",x"452813",x"472914",x"472913",x"482812",x"482711",x"472711",x"492811",x"472711",x"482711",x"4b2a13",x"452611",x"472811",x"492912",x"472811",x"472712",x"422410",x"452611",x"472812",x"442611",x"432510",x"462711",x"452711",x"4a2a13",x"4f2d15",x"492913",x"4a2a14",x"4a2913",x"492913",x"492a13",x"472712",x"452712",x"4a2a13",x"462712",x"422511",x"452611",x"482812",x"452610",x"442610",x"452610",x"482913",x"4b2a13",x"472811",x"482811",x"452610",x"472812",x"472813",x"4f2e15",x"4d2c14",x"462711",x"452610",x"452611",x"3f230e",x"482812",x"4a2912",x"482812",x"432611",x"492913",x"4d2c14",x"4d2c14",x"4c2b14",x"4a2a13",x"492913",x"4e2b14",x"4b2a13",x"462812",x"4a2911",x"4b2a12",x"4a2912",x"4b2912",x"4a2911",x"492811",x"4a2912",x"4b2b14",x"4a2913",x"472811",x"472812",x"4b2a13",x"4c2a14",x"4b2b14",x"452711",x"4a2a13",x"442611",x"482813",x"4a2a13",x"482812",x"482812",x"4c2a13",x"4a2912",x"4e2b14",x"4e2c15",x"502c14",x"4e2c14",x"462611",x"472712",x"462711",x"502e15",x"4b2913",x"492812",x"4a2912",x"4a2912",x"43240f",x"442510",x"482711",x"4b2912",x"482811",x"432410",x"4d2a12",x"4a2912",x"4b2912",x"482812",x"462611",x"492811",x"492812",x"4c2a12",x"4a2913",x"4d2b13",x"462610",x"462611",x"482712",x"4a2912",x"492812",x"4b2a13",x"4e2c14",x"512d15",x"492912",x"4a2912",x"482812",x"452611",x"4b2b13",x"4b2b14",x"4a2a13",x"4e2c14",x"4f2d15",x"522f16",x"4f2d14",x"4d2b13",x"4c2a13",x"4d2b13",x"4e2c14",x"4c2a14",x"4d2b14",x"4d2b14",x"4f2c13",x"4f2d14",x"482812",x"462610",x"452611",x"492912",x"472812",x"472711",x"4a2a13",x"492913",x"492a13",x"4c2b14",x"482812",x"432511",x"452611",x"452611",x"4c2b13",x"4d2c14",x"492913",x"512e15",x"492913",x"492812",x"4c2b14",x"4c2b14",x"4a2a13",x"492912",x"4a2813",x"4a2912",x"4b2912",x"4a2912",x"4c2b13",x"4a2a12",x"4d2b13",x"4f2d14",x"4b2c13",x"4b2c13",x"000000"),
(x"685646",x"685646",x"5c4e41",x"5e5043",x"564a3d",x"54483e",x"554a3f",x"584c40",x"574b40",x"584c41",x"574b3f",x"574c40",x"53483d",x"4e4338",x"4d4137",x"463c32",x"463b31",x"45392f",x"473c31",x"493d32",x"4a3d33",x"463a2f",x"4a3f35",x"4b3f34",x"4d4136",x"4f4338",x"4f4338",x"4b3e33",x"4c3f34",x"4d4136",x"4d4034",x"4a3e33",x"4a3e34",x"4a3f34",x"514439",x"574a3e",x"55483c",x"54473b",x"56493d",x"53463b",x"4e4237",x"4d4035",x"4b3e32",x"493d32",x"4d4136",x"4f4439",x"52463a",x"514539",x"54483d",x"524539",x"55493d",x"574a3e",x"54483c",x"574b3f",x"594d41",x"584c3f",x"5c4f43",x"5c5044",x"5d5145",x"5b4f43",x"5c5044",x"5c4f43",x"54473b",x"5a4e42",x"5b4f44",x"594c3f",x"584b3e",x"524538",x"4f4135",x"514336",x"4d4034",x"4e4034",x"514539",x"55493d",x"584c40",x"584d42",x"554a3f",x"4f4339",x"51463c",x"54473b",x"56483c",x"56483c",x"604e3d",x"604e3d",x"2d1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a140d",x"271e16",x"241d17",x"251f18",x"231c16",x"1f1912",x"1b150d",x"161009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a140d",x"3a2b1e",x"211b14",x"221c15",x"211b14",x"1f1811",x"19130c",x"160f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17100a",x"18120b",x"19130c",x"1b140e",x"1b140e",x"1b140e",x"1b150e",x"1d1710",x"1d1710",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1a0f",x"2a1a0f",x"412411",x"452813",x"472914",x"472913",x"482812",x"482711",x"472711",x"492811",x"472711",x"482711",x"4b2a13",x"452611",x"472811",x"492912",x"472811",x"472712",x"422410",x"452611",x"472812",x"442611",x"432510",x"462711",x"452711",x"4a2a13",x"4f2d15",x"492913",x"4a2a14",x"4a2913",x"492913",x"492a13",x"472712",x"452712",x"4a2a13",x"462712",x"422511",x"452611",x"482812",x"452610",x"442610",x"452610",x"482913",x"4b2a13",x"472811",x"482811",x"452610",x"472812",x"472813",x"4f2e15",x"4d2c14",x"462711",x"452610",x"452611",x"3f230e",x"482812",x"4a2912",x"482812",x"432611",x"492913",x"4d2c14",x"4d2c14",x"4c2b14",x"4a2a13",x"492913",x"4e2b14",x"4b2a13",x"462812",x"4a2911",x"4b2a12",x"4a2912",x"4b2912",x"4a2911",x"492811",x"4a2912",x"4b2b14",x"4a2913",x"472811",x"472812",x"4b2a13",x"4c2a14",x"4b2b14",x"452711",x"4a2a13",x"442611",x"482813",x"4a2a13",x"482812",x"482812",x"4c2a13",x"4a2912",x"4e2b14",x"4e2c15",x"502c14",x"4e2c14",x"462611",x"472712",x"462711",x"502e15",x"4b2913",x"492812",x"4a2912",x"4a2912",x"43240f",x"442510",x"482711",x"4b2912",x"482811",x"432410",x"4d2a12",x"4a2912",x"4b2912",x"482812",x"462611",x"492811",x"492812",x"4c2a12",x"4a2913",x"4d2b13",x"462610",x"462611",x"482712",x"4a2912",x"492812",x"4b2a13",x"4e2c14",x"512d15",x"492912",x"4a2912",x"482812",x"452611",x"4b2b13",x"4b2b14",x"4a2a13",x"4e2c14",x"4f2d15",x"522f16",x"4f2d14",x"4d2b13",x"4c2a13",x"4d2b13",x"4e2c14",x"4c2a14",x"4d2b14",x"4d2b14",x"4f2c13",x"4f2d14",x"482812",x"462610",x"452611",x"492912",x"472812",x"472711",x"4a2a13",x"492913",x"492a13",x"4c2b14",x"482812",x"432511",x"452611",x"452611",x"4c2b13",x"4d2c14",x"492913",x"512e15",x"492913",x"492812",x"4c2b14",x"4c2b14",x"4a2a13",x"492912",x"4a2813",x"4a2912",x"4b2912",x"4a2912",x"4c2b13",x"4a2a12",x"4d2b13",x"4f2d14",x"4b2c13",x"4b2c13",x"000000"),
(x"685645",x"685645",x"544638",x"584b3f",x"56483c",x"57493d",x"5c4e41",x"5d4e40",x"5b4c3e",x"605144",x"5e4f40",x"5f5144",x"5d4d40",x"564638",x"574739",x"534335",x"4e3e31",x"514134",x"544334",x"574637",x"584838",x"564639",x"584738",x"564535",x"574638",x"594739",x"554537",x"574637",x"554434",x"5c4a3a",x"524335",x"584636",x"4e3e31",x"534335",x"594739",x"58493b",x"5c4d3f",x"5e4e40",x"5f4f40",x"5e4e3f",x"5c4c3d",x"594838",x"594737",x"5a493a",x"5a493a",x"5b493a",x"5e4c3c",x"5f4e3f",x"5a493a",x"5c4a3a",x"5e4e3f",x"604f40",x"615142",x"605143",x"605143",x"5b4c3d",x"615245",x"635244",x"5f5042",x"615143",x"5a4a3c",x"635345",x"605144",x"625142",x"5b4d40",x"625141",x"5d4d3e",x"59483a",x"574738",x"584739",x"564435",x"544333",x"574638",x"584739",x"5c4d40",x"5a4b3d",x"5a4b3e",x"5b4c3e",x"57483a",x"57483b",x"58493b",x"5a4b3d",x"5b4b3d",x"5b4b3d",x"2d1a0b",x"4a3421",x"332316",x"2f2114",x"332416",x"2f2114",x"2d1f13",x"241b12",x"513c29",x"3d2e21",x"35281c",x"35281d",x"2f2217",x"2e2115",x"322216",x"2f2114",x"2e2013",x"2d1f13",x"2b1e12",x"2f2114",x"302215",x"312316",x"302215",x"312215",x"2b1e12",x"2d2013",x"302215",x"2d2013",x"281c10",x"2e2013",x"2e2013",x"332417",x"2c1e12",x"2d1f12",x"2d1f12",x"2d1f13",x"291c11",x"2b1e12",x"271b10",x"25190e",x"25190e",x"291c11",x"261a0e",x"25190e",x"24190e",x"21170c",x"281b10",x"21160c",x"21170c",x"21160c",x"24190e",x"20160d",x"21170d",x"20160d",x"21170d",x"20160c",x"21160d",x"21160d",x"23190f",x"1b140d",x"4a3524",x"443324",x"3f2f21",x"413123",x"3f2f20",x"3b2b1c",x"342516",x"352517",x"372718",x"362617",x"302114",x"382718",x"372718",x"39281a",x"302113",x"322315",x"2c1e11",x"312213",x"332416",x"302214",x"312214",x"312214",x"322215",x"332416",x"332417",x"312316",x"322416",x"2d1f13",x"2e2013",x"2d2013",x"2e2014",x"291d11",x"2a1d11",x"281c10",x"2a1d11",x"271b10",x"23180e",x"20160c",x"23180d",x"23180e",x"20160c",x"21160d",x"20150c",x"25190e",x"20160c",x"1e140b",x"1d130a",x"1d140b",x"1c120a",x"1e150d",x"20180f",x"1c140d",x"1d160f",x"1e160f",x"201811",x"241b13",x"201811",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150d",x"1c150d",x"1f150d",x"22160e",x"20140c",x"27180e",x"2e1b0e",x"311c0d",x"301b0c",x"321c0c",x"311c0c",x"351d0d",x"361e0d",x"351d0d",x"341c0c",x"311b0b",x"331c0c",x"331c0c",x"2e190b",x"2d190a",x"2e1a0b",x"2f1a0b",x"2c180a",x"2c180a",x"39200f",x"3d2310",x"3b2210",x"3d2210",x"39200e",x"351c0c",x"381f0d",x"3e230f",x"432713",x"3c220f",x"3f2411",x"3d220f",x"3c210f",x"3b2210",x"3f2512",x"442813",x"412612",x"422612",x"402511",x"3a210f",x"3b210f",x"381f0e",x"3e2310",x"381f0e",x"361f0e",x"331c0d",x"38200e",x"3a210f",x"422611",x"3e2310",x"412511",x"3a210f",x"3e2310",x"3d2310",x"3c2310",x"432712",x"422713",x"402612",x"3d2411",x"3d2310",x"3f2411",x"402612",x"402511",x"3f2410",x"3b210f",x"3b210e",x"3a200e",x"3d220f",x"3a210f",x"3c210f",x"3c210f",x"3b210f",x"371f0e",x"381f0e",x"39200f",x"351e0e",x"29170a",x"371f0d",x"402410",x"150e07",x"150e07",x"221409",x"231409",x"2c190b",x"351e0e",x"361e0e",x"351e0d",x"39200e",x"361e0e",x"361e0d",x"371f0e",x"361f0d",x"351e0d",x"331c0d",x"331d0d",x"39200f",x"38200e",x"39200e",x"39200e",x"371e0d",x"341c0c",x"271307",x"261207",x"2a1509",x"301a0b",x"311b0b",x"331c0c",x"341d0c",x"331c0c",x"341d0d",x"361e0d",x"3a210f",x"391f0d",x"381e0d",x"3b200e",x"351d0d",x"391f0e",x"351d0c",x"351d0c",x"381e0d",x"351d0c",x"331b0b",x"39200e",x"371f0e",x"3a210f",x"38200f",x"361e0d",x"2e190b",x"2f1a0b",x"361e0d",x"371f0e",x"3e2310",x"3d2310",x"412511",x"3b200e",x"3b210f",x"3f2511",x"3d2411",x"3b2210",x"3b2210",x"3e2411",x"3f2410",x"3c220f",x"391f0e",x"3c210f",x"3d220f",x"3c210f",x"391f0e",x"381f0e",x"3b210f",x"38200f",x"3d2310",x"3c220f",x"3a2210",x"3b2210",x"3b2210",x"3c2310",x"3f2511",x"3f2512",x"412712",x"402612",x"3d2310",x"402411",x"382110",x"392110",x"3f2410",x"3d2310",x"361f0e",x"40250f",x"3d230e",x"432710",x"41260f",x"422710",x"442810",x"4b2c12",x"442811",x"442811",x"000000"),
(x"6d5846",x"6d5846",x"594b3f",x"4f4337",x"55473a",x"57483c",x"594b3f",x"58483b",x"57483a",x"57483b",x"57493c",x"584a3d",x"4f4033",x"4e4033",x"4b3d31",x"4c3d31",x"4e3f32",x"4b3c2f",x"4b3d30",x"514234",x"544436",x"564436",x"4f3f31",x"4f3f31",x"534133",x"514133",x"4f3f30",x"514031",x"4f3e2f",x"4f3e30",x"4b3b2d",x"4c3d2f",x"4e3e2f",x"524233",x"4f3f32",x"554538",x"5a4a3b",x"5b4b3d",x"5c4a3b",x"5e4d3e",x"5a4839",x"574535",x"4f3e2f",x"554333",x"514032",x"554435",x"554537",x"544335",x"554435",x"564435",x"574637",x"564535",x"574738",x"554537",x"514235",x"574739",x"574739",x"554538",x"554538",x"544537",x"564638",x"564739",x"514234",x"554538",x"574738",x"504030",x"534233",x"4e3f31",x"4d3c2d",x"503f30",x"504032",x"503d2e",x"534131",x"513f2f",x"504133",x"504033",x"4d3f32",x"4b3d31",x"4c3f32",x"4d3f33",x"514336",x"554538",x"58483a",x"58483a",x"221409",x"4c3522",x"2f2114",x"2f2114",x"332416",x"2f2114",x"2e2015",x"1d1710",x"543d2a",x"3d2d21",x"33281d",x"32271c",x"302419",x"2a1e14",x"2d1f14",x"2b1d11",x"2f2013",x"322315",x"342416",x"342416",x"2d2013",x"2c1f12",x"291c10",x"2c1f12",x"322215",x"2c1e12",x"2d1f13",x"2e2013",x"2d1f13",x"2c1e12",x"2d1f12",x"2f2114",x"2d2013",x"2e2013",x"281c10",x"281c10",x"2d1f13",x"261a0f",x"261a0f",x"271a0f",x"281b10",x"2a1d11",x"25190e",x"271b0f",x"261a0e",x"20160c",x"25190f",x"1f150b",x"22170d",x"25190e",x"20160c",x"23180d",x"23180e",x"23180d",x"1f150b",x"20160c",x"20150c",x"1f150b",x"241910",x"1d1610",x"493626",x"403022",x"3c2d21",x"3f2f21",x"3e2e21",x"3b2b1d",x"362617",x"342416",x"372718",x"302214",x"302114",x"342416",x"362517",x"362617",x"2c1e11",x"2f2012",x"342415",x"2f2013",x"342416",x"302214",x"342416",x"312214",x"342416",x"322316",x"2d2013",x"312215",x"2b1e11",x"2e2013",x"2c1e12",x"2b1e11",x"2b1d11",x"2c1e12",x"2b1e12",x"281b10",x"271b10",x"291d11",x"251a0f",x"20160c",x"1f150b",x"21170d",x"22170d",x"261a0f",x"23180d",x"1d130a",x"20160c",x"1d140b",x"1e140b",x"1f150b",x"1c130a",x"1e150c",x"20170f",x"1e160f",x"221910",x"201811",x"231b13",x"241c14",x"211912",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211810",x"211810",x"1d1610",x"281a10",x"332012",x"332011",x"382212",x"3b2312",x"3c2411",x"3c2411",x"3c2311",x"3d2411",x"3d2411",x"3f2512",x"442914",x"432814",x"3e2411",x"3e2411",x"402612",x"3b2311",x"311d0d",x"38210f",x"361f0f",x"301c0c",x"2f1b0c",x"3a2210",x"3d2310",x"3c2210",x"472b15",x"492c15",x"4a2c15",x"402511",x"3c2311",x"402612",x"412712",x"442813",x"3e2310",x"3e220f",x"402410",x"432712",x"422712",x"412612",x"3e2310",x"3c220f",x"3d2310",x"3b220f",x"3b2210",x"3b2210",x"361f0e",x"3d2411",x"3d2410",x"381f0e",x"3f2411",x"3f2511",x"432713",x"3c220f",x"3c220f",x"39200f",x"39210f",x"3a2210",x"351f0f",x"3e2411",x"3d2411",x"3a2210",x"3c2310",x"3b2210",x"3b2310",x"3f2410",x"3c220f",x"3c2210",x"3c2210",x"3b210f",x"3c210f",x"402612",x"3d2310",x"3e2411",x"3e2311",x"3d2411",x"3e2511",x"38210f",x"25150a",x"3b210f",x"3e220f",x"150e07",x"150e07",x"150e07",x"29170b",x"2e1a0c",x"321c0d",x"341e0d",x"321c0c",x"311b0c",x"3a200e",x"341d0c",x"371f0d",x"3a210f",x"38200e",x"39200f",x"351e0e",x"3a200f",x"3b220f",x"3c2310",x"3e2411",x"412712",x"3f2512",x"3e2411",x"3c2310",x"3b2311",x"422712",x"3e2511",x"3c2411",x"422713",x"3f2512",x"402512",x"412713",x"432713",x"432814",x"492c16",x"462a14",x"452813",x"432813",x"462a14",x"422713",x"412612",x"452914",x"3f2410",x"3f2411",x"3e2310",x"3e2411",x"39200f",x"3c2311",x"402612",x"412612",x"412612",x"3e2411",x"402512",x"412712",x"412712",x"3d2310",x"381f0e",x"381f0e",x"39210f",x"3e2411",x"3c2310",x"3b220f",x"3b210f",x"3e2410",x"3c220f",x"3a210f",x"3b2210",x"3e2411",x"3a210f",x"3a220f",x"3f2411",x"3c2310",x"361f0e",x"402612",x"3c2210",x"3b210f",x"3a210f",x"3a210f",x"3b2210",x"3d2411",x"3c2311",x"402512",x"412612",x"412612",x"3e2310",x"402511",x"3e2411",x"3e230f",x"3c230f",x"402510",x"412610",x"412610",x"432910",x"492c12",x"472b11",x"4b2e13",x"452911",x"452911",x"000000"),
(x"705946",x"705946",x"524437",x"544639",x"514336",x"56473a",x"544639",x"534538",x"544538",x"534336",x"4d3e31",x"514234",x"4f4034",x"4a3c2f",x"483a2d",x"47392d",x"48392d",x"46382c",x"503f30",x"544334",x"544335",x"534233",x"514031",x"524032",x"554332",x"544131",x"524031",x"523f30",x"534031",x"4f3d2e",x"544233",x"503e30",x"513e2f",x"544131",x"544233",x"554335",x"554436",x"5a4939",x"5f4e3f",x"594839",x"544435",x"544233",x"503f30",x"534131",x"4e3d2e",x"4e3b2d",x"4e3d2d",x"503e2f",x"503e2d",x"49392b",x"4b3a2b",x"4f3d2e",x"4d3d2e",x"503e2f",x"503e2f",x"4e3e30",x"504031",x"4f3e2f",x"503e2e",x"503e30",x"503f30",x"4f3e30",x"524031",x"4f3e31",x"544233",x"534131",x"513f2f",x"513e2d",x"55402e",x"564230",x"503d2b",x"4f3c2d",x"4a3a2b",x"523f2f",x"503d2d",x"4b3a2d",x"4a3b2d",x"49382c",x"47382b",x"493c2f",x"4e3f32",x"4d4035",x"58483a",x"58483a",x"1e1209",x"4f3925",x"342416",x"342416",x"342516",x"332416",x"362617",x"1b140e",x"563f2b",x"3d2d20",x"3d2e22",x"30251a",x"35271a",x"332418",x"2a1d11",x"312215",x"302114",x"332416",x"352517",x"332416",x"2d2013",x"2c1e12",x"2a1d11",x"291c10",x"2d2013",x"2d1f13",x"271a0f",x"2b1e11",x"2a1d11",x"2d1f13",x"2e2013",x"2e1f13",x"2e2013",x"2e2014",x"281c10",x"2a1d11",x"2c1f12",x"2d1f13",x"291d11",x"281b10",x"281c10",x"291c10",x"2d2014",x"261a0f",x"281c10",x"251a0f",x"23180d",x"251a0f",x"22170d",x"24190e",x"21170d",x"20160c",x"23180e",x"23170d",x"20160c",x"1f150b",x"1f150b",x"1f150b",x"20170f",x"1d1710",x"493626",x"402f21",x"3e2f22",x"3e2e21",x"3f2f20",x"392a1b",x"362618",x"382718",x"382718",x"372718",x"3a291a",x"352517",x"382718",x"362517",x"362618",x"312214",x"362617",x"372718",x"362617",x"392818",x"322215",x"362618",x"342517",x"332416",x"322315",x"342416",x"312215",x"2c1e12",x"2d2013",x"2d1f13",x"2a1d11",x"291d11",x"291c10",x"291c11",x"261a0f",x"25190e",x"251a0f",x"291c11",x"23180d",x"23180d",x"23180d",x"23180e",x"21160d",x"20150c",x"23180d",x"1f150b",x"22170d",x"1c130a",x"1b130b",x"1c150d",x"20180f",x"221911",x"231a11",x"251c14",x"261d15",x"221a13",x"231b13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231911",x"231911",x"1d160f",x"271a11",x"2d1c11",x"321f12",x"372112",x"2a1a0d",x"3c2311",x"38210f",x"3a2110",x"3d2411",x"3b2310",x"3d2411",x"3e2411",x"3d2311",x"3c230f",x"3a2210",x"38200f",x"351e0d",x"361f0e",x"351f0e",x"3c2311",x"392110",x"361f0e",x"361f0e",x"3f2512",x"412613",x"422712",x"422713",x"3a2210",x"361f0e",x"39210f",x"3f2511",x"3f2511",x"3f2310",x"3d2310",x"3c210f",x"3e220f",x"3f2411",x"3d2310",x"3b210f",x"3b210f",x"3b210f",x"3a210f",x"3e2310",x"3e2311",x"3f2511",x"422712",x"422712",x"402612",x"432813",x"422713",x"402612",x"3e2411",x"3e2411",x"402511",x"3f2411",x"402511",x"3e2411",x"3b2210",x"3b210f",x"38200e",x"37200e",x"381f0e",x"361e0d",x"361f0d",x"3b210f",x"361f0e",x"351e0e",x"3d2310",x"3e2311",x"3d2310",x"3d2412",x"3d2412",x"372010",x"39210f",x"3a210f",x"39210f",x"321c0c",x"3b210f",x"3a200e",x"3f2410",x"3e230f",x"160e07",x"150e07",x"211309",x"28160a",x"2d190b",x"2f1a0b",x"301b0b",x"321c0c",x"311a0b",x"2e180a",x"2b170a",x"2e180a",x"2e190a",x"311b0b",x"341d0c",x"371f0e",x"39200e",x"361f0e",x"38200e",x"361e0e",x"371f0e",x"3a210f",x"321c0d",x"3c2210",x"38210f",x"3c2311",x"3e2411",x"432813",x"3e2411",x"402512",x"402612",x"412713",x"422712",x"412612",x"3f2411",x"412511",x"422612",x"3d220f",x"3f2410",x"432712",x"442813",x"452914",x"3d2310",x"3d2310",x"3e2411",x"412613",x"402612",x"3f2512",x"3e2511",x"3a210f",x"3b210f",x"3a2310",x"3d2410",x"3a210f",x"38200e",x"38200e",x"351d0d",x"361f0e",x"39200f",x"3a210f",x"3c220f",x"3b220f",x"3b220f",x"3e2410",x"3e2411",x"3d2310",x"422712",x"452914",x"412612",x"3f2512",x"412612",x"432813",x"3f2511",x"412612",x"38210f",x"39210f",x"3d2310",x"3f2411",x"3d2310",x"3a2110",x"3a210f",x"3c220f",x"3d220f",x"371f0e",x"38200d",x"3e230f",x"3f240f",x"402510",x"41260f",x"452a11",x"452a11",x"462a10",x"492b11",x"492c11",x"4c2e13",x"462911",x"462911",x"000000"),
(x"6b5542",x"6b5542",x"4d4035",x"4f4236",x"4b3e32",x"504235",x"524335",x"4f4032",x"514234",x"4e3f32",x"4e3f31",x"4c3e32",x"504032",x"4f4031",x"4f3f31",x"4e3d2f",x"4d3f31",x"4c3c2e",x"503f31",x"514133",x"4c3d2f",x"504031",x"4f3e2f",x"513f30",x"544131",x"523f2f",x"524030",x"554130",x"554131",x"5a4634",x"4e3c2d",x"523f2f",x"503e2e",x"4e3d2e",x"4c3b2b",x"544232",x"544334",x"574535",x"5a4838",x"5a4839",x"5a4838",x"514031",x"514130",x"534232",x"544132",x"584331",x"4f3d2d",x"4f3e2e",x"53402f",x"523f2f",x"4f3c2d",x"4f3c2d",x"4d3c2d",x"4d3b2c",x"514031",x"513e2e",x"4a3a2c",x"4a392b",x"4e3c2d",x"544132",x"524030",x"544232",x"4f3d2d",x"4f3e2f",x"543f2d",x"513d2b",x"503c2b",x"533f2e",x"503d2c",x"4d3c2b",x"523e2c",x"4f3d2c",x"503e2e",x"4c3b2c",x"503e2d",x"523f2e",x"4c3b2b",x"49382b",x"493a2c",x"4b3a2c",x"4e4032",x"514234",x"58483a",x"58483a",x"150e07",x"4a3421",x"392819",x"372718",x"342416",x"382718",x"342416",x"171009",x"5d442f",x"443223",x"33261a",x"2f2218",x"2e2014",x"2f2115",x"2b1d11",x"2d1f12",x"2a1d11",x"312215",x"312316",x"332416",x"2e2114",x"2b1f13",x"2b1f13",x"312316",x"352518",x"2e2014",x"2f2114",x"2e2013",x"302214",x"2f2114",x"2c1e12",x"2f2014",x"2c1f12",x"2a1d11",x"2b1e12",x"2d1f13",x"2d1f12",x"2e2013",x"261a0f",x"2c1e12",x"2c1f13",x"271b10",x"281c10",x"291c10",x"271b10",x"271a0f",x"23180d",x"22170d",x"261a0f",x"271b10",x"291c11",x"21170d",x"21170d",x"1d140b",x"24190e",x"20160d",x"21170d",x"21170d",x"21180e",x"1d1710",x"503b29",x"453424",x"403123",x"403023",x"3c2c1f",x"38281b",x"3e2c1c",x"372718",x"3a2919",x"3b2919",x"3b2a1a",x"382819",x"3a2a1a",x"3c2a1b",x"382818",x"342516",x"352517",x"2e2013",x"342415",x"352517",x"312214",x"352517",x"352517",x"39291a",x"332517",x"302316",x"302215",x"322517",x"302215",x"2e2114",x"2f2114",x"302214",x"2c1f12",x"2b1e12",x"281b10",x"271b0f",x"24180e",x"281c10",x"251a0f",x"20160c",x"20160c",x"23180d",x"23180e",x"24180e",x"21170d",x"21170d",x"20160c",x"1d140b",x"1f160d",x"20170e",x"241a11",x"231a12",x"231a12",x"251c14",x"211912",x"261e15",x"221b14",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"241a12",x"241a12",x"1e1711",x"1e1711",x"291b10",x"2d1c11",x"311e10",x"2d1b0d",x"311c0c",x"351e0e",x"39200f",x"331d0d",x"39200f",x"37200e",x"351e0d",x"371e0d",x"341d0d",x"321c0c",x"331c0c",x"351d0d",x"331c0d",x"331c0c",x"2e190b",x"2d190b",x"2f1a0b",x"2e190b",x"351d0d",x"311a0b",x"321b0b",x"371e0d",x"361f0e",x"361f0e",x"321c0c",x"351d0d",x"3e2311",x"402511",x"402512",x"402612",x"462914",x"432813",x"422612",x"3d2210",x"391f0e",x"371e0d",x"381f0e",x"381f0e",x"391f0e",x"361d0d",x"311b0c",x"3a210f",x"39210f",x"3f2411",x"3b2311",x"422713",x"412713",x"412613",x"402512",x"3e2512",x"462914",x"422713",x"412713",x"422813",x"412713",x"321d0e",x"3b210f",x"3f2511",x"412612",x"3e2410",x"442813",x"452a14",x"462914",x"472a14",x"412612",x"442814",x"412713",x"3b2211",x"3c2311",x"39200e",x"3a210f",x"361f0e",x"3f2410",x"3d230f",x"3f2410",x"3e220f",x"381f0e",x"160e07",x"241509",x"231409",x"29170a",x"2e1a0b",x"321b0c",x"321c0c",x"331c0c",x"341d0c",x"341d0c",x"311b0c",x"341c0c",x"361e0d",x"351e0d",x"371e0d",x"351e0d",x"361e0d",x"371f0e",x"361e0d",x"341d0d",x"39200f",x"39200f",x"361f0e",x"39200f",x"371f0e",x"371f0e",x"3b210f",x"3a210f",x"3a210f",x"3d2310",x"3e2310",x"39200e",x"391f0e",x"3a200e",x"39200d",x"351d0c",x"361e0d",x"3c220f",x"391f0e",x"371e0d",x"331b0b",x"341d0c",x"361e0d",x"341c0c",x"341c0c",x"341c0b",x"321b0c",x"361f0e",x"38200f",x"38200e",x"331c0c",x"39200f",x"3d2310",x"39200f",x"3f2512",x"3e2511",x"3b2311",x"3c2311",x"3b2210",x"3a200e",x"351d0d",x"381f0d",x"3b200f",x"351d0d",x"361d0d",x"361d0d",x"381f0e",x"3f2412",x"3f2512",x"3e2512",x"432813",x"442813",x"382110",x"402612",x"452914",x"412612",x"402512",x"402612",x"432814",x"432814",x"412612",x"3f230f",x"3b220f",x"462912",x"442811",x"452912",x"4a2d15",x"4b2e15",x"4b2d14",x"4a2c13",x"4a2d12",x"4b2e13",x"462a11",x"4a2c11",x"442811",x"442811",x"000000"),
(x"6e5743",x"6e5743",x"4d3f31",x"493b2f",x"493b2d",x"4a3c2f",x"4e3e30",x"4f3f32",x"514132",x"4e3e2f",x"4a3b2e",x"4d3d30",x"4e3e2f",x"4d3e2f",x"4a392b",x"513f31",x"4d3c2e",x"503f2f",x"524031",x"514030",x"4d3c2e",x"4f3d2f",x"4e3c2e",x"534030",x"4f3c2d",x"503e2e",x"523f2e",x"4e3c2d",x"544131",x"55402f",x"513c2b",x"54402e",x"564230",x"564130",x"584331",x"56412d",x"584332",x"574333",x"594534",x"5e4936",x"5b4735",x"564231",x"58422f",x"574330",x"544130",x"534130",x"53402f",x"513e2d",x"564131",x"513f2e",x"523e2e",x"4f3d2d",x"513e2e",x"503d2d",x"4e3c2b",x"4f3c2d",x"503d2d",x"4c3b2b",x"4e3c2d",x"4f3c2d",x"513f2f",x"4f3d2e",x"4f3c2d",x"4f3e2c",x"594430",x"55402e",x"533f2e",x"543f2c",x"503d2c",x"4d3b2c",x"513e2d",x"513f2d",x"4e3b2b",x"533f2d",x"4f3d2d",x"4f3c2a",x"523f2d",x"4b392b",x"483a2c",x"4a3b2d",x"4a3d31",x"534437",x"5b4a3b",x"5b4a3b",x"150e07",x"4e3723",x"392819",x"362618",x"372618",x"392819",x"352517",x"171009",x"5f462f",x"3d2c1c",x"342518",x"352618",x"2f2114",x"302114",x"2d1f12",x"2d1f12",x"332315",x"2b1d11",x"322316",x"312316",x"322416",x"312215",x"332417",x"302215",x"322315",x"312215",x"2d2013",x"312214",x"2f2114",x"312215",x"322315",x"302114",x"2d1f12",x"2d1f12",x"2d1f12",x"2c1f12",x"291c10",x"2d1f13",x"2b1e12",x"2a1d11",x"2c1f13",x"23180d",x"281c10",x"291c10",x"2b1e12",x"261a0f",x"291c10",x"251a0e",x"25190e",x"25190f",x"2c1e12",x"241a0f",x"251a0f",x"21170d",x"24190f",x"21170d",x"21160c",x"20160c",x"23180f",x"1d160f",x"4e3a29",x"463424",x"423123",x"433223",x"3d2d1f",x"3d2c1d",x"382718",x"3b291a",x"382818",x"392819",x"382718",x"352517",x"392819",x"392818",x"3d2a1b",x"382818",x"352517",x"362617",x"372617",x"3a2919",x"362617",x"382718",x"362618",x"352719",x"372719",x"352618",x"2f2114",x"302215",x"342416",x"2e2013",x"322316",x"2e2013",x"2f2114",x"281c10",x"2d1f13",x"2a1d11",x"271b10",x"271b10",x"24190e",x"23180d",x"251a0f",x"23180e",x"21160d",x"20150c",x"24190e",x"21160c",x"23180d",x"1d140b",x"22170e",x"221910",x"221a11",x"201810",x"221a13",x"251c14",x"261d15",x"231c15",x"251d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"251c14",x"251c14",x"201912",x"1f1811",x"241910",x"291b11",x"321e11",x"3b2110",x"371f0d",x"3e230f",x"422510",x"412410",x"402410",x"3b200e",x"3d220f",x"432611",x"3b200e",x"3a200d",x"3a1f0d",x"3c210e",x"412410",x"422511",x"3e220f",x"3d220f",x"402410",x"3a200e",x"3d220f",x"3c210e",x"442611",x"452711",x"452812",x"462812",x"492a13",x"4c2c15",x"4b2b14",x"452611",x"3f230f",x"462712",x"4c2c14",x"482812",x"482913",x"4c2c14",x"482913",x"462611",x"432410",x"41230f",x"3a1f0d",x"3c200d",x"412310",x"472913",x"422611",x"472914",x"472912",x"472812",x"482a13",x"472913",x"4c2c15",x"4d2d15",x"4c2d15",x"4a2b14",x"4a2b14",x"482914",x"482a14",x"492b15",x"4a2b14",x"4a2a14",x"502f17",x"4b2c16",x"472913",x"472913",x"4e2e16",x"4b2b14",x"4f2f17",x"56341a",x"4f3018",x"54341a",x"482b15",x"442915",x"3c2311",x"341f0f",x"371e0d",x"361e0d",x"371f0e",x"402511",x"432712",x"180f07",x"160e07",x"24150a",x"3d2410",x"432712",x"432711",x"402410",x"432611",x"432611",x"472812",x"452712",x"472812",x"462712",x"472912",x"452712",x"462813",x"472912",x"452711",x"432611",x"432611",x"442611",x"452611",x"412310",x"3e220e",x"3c210e",x"412410",x"3f230f",x"412410",x"422510",x"40230f",x"3f220f",x"41240f",x"442611",x"432511",x"3e210e",x"42240f",x"41240f",x"452611",x"432611",x"482913",x"432511",x"442611",x"462711",x"422410",x"40230f",x"452711",x"452711",x"482a13",x"452712",x"4a2a14",x"482a14",x"462813",x"462712",x"442510",x"442611",x"492a13",x"482913",x"442611",x"482913",x"432611",x"442611",x"402310",x"3f220f",x"3f220e",x"3b200d",x"3d210e",x"482915",x"4a2b15",x"4a2b15",x"472913",x"311c0d",x"3c220f",x"3c2310",x"3c2310",x"3b2210",x"3b2210",x"3a2110",x"3a2210",x"3b2210",x"3a2110",x"412612",x"4a2b15",x"4a2a13",x"462912",x"4d2f15",x"4b2c15",x"4d2e15",x"4d2d14",x"4d2e14",x"4d2e13",x"4c2e14",x"513115",x"543416",x"533317",x"4f3016",x"51311d",x"51311d"),
(x"6b5440",x"6b5440",x"493b2e",x"46392c",x"473a2e",x"493b2f",x"46382b",x"4e3e30",x"4d3c2f",x"4d3d2f",x"4b3c2f",x"483a2d",x"534133",x"4d3c2d",x"524133",x"554334",x"4d3e31",x"4c3c2e",x"4b3a2c",x"503f2f",x"4e3d2d",x"4f3e2f",x"4e3d2d",x"4f3d2d",x"49392a",x"513e2f",x"503e2e",x"553f2e",x"543f2d",x"574130",x"56412f",x"55412f",x"59432f",x"594430",x"56412f",x"513d2c",x"513e2d",x"533f2e",x"564130",x"5b4533",x"594431",x"5c4533",x"5b4531",x"5a4431",x"5d4632",x"55402e",x"584331",x"584330",x"584331",x"57422f",x"533f2e",x"52402e",x"55402f",x"543f2e",x"54402f",x"53402e",x"4f3d2b",x"4d3b2c",x"4b3a2a",x"513d2d",x"4e3c2c",x"503e2e",x"553f2e",x"513d2b",x"4e3b2b",x"533f2c",x"553f2b",x"513e2a",x"4e3b2a",x"4c3929",x"4a3829",x"4c3b2b",x"4f3d2d",x"4c3b2b",x"4f3c2b",x"4c3a2a",x"503e2d",x"523e2c",x"523f2f",x"4c3d2f",x"504133",x"554638",x"5a4a3b",x"5a4a3b",x"150e07",x"493421",x"3b2a1a",x"362617",x"342415",x"342416",x"322315",x"171009",x"61452d",x"3b2a1a",x"312216",x"342417",x"312215",x"312214",x"302114",x"2a1d11",x"281b0f",x"2d1f12",x"2d1f12",x"322316",x"342416",x"312216",x"352518",x"2e2014",x"352618",x"2f2114",x"2f2114",x"352617",x"342518",x"312215",x"312214",x"2f2014",x"312215",x"312215",x"2e2013",x"2d1f12",x"2c1e12",x"271b0f",x"291c10",x"281c10",x"281c10",x"281c10",x"281b10",x"22170d",x"281c10",x"25190e",x"24190e",x"21170c",x"1f150b",x"21160c",x"281b10",x"261a0f",x"261a0f",x"22170d",x"1e150c",x"20160c",x"24190f",x"21160d",x"22180f",x"1b140d",x"4d3a28",x"4b3827",x"3e2f22",x"3f2f22",x"402f21",x"3d2c1d",x"382718",x"3c2a1a",x"3a2819",x"372617",x"322315",x"3a2819",x"382718",x"3c2a1b",x"322215",x"352517",x"372718",x"332416",x"352517",x"312214",x"2c1d11",x"322214",x"332316",x"382718",x"362617",x"362618",x"352518",x"312215",x"312215",x"2d2013",x"332417",x"312215",x"2f2115",x"2d1f12",x"2a1d11",x"251a0f",x"2a1d11",x"23180d",x"25190f",x"24180e",x"24180d",x"22170d",x"22170d",x"23180d",x"23180d",x"20160c",x"20150c",x"1d140b",x"1f160d",x"221911",x"241b13",x"241c14",x"231a12",x"231b14",x"271e16",x"271d15",x"251d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"261d15",x"261d15",x"291c13",x"2d1e15",x"301f14",x"352013",x"2f1b0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17100a",x"171009",x"1a130c",x"19130c",x"19120c",x"462812",x"3b2211",x"371f0e",x"311c0d",x"361f0e",x"402511",x"371f0e",x"3e2310",x"3c2210",x"170f07",x"180f08",x"25160a",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"1c150e",x"1f1811",x"221a13",x"221a12",x"4f2e15",x"3a200f",x"2f1a0b",x"301a0b",x"351d0c",x"341d0c",x"331c0c",x"2e180a",x"321c0c",x"2f1a0b",x"39200f",x"3b220f",x"241409",x"150e07",x"150e07",x"4e3f32",x"41372e",x"150e07",x"1c1108",x"201309",x"382e25",x"3f372f",x"26160a",x"311c0d",x"341d0f",x"3e2310",x"4f3b2d",x"4f3b2d"),
(x"705741",x"705741",x"4e3f32",x"4d3e31",x"48392c",x"4c3d30",x"4f3e2f",x"4d3e30",x"514133",x"4d3d2e",x"534233",x"504032",x"4b3c2f",x"4d3d2f",x"4c3e32",x"4d3e30",x"503f30",x"503e2f",x"4d3c2d",x"523f2f",x"4f3d2e",x"4c3c2d",x"4b3a2b",x"523f2e",x"523f2f",x"503d2d",x"55412f",x"58422f",x"5b4532",x"5d4632",x"5f4733",x"604a34",x"644a34",x"5e4933",x"5a4532",x"5a4431",x"55402d",x"57412f",x"56412f",x"5a4531",x"5c4632",x"5b4531",x"5f4733",x"59432f",x"553f2d",x"543f2d",x"543f2c",x"56412f",x"584330",x"523e2d",x"58422f",x"55412f",x"56412e",x"56422f",x"543f2e",x"554130",x"574230",x"4f3c2b",x"543f2d",x"55412e",x"544030",x"54402f",x"523f2f",x"564230",x"564231",x"54402e",x"56422f",x"584332",x"513e2e",x"4d3b2b",x"513e2d",x"4e3c2d",x"4d3c2d",x"53402f",x"523f2e",x"4f3e2e",x"4b3a2a",x"493929",x"4b3a2c",x"4a3b2d",x"4f4032",x"564638",x"5a4a3c",x"5a4a3c",x"150e07",x"4f3925",x"392819",x"3a2819",x"352517",x"322314",x"342416",x"171009",x"664a32",x"453121",x"38291c",x"342517",x"39291a",x"392819",x"312215",x"312316",x"342516",x"2f2013",x"342517",x"342417",x"302114",x"332517",x"332416",x"312315",x"302114",x"2f2013",x"2b1e11",x"302114",x"342416",x"312215",x"322316",x"2e2013",x"2e2013",x"2f2114",x"322315",x"2e2013",x"312215",x"271b0f",x"281c10",x"2d2013",x"2b1e12",x"2a1d11",x"271b10",x"2c1f13",x"2c1f13",x"24190e",x"271b10",x"2b1e12",x"251a0f",x"20160c",x"2b1e12",x"2a1d11",x"21170d",x"21170d",x"21170d",x"20160c",x"1f150b",x"22170d",x"21170e",x"1d160f",x"4a3727",x"473524",x"463425",x"402f22",x"3e2d1f",x"3b2b1c",x"392819",x"3d2b1b",x"392819",x"372617",x"382718",x"3a281a",x"3e2c1c",x"3b2a1b",x"3b2a1b",x"392819",x"3b2a1a",x"362718",x"342517",x"382819",x"342516",x"332416",x"3c2b1b",x"3b2a1b",x"362618",x"352618",x"352517",x"332416",x"2f2013",x"2c1e12",x"312215",x"322315",x"322316",x"2e2013",x"2b1e12",x"2b1d11",x"281c10",x"261a0f",x"25190e",x"25190e",x"24190e",x"20150b",x"20160c",x"23180e",x"21160d",x"21160d",x"21170d",x"21160d",x"20170d",x"231a11",x"281d14",x"261d15",x"251c14",x"261d14",x"231c15",x"231b14",x"271e15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"261d15",x"261d15",x"2c1f16",x"2e1f15",x"2f1e12",x"342114",x"26170b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"1c1108",x"1f1209",x"1a1008",x"170f07",x"170f07",x"170f07",x"1d1108",x"201309",x"1a1008",x"1b1008",x"1d1108",x"1d1108",x"1e1208",x"201309",x"1d1108",x"1d1108",x"1a1008",x"150e07",x"1f1208",x"1c1108",x"1f1309",x"1b1108",x"221409",x"1f1309",x"150e07",x"1d1208",x"1e1208",x"24150a",x"150e07",x"1d1208",x"1d1108",x"190f07",x"150e07",x"150e07",x"201308",x"1e1208",x"1f1309",x"1c1108",x"1c1108",x"191008",x"17110a",x"171009",x"1a130c",x"19130c",x"19130c",x"462914",x"351e0f",x"371f0e",x"301c0d",x"341e0e",x"402512",x"412611",x"3e2410",x"3a210f",x"1a1008",x"1c1108",x"28170b",x"1b1007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"1b150e",x"201811",x"221a12",x"221a12",x"4c2c14",x"331d0d",x"301a0b",x"2e190b",x"361e0d",x"341d0c",x"29170a",x"2b1609",x"331c0c",x"2e190b",x"301a0b",x"38200e",x"26160a",x"150e07",x"150e07",x"4d3726",x"271e17",x"150e07",x"1d1108",x"211409",x"332318",x"261f18",x"27160a",x"2d1a0b",x"1d1108",x"3a200e",x"453124",x"4c392d"),
(x"6c543f",x"6c543f",x"4c3d30",x"45372b",x"46382b",x"47392d",x"4d3d30",x"4e3e30",x"504134",x"4d3f32",x"4e3f32",x"4d3e31",x"4d3e31",x"4f3f33",x"504032",x"4c3c2f",x"4c3b2d",x"4b3a2b",x"4d3b2d",x"4d3b2d",x"4c3a2c",x"4f3c2e",x"513f2e",x"4f3d2d",x"54402e",x"54402d",x"5b4532",x"5a4330",x"5d4631",x"5e4733",x"604833",x"604935",x"604834",x"5c4532",x"58432f",x"533e2d",x"513e2c",x"56412f",x"58422f",x"5b4431",x"56402d",x"59422d",x"57412d",x"553f2d",x"533f2d",x"523d2c",x"57412d",x"57422f",x"503e2b",x"54402e",x"56402e",x"523d2b",x"543f2c",x"53402d",x"513f2e",x"54412e",x"56422e",x"503c2a",x"523f2e",x"56412f",x"56412f",x"56412e",x"594431",x"594432",x"56422f",x"58422f",x"543f2d",x"533f2e",x"513d2c",x"4b3a2b",x"4d3b2b",x"4f3d2e",x"51402f",x"503e2e",x"4f3d2d",x"4d3c2e",x"4f3e2d",x"4d3b2c",x"4d3c2d",x"4c3d30",x"504235",x"524335",x"574738",x"574738",x"150e07",x"4b3522",x"372718",x"362517",x"382818",x"352517",x"352517",x"1b130b",x"674b32",x"42301f",x"35261a",x"372719",x"382819",x"362517",x"342416",x"312214",x"2c1e12",x"2d1f13",x"2e2013",x"362517",x"2e2013",x"322315",x"2a1d11",x"2e2013",x"2b1e11",x"2b1d11",x"2f2014",x"2c1e12",x"2e2013",x"2e2013",x"2e1f13",x"2e2013",x"2f2013",x"2e2013",x"2c1e12",x"2d1f12",x"2d1f13",x"2c1e11",x"2b1e12",x"2c1f12",x"2d2013",x"2c1f12",x"2e2013",x"291c11",x"261a0f",x"25190e",x"25190f",x"24180e",x"271a0f",x"23180d",x"25190e",x"25190e",x"281c10",x"20160c",x"1f150b",x"1f150b",x"1f150c",x"1f140b",x"21170e",x"1c160f",x"413122",x"463525",x"3f2e20",x"423123",x"3d2c1e",x"3b2a1b",x"372718",x"382718",x"3c2a1a",x"372617",x"3a291a",x"382718",x"3c2b1b",x"3b2a1b",x"3a2819",x"392819",x"382819",x"342416",x"2e2013",x"322315",x"302114",x"342416",x"342416",x"372718",x"362617",x"362617",x"2f2114",x"312215",x"2d1f12",x"2f2013",x"2f2114",x"2c1e12",x"2e2013",x"2a1d11",x"291c10",x"2a1d11",x"291c10",x"261a0f",x"261a0f",x"271b10",x"22170d",x"20150c",x"251a0f",x"25190f",x"261a0f",x"261a0f",x"23180d",x"1e140b",x"23180f",x"221911",x"231a12",x"241b13",x"201912",x"251c14",x"261d15",x"261d15",x"271d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281e16",x"281e16",x"2d2016",x"302117",x"312015",x"382416",x"22140a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"191008",x"170f07",x"25160a",x"1d1208",x"1f1209",x"1a1008",x"211409",x"231409",x"1e1208",x"1c1108",x"150e07",x"1c1108",x"180f08",x"26160a",x"26160a",x"221409",x"1c1108",x"1c1208",x"180f08",x"1c1108",x"1b1108",x"1c1108",x"26160a",x"28170a",x"27160a",x"25150a",x"26160a",x"29170a",x"27160a",x"26160a",x"29180b",x"29180b",x"2a190b",x"25160a",x"29180b",x"26160a",x"321d0e",x"29180b",x"26160a",x"1e1209",x"26170b",x"27170a",x"28170b",x"27170a",x"26160a",x"26160a",x"241409",x"211309",x"26160a",x"1b1108",x"261609",x"26160a",x"26160a",x"27160a",x"1e1208",x"231409",x"23150b",x"1c120b",x"19130c",x"171009",x"482a15",x"331d0f",x"372010",x"311d0d",x"3b2210",x"3a2110",x"412612",x"3b210f",x"3a210f",x"1d1208",x"1f1309",x"201309",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"150e07",x"150e07",x"170f07",x"1a1008",x"170f07",x"1d1108",x"180f08",x"1d1108",x"1a1008",x"211409",x"1b1008",x"1d1108",x"1e1208",x"24150a",x"1d1108",x"211409",x"231409",x"211409",x"1f1309",x"211409",x"191008",x"1f1309",x"201309",x"201309",x"1c1108",x"201309",x"1f1309",x"211409",x"231409",x"1f1209",x"1f1208",x"1f1208",x"1e1208",x"211409",x"201309",x"1d1108",x"201309",x"150e07",x"211409",x"1f1309",x"1e1208",x"1c1208",x"1b1108",x"1f1208",x"201309",x"211309",x"1d1108",x"1c1108",x"1a1008",x"221409",x"1c1108",x"1c1108",x"171009",x"1b140e",x"1e170f",x"211912",x"231b14",x"4f2e16",x"321c0c",x"321c0c",x"341c0c",x"351d0d",x"361e0d",x"321b0c",x"2f190b",x"28160a",x"2f1a0b",x"2f1a0a",x"361f0d",x"2e190b",x"150e07",x"150e07",x"473020",x"201810",x"150e07",x"1e1108",x"221409",x"332215",x"2a231c",x"28160a",x"271609",x"1d1108",x"371e0d",x"483427",x"483427"),
(x"6c543f",x"6c543f",x"4b3c2f",x"493a2d",x"4a3b2e",x"4a3c30",x"4e3f33",x"4f4134",x"4c3e31",x"4f4032",x"514235",x"504134",x"4f4032",x"504033",x"503e30",x"4c3d2f",x"47372a",x"48392c",x"48382b",x"4c3d2e",x"4e3e30",x"4e3d2d",x"544231",x"53402f",x"574331",x"574330",x"5a4330",x"5c4430",x"5b442f",x"5f4733",x"614a35",x"604934",x"5c4532",x"5d4631",x"5b4532",x"564231",x"594331",x"594331",x"55402d",x"543f2d",x"58412e",x"58412e",x"5a432f",x"55402e",x"543f2c",x"5a4431",x"56402e",x"55412d",x"55402d",x"56412e",x"543e2a",x"55412e",x"523d2b",x"513c2a",x"56412e",x"543d29",x"503d2c",x"533f2c",x"53402f",x"58422f",x"574130",x"584331",x"594432",x"594432",x"584231",x"574332",x"55402f",x"524130",x"524233",x"544231",x"4e3e2e",x"4e3c2e",x"4c3b2d",x"4f3d2d",x"513f30",x"4e3e2f",x"503e2f",x"53402e",x"554130",x"4c3c2d",x"4f4033",x"544435",x"58483b",x"58483b",x"150e07",x"47321e",x"312214",x"352416",x"342416",x"332415",x"332416",x"1c150d",x"664a32",x"423020",x"3b2c1d",x"38291b",x"372618",x"362618",x"3a2819",x"2f2114",x"332416",x"312215",x"2e2013",x"2d2013",x"342315",x"302114",x"2e2013",x"312215",x"312214",x"322316",x"2f2114",x"2f2013",x"2b1d11",x"2f2013",x"2c1e12",x"2f2014",x"2b1e12",x"291c10",x"2e2013",x"2b1d11",x"291c11",x"2e2013",x"2e1f13",x"2e1f13",x"2c1f12",x"281c10",x"2b1d12",x"2c1f12",x"281b10",x"25190f",x"281c10",x"251a0f",x"251a0f",x"25190f",x"21170c",x"21160c",x"26190e",x"24190e",x"21160c",x"1d140b",x"21170c",x"23180d",x"23190f",x"1d160f",x"433223",x"493626",x"3b2d1f",x"3c2d20",x"3b2b1d",x"372618",x"392819",x"322214",x"342416",x"352516",x"382718",x"392818",x"3b291a",x"3e2c1c",x"3d2b1c",x"3a2819",x"332416",x"322315",x"362618",x"342416",x"332416",x"3b291a",x"352516",x"332315",x"302113",x"372718",x"312214",x"312215",x"2f2114",x"322316",x"312215",x"2f2013",x"2f2114",x"2f2013",x"2e2013",x"2b1d11",x"23180d",x"26190e",x"271a0f",x"26190e",x"21160c",x"261a0f",x"25190e",x"25190e",x"23180d",x"23180d",x"20160c",x"20160c",x"21180e",x"221911",x"231a12",x"241b13",x"251c14",x"261d15",x"251d15",x"251d15",x"251d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"271e16",x"271e16",x"2f2117",x"2f2116",x"332115",x"362215",x"22150b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"180f08",x"180f08",x"201309",x"1f1309",x"1f1209",x"201309",x"211309",x"1f1209",x"211409",x"241509",x"150e07",x"211409",x"180f08",x"1d1208",x"24150a",x"24160a",x"26160a",x"251509",x"221409",x"27170a",x"231409",x"211409",x"231409",x"231409",x"211309",x"231409",x"241509",x"221409",x"28170a",x"27160a",x"28170b",x"26160a",x"27170a",x"26160a",x"2b190b",x"2c1a0c",x"2a190b",x"2b190b",x"28180b",x"2b1a0c",x"291a0c",x"291a0c",x"29190b",x"28180b",x"2a190b",x"28170b",x"27170b",x"2b190c",x"2e1c0d",x"2f1d0d",x"24150a",x"28170b",x"2d1b0c",x"2f1d0d",x"2b1a0c",x"2f1b0d",x"24150a",x"1f140a",x"1e130a",x"171009",x"17110a",x"432613",x"28180c",x"2d1a0d",x"2b190b",x"3b2310",x"392110",x"3c2310",x"3f2411",x"3a200e",x"201309",x"221409",x"211409",x"1e1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"221409",x"201309",x"1e1208",x"211309",x"221409",x"231409",x"1d1108",x"231409",x"251509",x"1f1309",x"26160a",x"1d1208",x"27170b",x"27170a",x"221409",x"221409",x"26160a",x"231409",x"26160a",x"26160a",x"2b190b",x"2a180b",x"23150a",x"27170a",x"1e1208",x"201309",x"201309",x"25160a",x"28170a",x"29170a",x"29170a",x"25160a",x"241509",x"27160a",x"25160a",x"28170a",x"29180b",x"2c1a0c",x"2b190b",x"241509",x"241509",x"26160a",x"251509",x"27160a",x"25150a",x"27160a",x"26150a",x"231409",x"221409",x"251509",x"27160a",x"24150a",x"26160a",x"27170a",x"27180c",x"27190e",x"261a11",x"291d13",x"211911",x"502f18",x"351d0d",x"311b0b",x"331c0c",x"341d0d",x"2c190b",x"2f1a0b",x"2d190a",x"371e0d",x"2e190b",x"331b0c",x"361d0d",x"351d0d",x"150e07",x"150e07",x"402c21",x"272019",x"160f08",x"1f1208",x"241509",x"322216",x"352d26",x"29170a",x"27160a",x"201309",x"3a200e",x"483325",x"483325"),
(x"6d5542",x"6d5542",x"4c3e32",x"4a3b2f",x"493b2f",x"4b3e32",x"4f4134",x"4c3e31",x"4e3f33",x"554436",x"544435",x"514134",x"544435",x"4f3f30",x"504033",x"4e3d2f",x"4f3e2f",x"503f31",x"544333",x"514031",x"544334",x"554332",x"594534",x"564230",x"594331",x"5b4632",x"5c4633",x"594431",x"5b4530",x"5e4833",x"644c36",x"634b35",x"604933",x"5d4633",x"5a4532",x"584332",x"533f2d",x"564230",x"574331",x"56412d",x"5b4431",x"5d4531",x"5d4631",x"57402d",x"5b4330",x"5b4531",x"5a4531",x"5a4431",x"5e4732",x"5a432f",x"5d4631",x"56412e",x"574130",x"5a4431",x"5c4531",x"55402e",x"5a4331",x"56412f",x"53402f",x"503c2c",x"54402d",x"59432f",x"584331",x"5a4532",x"5a442f",x"594533",x"594535",x"544030",x"534233",x"524132",x"534132",x"4f3e2f",x"514132",x"544232",x"564434",x"523f2f",x"534131",x"503e2e",x"513e2e",x"4f3e30",x"524234",x"544538",x"5c4b3c",x"5c4b3c",x"150e07",x"483321",x"392819",x"382719",x"372618",x"362617",x"342516",x"1b140e",x"5c432d",x"433121",x"382a1c",x"3d2e1f",x"38291a",x"332416",x"372718",x"302114",x"2f2013",x"2f2114",x"2c1f12",x"312214",x"322315",x"342517",x"322316",x"322315",x"342416",x"322316",x"2e1f13",x"322316",x"2d1f13",x"322215",x"302114",x"312213",x"2c1f12",x"2e2013",x"312114",x"2d1f12",x"291c11",x"2d1f12",x"2a1d11",x"281b10",x"2a1d11",x"2c1e12",x"2d1f12",x"2a1d12",x"251a0f",x"281b10",x"251a0f",x"281b10",x"271a0f",x"24190e",x"24180e",x"21160c",x"1f150b",x"24190e",x"23180e",x"20160c",x"20160c",x"20160c",x"21180e",x"1d160f",x"433223",x"4b3827",x"413123",x"403021",x"3c2c1e",x"3b2a1b",x"3c2a1a",x"382719",x"382719",x"382819",x"342416",x"332315",x"362617",x"392819",x"3b2a1a",x"39291a",x"342516",x"322315",x"382819",x"342416",x"2f2014",x"362617",x"342416",x"342416",x"322315",x"342517",x"362617",x"342416",x"362618",x"362618",x"322315",x"362618",x"332416",x"322215",x"342517",x"2b1d11",x"291c10",x"2e2013",x"2a1d11",x"2b1d11",x"24180e",x"22170d",x"1f150b",x"22170d",x"24180e",x"23180d",x"20160c",x"1e150c",x"22180e",x"211910",x"221911",x"251b12",x"261d15",x"261c14",x"251c14",x"261c13",x"271d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291f18",x"291f18",x"2e2016",x"302218",x"332218",x"362315",x"28190c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1008",x"180f08",x"180f07",x"1d1108",x"1b1108",x"1c1108",x"1a1008",x"1f1209",x"231409",x"211309",x"1d1108",x"180f07",x"150e07",x"150e07",x"150e07",x"231509",x"25150a",x"1c1108",x"211309",x"231409",x"201309",x"231509",x"231509",x"201309",x"1e1208",x"25160a",x"25160a",x"221409",x"1c1108",x"1e1208",x"27170a",x"27160a",x"231409",x"27160a",x"29170a",x"231409",x"241509",x"241509",x"221409",x"25150a",x"26160a",x"201309",x"27170a",x"27170a",x"201309",x"25150a",x"24150a",x"231509",x"29170b",x"29170a",x"26160a",x"27160a",x"25160a",x"28170b",x"27170a",x"27170b",x"2b190b",x"29180b",x"27180c",x"24160b",x"1e130a",x"23150b",x"54331b",x"321d0e",x"321d0f",x"2b180b",x"361f0e",x"361e0d",x"3d2310",x"3a210f",x"38200e",x"211409",x"231409",x"29180b",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"1f1208",x"1d1108",x"1d1208",x"1f1208",x"1c1108",x"1d1108",x"251509",x"211309",x"231409",x"221409",x"211409",x"25150a",x"211409",x"241509",x"26160a",x"29180b",x"27170a",x"231409",x"241409",x"211308",x"231409",x"211309",x"241509",x"25160a",x"28170b",x"221409",x"211309",x"1e1108",x"26160a",x"241409",x"28170a",x"2b190b",x"28170a",x"251509",x"261509",x"241509",x"27170a",x"29180b",x"29180b",x"29180b",x"241509",x"221309",x"231509",x"2c190b",x"1f1309",x"25160a",x"25150a",x"29180b",x"28180b",x"29190b",x"26160a",x"241509",x"27160a",x"26160a",x"231409",x"221409",x"28170a",x"28190c",x"2f1d11",x"2a1c12",x"241911",x"3e220f",x"381e0d",x"301a0b",x"341d0c",x"3a210f",x"321c0c",x"321c0c",x"281609",x"321b0b",x"29170a",x"351d0d",x"39200e",x"361e0d",x"150e07",x"160e07",x"48372b",x"28221b",x"161009",x"201308",x"26160a",x"402f22",x"332b24",x"2a170a",x"28170a",x"1e1208",x"3a200e",x"463123",x"463123"),
(x"5e4a3a",x"5e4a3a",x"4a3d31",x"4b3c2f",x"4a3b2e",x"4d3e30",x"4d3e31",x"504033",x"4d3d30",x"4e3e31",x"4e3e30",x"534335",x"554436",x"534332",x"504030",x"514031",x"554232",x"554333",x"514131",x"534233",x"574535",x"584535",x"574330",x"544231",x"5a4532",x"5a4431",x"5f4832",x"5a452f",x"5b4532",x"604730",x"5a432e",x"5b432f",x"513d2d",x"4e3b28",x"544130",x"564130",x"554130",x"574231",x"584332",x"584231",x"58422e",x"594331",x"5b4430",x"5e4733",x"594431",x"644c35",x"5f4733",x"5f4832",x"614934",x"5b4530",x"5c4632",x"58412d",x"5c4633",x"5f4632",x"5a432f",x"57422f",x"55402e",x"594432",x"594331",x"55412e",x"57422f",x"56412f",x"55402f",x"523d29",x"4e3a2a",x"503c2a",x"554231",x"594535",x"574332",x"544232",x"554233",x"534232",x"503e2e",x"534233",x"524030",x"534130",x"503d2e",x"53402f",x"544130",x"503e2f",x"524233",x"504134",x"584739",x"584739",x"150e07",x"483321",x"3a2919",x"372617",x"362617",x"382718",x"38271a",x"1d1710",x"5e432d",x"402f20",x"37281c",x"38281b",x"2c1e13",x"22160a",x"362617",x"352517",x"302114",x"322316",x"312215",x"2f2114",x"342415",x"332416",x"372718",x"352517",x"342416",x"352517",x"322316",x"2e2013",x"352517",x"312215",x"352517",x"2e2013",x"2e2013",x"302114",x"2f2013",x"2d1f12",x"2c1e12",x"2d1f13",x"2e1f13",x"2c1e12",x"281b10",x"2c1d11",x"291c10",x"25190e",x"1f140a",x"1f1309",x"261a0f",x"24190e",x"24190e",x"281c10",x"24190e",x"23180d",x"23180d",x"23180e",x"23180e",x"21170d",x"23180e",x"21170d",x"23180f",x"1f1912",x"3f2f21",x"4f3b29",x"433224",x"3e2e20",x"413020",x"3d2c1d",x"3b2a1a",x"3a291a",x"372718",x"3a2819",x"372718",x"352516",x"392718",x"362516",x"3a2818",x"322315",x"281a0d",x"27180b",x"2f2113",x"382718",x"3a2819",x"322316",x"352517",x"382718",x"342415",x"352517",x"352517",x"342517",x"382719",x"392819",x"362618",x"382819",x"352517",x"302114",x"2c1e12",x"2d1f12",x"2a1d11",x"2c1e12",x"2a1d11",x"271b0f",x"23180d",x"24190e",x"281b10",x"23180d",x"1e140b",x"22170d",x"1c130a",x"1e140b",x"1b120a",x"1c140c",x"231a10",x"261b13",x"261c13",x"231b12",x"241c13",x"261d15",x"261d15",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2018",x"2a2018",x"31231a",x"302117",x"312116",x"2b1a0d",x"28180c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"190f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f08",x"191008",x"150e07",x"160e07",x"160f07",x"150e07",x"1a1008",x"150e07",x"170f07",x"160f07",x"1a1008",x"150e07",x"170f08",x"160f07",x"170f07",x"1e1308",x"1a1008",x"1a1008",x"1a1008",x"1c1108",x"191008",x"170f08",x"191008",x"180f08",x"191008",x"1c1108",x"170f07",x"180f08",x"1c1108",x"170f08",x"180f08",x"180f08",x"180f08",x"191008",x"160f07",x"1c1108",x"150e07",x"1a1108",x"170f07",x"170f07",x"190f08",x"27160a",x"2d1a0c",x"28180c",x"2a1a0f",x"23160d",x"25180e",x"3e2312",x"331d0e",x"351f10",x"2a180b",x"361e0d",x"351d0d",x"3a200f",x"3c210f",x"3e2410",x"221409",x"241509",x"25150a",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"26160a",x"191008",x"1b1108",x"180f08",x"1e1209",x"1b1108",x"221409",x"191008",x"201409",x"211409",x"22140a",x"1d1209",x"1d1209",x"22140a",x"23150a",x"25160a",x"211409",x"28170b",x"180f08",x"231509",x"1c1108",x"211409",x"25160a",x"1d1209",x"201309",x"180f07",x"1c1108",x"1a1008",x"221409",x"201309",x"201309",x"201309",x"241509",x"25160a",x"23150a",x"201309",x"23150a",x"201309",x"24150a",x"211309",x"1e1108",x"201208",x"1b1108",x"211309",x"1e1108",x"1c1108",x"1d1208",x"1e1208",x"1d1108",x"1d1108",x"221409",x"1c1108",x"221409",x"231409",x"211409",x"1e1108",x"251509",x"27170c",x"27190d",x"2a1a10",x"231911",x"231911",x"442611",x"331c0c",x"331c0c",x"381f0e",x"2e1a0b",x"311b0c",x"301b0b",x"331c0c",x"2e190a",x"331c0c",x"371f0e",x"39200f",x"160e07",x"170f07",x"341d0d",x"281f17",x"18110a",x"241509",x"261509",x"472e1d",x"322b23",x"29170b",x"28160a",x"1c1108",x"3f2310",x"453124",x"453124"),
(x"6b5440",x"6b5440",x"4d4034",x"493b2e",x"493b2e",x"4e3f32",x"4e3d2f",x"4d3d2f",x"4e3d2f",x"4d3c2e",x"52402f",x"524031",x"544333",x"514131",x"524233",x"534132",x"534030",x"503f31",x"524132",x"574435",x"564333",x"524030",x"574432",x"5a4533",x"5e4835",x"5e4833",x"614a36",x"604935",x"5e4732",x"644b36",x"604934",x"5c4632",x"5d4732",x"5a4532",x"574331",x"564230",x"584331",x"564130",x"56422e",x"5a4430",x"5b4531",x"5b4530",x"5f4732",x"644b35",x"5f4732",x"624b34",x"5d4530",x"614731",x"5a422d",x"5b432e",x"5a432d",x"5e4631",x"5a432d",x"59432d",x"5a4431",x"574230",x"594330",x"5b4431",x"5d4531",x"5e4630",x"604631",x"604832",x"5d4630",x"5b432f",x"5b4532",x"5e4733",x"5a4431",x"594533",x"5a4635",x"554231",x"574433",x"554333",x"554233",x"544332",x"4f3f2e",x"584230",x"503e2f",x"513f30",x"4a392b",x"4c3a2b",x"514132",x"534335",x"594738",x"594738",x"150e07",x"45311e",x"392819",x"392819",x"3b2a1a",x"3a2819",x"3c2b1c",x"1d1610",x"674b33",x"4a3725",x"3f2f20",x"37281b",x"38281b",x"382818",x"382718",x"2f2014",x"322315",x"362517",x"372718",x"382718",x"382718",x"342516",x"372718",x"362617",x"352517",x"362718",x"322315",x"2e2013",x"342416",x"362618",x"2b1d11",x"322315",x"2c1e12",x"302114",x"302114",x"2b1e11",x"2d1f12",x"2e2013",x"2e2013",x"2d1f12",x"2e1f13",x"2d1f12",x"271a0f",x"2a1d11",x"2b1d11",x"2b1d11",x"291c11",x"271b10",x"281c10",x"24180e",x"22170d",x"281c10",x"25190e",x"23180d",x"23180e",x"23180e",x"23180e",x"21170d",x"231910",x"201913",x"3b2c20",x"4c3828",x"433324",x"433224",x"453223",x"3d2c1c",x"362617",x"3d2a1a",x"422f1d",x"3e2b1b",x"3a2819",x"3a2919",x"392818",x"3b291a",x"372617",x"332315",x"372617",x"372718",x"342416",x"352517",x"3a2919",x"352517",x"322315",x"392819",x"3a2819",x"372718",x"372718",x"3a291a",x"382718",x"332416",x"322315",x"312215",x"332316",x"312214",x"2d1f12",x"2c1f12",x"281b10",x"291c10",x"291d11",x"2b1e11",x"291c10",x"25190e",x"281c10",x"291c10",x"22170d",x"23180d",x"1f150b",x"1e140b",x"20170d",x"20180f",x"20170e",x"241a11",x"241a11",x"261c13",x"261c13",x"251c13",x"251c13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2018",x"2a2018",x"2f2117",x"2f2118",x"302016",x"321e10",x"321e10",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"1a1008",x"422511",x"2f1b0c",x"311c0d",x"321d0d",x"331d0d",x"341e0e",x"38200f",x"361f0e",x"301c0c",x"351d0d",x"2d190b",x"301b0c",x"28170a",x"2f1b0c",x"331d0d",x"361f0e",x"351e0e",x"351e0d",x"2f1a0c",x"331c0d",x"361f0e",x"361f0e",x"351e0d",x"331d0d",x"2e1a0b",x"341d0c",x"331d0c",x"361e0d",x"361e0d",x"311c0d",x"371f0e",x"39200e",x"361f0e",x"351e0d",x"3a210f",x"361f0e",x"39200e",x"3a200f",x"3c210f",x"39200f",x"3a210f",x"371f0e",x"39210f",x"3b2210",x"3a2210",x"3c2311",x"3a2210",x"3b220f",x"39200e",x"38200f",x"361f0e",x"38200f",x"3e2411",x"3d2310",x"3c2311",x"3c2311",x"402512",x"1f1309",x"1c1108",x"351f10",x"2b1a0e",x"26180e",x"2b1a0f",x"3f2412",x"392010",x"341e0e",x"2f1b0c",x"37200e",x"321d0d",x"39210f",x"371f0e",x"3c220f",x"231409",x"27170a",x"28170b",x"17100a",x"171009",x"150e07",x"150e07",x"150e07",x"1f1309",x"462914",x"432813",x"482b15",x"4c2e17",x"4b2d15",x"472a14",x"4c2f17",x"4a2c15",x"462914",x"452813",x"3c220f",x"402511",x"452913",x"472914",x"412612",x"3d220f",x"412511",x"462914",x"4b2c16",x"412510",x"442812",x"3b210f",x"432612",x"3f2411",x"432712",x"432713",x"422612",x"402511",x"3f2511",x"3b220f",x"3d220f",x"3a200e",x"3b210f",x"3a200e",x"3d2310",x"3f2310",x"402510",x"3f2411",x"3d2411",x"402612",x"452813",x"3e2310",x"422612",x"412611",x"3d2210",x"3e2310",x"3f2410",x"381f0d",x"2e190a",x"371e0c",x"2e1a0a",x"351d0c",x"361e0d",x"422611",x"3f2410",x"150e07",x"29180b",x"24170b",x"2a1a0f",x"24180f",x"20160e",x"452711",x"351d0c",x"341c0c",x"2c190b",x"2a170a",x"341d0d",x"311b0c",x"301b0b",x"2a170a",x"321c0c",x"38200e",x"38200e",x"160e07",x"191008",x"351e0d",x"29221a",x"18110a",x"27160a",x"271609",x"362213",x"373028",x"29170b",x"27160a",x"1e1208",x"3b210f",x"443125",x"443125"),
(x"6e5642",x"6e5642",x"514235",x"4b3d31",x"4d3d2f",x"4f3e2f",x"4f3e2f",x"4e3d2d",x"48382a",x"523f2e",x"4d3c2d",x"503f2f",x"523f2f",x"554433",x"534232",x"534231",x"503f2f",x"544130",x"544231",x"564333",x"584433",x"5c4735",x"584432",x"584432",x"5b4634",x"624b38",x"614b36",x"654d39",x"634b36",x"5f4935",x"614832",x"654d37",x"634b36",x"614934",x"5e4732",x"5a4531",x"5f4935",x"604934",x"5d4733",x"624a35",x"5a442f",x"5d442f",x"604732",x"5d4630",x"62472f",x"5d452e",x"624831",x"5f4731",x"614933",x"654a32",x"604730",x"614933",x"5d4531",x"634a33",x"604831",x"59432f",x"5b4330",x"5e4631",x"614832",x"614833",x"614831",x"604831",x"614933",x"614833",x"5f4732",x"5d4632",x"614936",x"5a4533",x"5a4632",x"594432",x"594534",x"564434",x"564333",x"544232",x"4e3d2f",x"533f2e",x"523f2f",x"4d3d2d",x"523f2f",x"503e2f",x"4e3e30",x"544435",x"564536",x"564536",x"150e07",x"4b3623",x"3b2a1a",x"362617",x"382718",x"3b2a1a",x"3d2d1d",x"201911",x"6a4e36",x"493725",x"402f20",x"3b2b1d",x"3d2c1d",x"372718",x"332416",x"312214",x"362718",x"382718",x"382819",x"3b2a1a",x"382718",x"362618",x"382718",x"322315",x"362517",x"352517",x"322315",x"322315",x"312215",x"322315",x"322316",x"342416",x"2f2114",x"332416",x"2e2013",x"2c1e12",x"2b1e11",x"322316",x"2d2013",x"2d2013",x"2d1f13",x"2c1f12",x"2b1d11",x"2d1f12",x"2b1d11",x"2b1d11",x"291c10",x"281c10",x"291c10",x"25190e",x"2c1f12",x"2b1e12",x"25190e",x"25190f",x"20150c",x"20150c",x"22170d",x"20150c",x"241911",x"221b14",x"3b2d20",x"5d4531",x"423123",x"463424",x"433223",x"412f20",x"3b291a",x"3c2a1a",x"3b2a1a",x"3d2b1b",x"3d2b1b",x"402d1d",x"3c2a1b",x"402e1d",x"402d1c",x"402d1c",x"3a2919",x"392818",x"392818",x"362616",x"3a2919",x"382718",x"3a291a",x"3a281a",x"342416",x"3a2819",x"322215",x"362617",x"342416",x"322315",x"352517",x"2f2114",x"332416",x"322315",x"342416",x"322316",x"291d11",x"2e2013",x"2a1d11",x"271a0f",x"271b10",x"261a0f",x"261a0f",x"23180e",x"20160c",x"21170d",x"20160c",x"1e140b",x"20160c",x"20160d",x"231910",x"22190f",x"251b12",x"221911",x"251c12",x"261b13",x"231b12",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291f18",x"291f18",x"302218",x"2f2016",x"332318",x"362112",x"362112",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"3e2310",x"2e1a0b",x"2d190b",x"2f1a0c",x"341d0d",x"301a0b",x"331c0d",x"361f0e",x"341d0d",x"341d0d",x"2d190b",x"2c190b",x"301c0c",x"2e1b0c",x"321c0d",x"351e0e",x"39210f",x"331d0d",x"311b0c",x"311a0b",x"311b0c",x"351d0d",x"351e0e",x"38200e",x"2f1b0c",x"301b0c",x"2c180b",x"301a0c",x"311b0b",x"2e1a0b",x"321c0c",x"351d0d",x"351d0d",x"321c0c",x"39200e",x"39200f",x"3b2310",x"3b2211",x"331e0e",x"3a2210",x"3c2310",x"39200f",x"3a210f",x"38200f",x"3a200f",x"381f0e",x"371f0d",x"371e0d",x"371e0d",x"38200e",x"351d0d",x"371f0e",x"3b2210",x"3d2411",x"3b2210",x"3d2411",x"382110",x"1e1209",x"321e0f",x"291b0f",x"342011",x"27190e",x"291a0e",x"402412",x"381f0f",x"2d1a0c",x"2e1b0c",x"38200f",x"351d0d",x"3b2310",x"381f0e",x"39200f",x"241509",x"27170a",x"28170b",x"19130c",x"1a130c",x"171009",x"180f08",x"1d1208",x"211409",x"2f1b0c",x"2f1b0c",x"321c0d",x"361f0e",x"37200f",x"351e0e",x"351e0e",x"311c0d",x"341e0e",x"392110",x"3c2311",x"3d2411",x"37200f",x"3a210f",x"37200f",x"331d0e",x"392110",x"3d2411",x"3c2311",x"341e0e",x"37200f",x"331d0e",x"2f1b0c",x"2e1a0b",x"321c0c",x"311c0c",x"351d0d",x"351d0d",x"39210f",x"3c220f",x"371f0e",x"381f0e",x"331c0c",x"39200f",x"3a210f",x"39200e",x"38200e",x"36200f",x"37200f",x"341d0d",x"321b0c",x"321c0c",x"331c0d",x"39200f",x"39200f",x"351e0e",x"351d0d",x"351d0d",x"361e0d",x"331c0c",x"341d0c",x"361e0d",x"361e0d",x"351d0d",x"361e0d",x"150e07",x"28170b",x"331e10",x"2f1e0f",x"2c1b0f",x"281a0f",x"472913",x"331c0c",x"381f0e",x"321c0c",x"321c0c",x"361e0d",x"311c0c",x"311c0c",x"2f1a0b",x"371e0d",x"371f0e",x"361e0d",x"160e07",x"170f07",x"4b3628",x"2d231b",x"18110a",x"241409",x"271609",x"3a2313",x"383129",x"29170b",x"251509",x"1f1209",x"3b2110",x"473327",x"473327"),
(x"66513e",x"66513e",x"4c3e32",x"4d3f32",x"4f3f31",x"4b3b2d",x"4d3c2d",x"4f3d2c",x"4b3a2b",x"4f3c2a",x"503e2d",x"544131",x"564332",x"564333",x"534132",x"5a4634",x"544131",x"564333",x"5b4635",x"594635",x"5a4634",x"5d4936",x"604a37",x"624b38",x"624b38",x"624b36",x"624c38",x"614a35",x"5e4936",x"644c39",x"614a36",x"614a35",x"604a35",x"5f4732",x"5d4632",x"5e4731",x"5d4631",x"5b4431",x"5b4531",x"5f4632",x"5d452f",x"5d442e",x"654a32",x"624933",x"614932",x"684d34",x"644933",x"664c35",x"624931",x"664c33",x"664b34",x"634931",x"614933",x"684e38",x"634a35",x"644c37",x"644c36",x"624a33",x"5f4832",x"5e4732",x"614831",x"634a32",x"614933",x"5d4632",x"614933",x"5f4732",x"5b4734",x"5b4532",x"584330",x"544030",x"54412f",x"534132",x"554334",x"574433",x"534030",x"574433",x"554130",x"534131",x"513e2d",x"544232",x"514132",x"574536",x"594738",x"594738",x"150e07",x"4c3725",x"402e1e",x"402e1e",x"3d2c1d",x"3b2a1a",x"3d2d1e",x"201810",x"654932",x"483523",x"412f20",x"3a2b1b",x"39291a",x"352517",x"302114",x"362617",x"382718",x"312215",x"342415",x"342416",x"322315",x"332416",x"352617",x"3a291a",x"362718",x"3a291a",x"362617",x"3a291a",x"342416",x"372719",x"362618",x"342516",x"352517",x"372719",x"322416",x"372719",x"382819",x"342516",x"2f2214",x"2a1d11",x"2e2013",x"2d2013",x"2e2013",x"2b1d11",x"2c1e11",x"291c11",x"271a0f",x"271a0f",x"281b10",x"24190e",x"21170c",x"281c10",x"291c10",x"281b10",x"23180e",x"24190e",x"21170d",x"21170d",x"281c13",x"221b15",x"382b1f",x"604834",x"483628",x"413123",x"463524",x"443122",x"423020",x"3e2d1d",x"3c2b1c",x"3b2a1a",x"3a291a",x"3b291a",x"3a2819",x"3d2b1b",x"3e2b1b",x"3b2a1a",x"352517",x"392819",x"382718",x"352516",x"352517",x"332315",x"342415",x"382718",x"382617",x"352517",x"392819",x"392819",x"392819",x"3c2a1b",x"322316",x"352618",x"2f2114",x"352618",x"312215",x"332416",x"332416",x"312216",x"2e2014",x"2d2014",x"2f2115",x"2c1e12",x"291d11",x"25190f",x"23180d",x"23180e",x"281c10",x"20160c",x"20150c",x"22170e",x"20170d",x"21170d",x"20180f",x"231810",x"211810",x"251b12",x"211911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2018",x"2a2018",x"31241a",x"312218",x"312116",x"352011",x"352011",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"180f08",x"38200f",x"321d0e",x"2e1b0c",x"2f1a0b",x"37200e",x"311c0c",x"341d0d",x"351e0e",x"321d0d",x"341e0d",x"321c0d",x"2d1a0b",x"301b0c",x"2f1a0b",x"28170a",x"341e0d",x"2e1a0c",x"311c0d",x"2f1a0b",x"351d0d",x"39210f",x"2d1a0b",x"361f0e",x"38200f",x"3a2210",x"38200f",x"37200f",x"361f0f",x"351e0e",x"351e0e",x"361f0e",x"37200f",x"361f0e",x"39200f",x"3a210f",x"38200e",x"351e0e",x"371f0e",x"3c2311",x"3f2512",x"3b2311",x"3c2310",x"39210f",x"3b2210",x"39200f",x"39200f",x"361f0e",x"38200e",x"371f0e",x"3b210f",x"361e0d",x"381f0e",x"3a210f",x"392110",x"331d0e",x"412713",x"3e2411",x"191008",x"321d0f",x"342011",x"291a0f",x"2c1b0f",x"291a0f",x"3d2211",x"301b0d",x"29180b",x"241509",x"2c180b",x"3a210f",x"331d0d",x"361f0e",x"39200e",x"241509",x"27170a",x"27170a",x"1a130c",x"1a130c",x"17110a",x"150e07",x"191008",x"1a1008",x"2e190b",x"2c190b",x"2d190b",x"2f1a0b",x"351e0e",x"3a2210",x"341e0e",x"2f1b0c",x"341e0e",x"341f0e",x"341d0d",x"351f0e",x"38200f",x"38200f",x"2c190b",x"371f0e",x"3d2310",x"3a210f",x"3a210f",x"37200f",x"341e0e",x"36200f",x"3d2411",x"3a210f",x"311b0c",x"351e0d",x"371f0e",x"361e0d",x"39200f",x"371f0e",x"38200f",x"38200e",x"3b220f",x"371f0e",x"3b220f",x"3a200f",x"39210f",x"38200f",x"3c2210",x"371f0e",x"361e0d",x"37200e",x"38200e",x"351d0d",x"3c2310",x"3a2210",x"3a2110",x"3b2310",x"3c2311",x"39210f",x"3b2210",x"3d2410",x"38200e",x"38200e",x"39210f",x"150e07",x"28170b",x"2d1a0d",x"2f1c0f",x"28190e",x"21160d",x"4b2b14",x"301a0b",x"381f0e",x"351d0d",x"361e0d",x"351d0d",x"351e0d",x"331c0c",x"351d0d",x"311b0c",x"361e0d",x"341d0d",x"160e07",x"180f07",x"3e291b",x"2a2018",x"18120b",x"261509",x"281709",x"362111",x"332b23",x"28170b",x"241509",x"211409",x"392010",x"4d3a2d",x"4d3a2d"),
(x"6c5542",x"6c5542",x"514337",x"4b3d31",x"483a2e",x"4d3b2c",x"4b3a29",x"4f3c2b",x"4c3a2a",x"4a382a",x"493828",x"463527",x"503e2e",x"544030",x"5b4633",x"554131",x"574331",x"554130",x"574332",x"5a4634",x"614c39",x"5e4a37",x"5f4936",x"5d4734",x"614b37",x"604b37",x"604a37",x"5d4633",x"5a4634",x"5f4b37",x"604b37",x"614a37",x"614937",x"624a36",x"5f4733",x"5d4532",x"5b4632",x"604732",x"5f4830",x"604730",x"5e4631",x"5c432e",x"563d26",x"573e27",x"5a422c",x"624831",x"674c32",x"664a31",x"614830",x"664a31",x"61472f",x"604731",x"664d35",x"644b35",x"664c35",x"684d36",x"5f4833",x"604832",x"624933",x"614831",x"59432d",x"5d4732",x"5a4532",x"5f4835",x"5e4733",x"5f4733",x"5e4936",x"5c4633",x"584431",x"584330",x"513f2e",x"534131",x"584736",x"534131",x"493a2d",x"46372a",x"534131",x"524031",x"54412f",x"4f3d2f",x"4e3e30",x"544436",x"554436",x"554436",x"150e07",x"493422",x"3b2a1a",x"3b291a",x"3c2a1b",x"382718",x"38281a",x"1f1710",x"543c29",x"413020",x"3c2c1e",x"3c2b1d",x"392a1b",x"312215",x"312215",x"342416",x"342416",x"2f2114",x"342415",x"352516",x"372617",x"332315",x"25180b",x"27190d",x"332215",x"392818",x"362617",x"3a281a",x"382819",x"312215",x"322315",x"362618",x"302215",x"322316",x"2e2013",x"322316",x"342416",x"302114",x"312214",x"2a1d11",x"281b0f",x"2f2114",x"2b1d11",x"2d1f13",x"2d1f13",x"271b10",x"24180e",x"281b10",x"261a0f",x"291c11",x"271a0f",x"281b0f",x"271b0f",x"22170d",x"1d1309",x"1b1109",x"21160c",x"20160c",x"2b1f15",x"231d16",x"382b20",x"5d4531",x"463526",x"463425",x"453424",x"453222",x"3e2c1c",x"3d2b1b",x"3f2c1c",x"392819",x"342416",x"362516",x"312214",x"362617",x"3a291a",x"392819",x"3c2a1b",x"3d2b1b",x"3a2919",x"332315",x"332315",x"352517",x"352516",x"352516",x"382718",x"342315",x"291a0b",x"27190d",x"332315",x"392819",x"3b2a1a",x"362617",x"332416",x"332416",x"2f2114",x"322316",x"352517",x"2d2013",x"281c10",x"2a1d11",x"2a1d11",x"271b10",x"261a0f",x"22170d",x"1f150b",x"21170c",x"1f150c",x"20150c",x"1d140b",x"20150c",x"20170d",x"1d150c",x"20170d",x"231810",x"22190f",x"1f170e",x"20170f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b2119",x"2b2119",x"302218",x"312319",x"342417",x"331e10",x"331e10",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"3b210f",x"351f0e",x"331e0e",x"351f0f",x"36200f",x"392110",x"37200f",x"351f0f",x"38200f",x"38210f",x"2a180b",x"301c0d",x"321d0d",x"37200f",x"301c0d",x"361f0f",x"3b2210",x"392110",x"392110",x"311d0d",x"38210f",x"361f0e",x"38200e",x"371f0f",x"361f0e",x"38200f",x"361f0e",x"321c0c",x"361f0e",x"2f1c0d",x"321d0d",x"331d0d",x"3a200f",x"371f0e",x"371f0e",x"3e2310",x"371f0e",x"38200e",x"392110",x"3b2310",x"3e2511",x"3c2311",x"39210f",x"37200f",x"371f0e",x"351e0d",x"3a200f",x"371f0e",x"3a210f",x"3c2311",x"3f2411",x"3c2311",x"3a2110",x"38200f",x"3d2411",x"412612",x"3d2411",x"211409",x"331e10",x"362010",x"382112",x"301e11",x"301d10",x"3f2411",x"331d0e",x"2f1a0c",x"1f1208",x"2c180b",x"37200f",x"321d0d",x"311c0d",x"371f0e",x"241509",x"28170b",x"26160a",x"19130c",x"19130c",x"17110a",x"171009",x"201309",x"201409",x"341e0e",x"321d0e",x"321d0e",x"341e0e",x"351f0e",x"3b2210",x"38200f",x"38200f",x"311c0d",x"321c0c",x"321d0d",x"3d2411",x"3b2310",x"36200f",x"36200f",x"3a210f",x"3b220f",x"38200f",x"3b210f",x"341d0d",x"2e1a0b",x"2d190b",x"311d0d",x"392110",x"36200f",x"392110",x"392110",x"3b2310",x"3a2110",x"3f2512",x"3c2310",x"3a210f",x"3a210f",x"39200f",x"3c2210",x"3c2310",x"3c2311",x"3e2511",x"412712",x"3c2311",x"3d2411",x"3b2310",x"3d2310",x"3a210f",x"3a210f",x"3b2310",x"3a2110",x"3c2310",x"3c220f",x"38200e",x"3c2311",x"3c2311",x"39200e",x"38200e",x"381f0e",x"150e07",x"27160a",x"2b190d",x"2c1b0f",x"28190e",x"22160d",x"432611",x"351e0d",x"381f0e",x"2f1b0c",x"321c0c",x"321c0c",x"311b0c",x"341c0c",x"341d0c",x"311c0c",x"321c0c",x"321c0c",x"160e07",x"190f07",x"3d281b",x"271e16",x"19120b",x"27160a",x"28160a",x"412917",x"28211a",x"28170b",x"221309",x"24150a",x"3d2210",x"4a362a",x"4a362a"),
(x"6c5643",x"6c5643",x"524437",x"4f3f31",x"4e3f31",x"4c3b2d",x"4d3b2a",x"52402f",x"584330",x"54402d",x"513e2c",x"513e2d",x"4e3d2e",x"4d3c2d",x"513e2f",x"513f2d",x"523e2e",x"544030",x"574433",x"574230",x"5a4534",x"5c4835",x"614b38",x"604a37",x"5f4a36",x"644d38",x"644d39",x"654e3a",x"634d39",x"664f3b",x"644d39",x"654e3a",x"644c39",x"644d39",x"664d39",x"634a34",x"614934",x"614933",x"614934",x"644b34",x"634b35",x"654a32",x"5c432c",x"5c442e",x"5b422b",x"5b422b",x"5e432c",x"62482f",x"654b33",x"634a31",x"654932",x"614830",x"614730",x"5d4631",x"624933",x"664c34",x"644a33",x"644b34",x"614832",x"604833",x"644c36",x"644c36",x"604a35",x"604732",x"5f4936",x"634c38",x"5e4733",x"5e4835",x"5d4835",x"594432",x"544130",x"503d2e",x"5b4836",x"544132",x"524031",x"4f3d2e",x"4d3c2c",x"4b3a2c",x"48382a",x"4c3b2b",x"4a3b2d",x"4e3f32",x"4e3f33",x"4e3f33",x"150e07",x"44311e",x"3c2a1a",x"3c2a1b",x"3d2b1b",x"3a2919",x"392819",x"201911",x"5b432d",x"4c3826",x"3d2c1e",x"3d2b1d",x"3d2c1d",x"372718",x"362517",x"362617",x"332316",x"352517",x"362517",x"342416",x"3b2a1a",x"372617",x"342415",x"312214",x"312114",x"2b1d11",x"302114",x"342415",x"342416",x"332416",x"312215",x"2f2014",x"322215",x"302214",x"322315",x"302114",x"332416",x"312214",x"2f2013",x"312215",x"2c1f12",x"322316",x"2d1f13",x"2c1f12",x"2b1d12",x"2b1e12",x"281b10",x"281c10",x"281b10",x"291c11",x"24180e",x"23180e",x"2b1e12",x"271a0f",x"21160c",x"20150c",x"1d130a",x"1d130a",x"241b12",x"241d16",x"33271d",x"543f2d",x"3f3123",x"423224",x"3f2f20",x"3e2d1d",x"402d1c",x"3d2b1b",x"372718",x"3c2a1b",x"3a2919",x"3f2c1c",x"3a2819",x"3b2a1b",x"392819",x"3e2c1c",x"3f2c1c",x"3c2a1b",x"3c2a1b",x"3c2a1b",x"352517",x"352517",x"342417",x"352517",x"3b2a1b",x"362616",x"352515",x"332315",x"2e2012",x"312014",x"302114",x"322314",x"332315",x"2e2013",x"312215",x"322315",x"322315",x"2c1f12",x"2d1f13",x"2a1d11",x"291c11",x"25190e",x"271b10",x"251a0f",x"23180d",x"21170d",x"20160c",x"20160c",x"1d140b",x"1e140b",x"20160c",x"21180e",x"21180e",x"21170e",x"22180f",x"20170f",x"20180f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2119",x"2a2119",x"2e2218",x"302218",x"332318",x"372012",x"372012",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a0f07",x"412511",x"2e190b",x"2d190b",x"2d190b",x"2d1a0b",x"2f1a0b",x"2f1b0c",x"2c190b",x"2e1a0b",x"311b0c",x"2a180a",x"2f1a0b",x"27160a",x"29160a",x"28160a",x"2b180b",x"2d190b",x"2e190b",x"331d0d",x"331d0d",x"321c0c",x"351e0e",x"2f1b0c",x"331d0d",x"38200f",x"361f0e",x"39200f",x"351e0e",x"311c0d",x"331d0d",x"361f0e",x"39210f",x"37200f",x"3e2512",x"3b2310",x"3e2511",x"3e2511",x"382110",x"3a2210",x"392110",x"402512",x"3f2512",x"3e2512",x"3c2311",x"3b2210",x"3b2210",x"371f0e",x"351d0d",x"361e0d",x"3b2210",x"3f2512",x"432813",x"3a2311",x"3e2512",x"3f2613",x"402713",x"402612",x"191008",x"2d1a0c",x"2d1a0d",x"321d0f",x"24180e",x"24170c",x"3e2210",x"351e0e",x"201308",x"251509",x"351c0c",x"3c2310",x"2f1b0c",x"311c0d",x"341d0d",x"221409",x"26170a",x"25160a",x"19130c",x"19130c",x"171009",x"17110a",x"150e07",x"1d1108",x"29170a",x"2d190b",x"2f1a0b",x"2e1a0b",x"311b0c",x"38200e",x"341d0d",x"341d0d",x"351d0d",x"311b0c",x"311b0c",x"341d0d",x"331c0c",x"2d190b",x"361e0d",x"351e0d",x"371f0e",x"361e0d",x"331d0d",x"2e190b",x"251408",x"29160a",x"29170a",x"2c180b",x"2a170a",x"2d1a0b",x"2f1b0b",x"341d0c",x"351d0d",x"361e0d",x"361e0d",x"341d0d",x"331d0d",x"351d0d",x"311b0b",x"2f1a0b",x"331c0c",x"301a0b",x"2f1a0b",x"331c0c",x"371f0e",x"321c0d",x"351e0e",x"3c230f",x"3a210f",x"361e0e",x"3d2310",x"3d2310",x"3d2310",x"3d2310",x"3a220f",x"3a210f",x"3d2311",x"3a2210",x"3e2511",x"150e07",x"2b1a0c",x"321e0f",x"342011",x"2f1e11",x"281a10",x"442611",x"361e0d",x"351d0d",x"3a210f",x"381f0d",x"331c0c",x"2f1a0b",x"331c0c",x"341d0c",x"331c0c",x"341d0d",x"351e0d",x"160e07",x"1a1008",x"3c281c",x"2f2319",x"18110a",x"27160a",x"28160a",x"3c2516",x"2b2119",x"26160a",x"221409",x"27170b",x"382010",x"4b3629",x"4b3629"),
(x"675341",x"675341",x"574739",x"504134",x"514032",x"524031",x"53402e",x"58422f",x"503c2b",x"4e3b2a",x"57422f",x"564230",x"574433",x"594635",x"5a4635",x"584431",x"5f4936",x"5d4733",x"5e4935",x"624c39",x"644f3c",x"654f3b",x"69513d",x"644d38",x"644c38",x"614a38",x"5e4834",x"594433",x"624c39",x"5e4835",x"624c38",x"604a37",x"614b38",x"654e39",x"664e38",x"644c36",x"644c37",x"6a513a",x"664c37",x"624a34",x"614932",x"614730",x"664c34",x"614932",x"664c34",x"674c34",x"654b34",x"694d33",x"684d33",x"664c34",x"644b32",x"6b4f35",x"664d34",x"664c34",x"6a4f37",x"674e37",x"634932",x"614731",x"5b4531",x"543f2d",x"594331",x"604935",x"5f4935",x"634b36",x"624c3a",x"624a36",x"624c37",x"604b37",x"614a36",x"5c4734",x"5e4836",x"5a4634",x"564534",x"554333",x"564333",x"554331",x"544131",x"513f2f",x"513f30",x"524030",x"534131",x"584637",x"524133",x"524133",x"150e07",x"4e3926",x"412f1f",x"3f2d1d",x"3c2a1b",x"362617",x"362517",x"1f1711",x"563e29",x"473423",x"3e2d1f",x"39291c",x"3b2a1c",x"332416",x"3a2a1b",x"3a2919",x"3b2a1a",x"3d2b1c",x"382819",x"3a291a",x"342415",x"322214",x"3a2919",x"3d2b1c",x"3c2b1b",x"3b2a1a",x"382819",x"382819",x"3a291a",x"362719",x"382819",x"362618",x"362719",x"372719",x"372819",x"362618",x"322315",x"2d1f13",x"2c1e12",x"25180c",x"2a1c11",x"2d1f12",x"2c1e12",x"2e1f13",x"2d1f13",x"2d1f13",x"2c1f13",x"281c10",x"291c11",x"2a1d11",x"2c1e13",x"2a1d11",x"23180d",x"261a0f",x"24190e",x"24190e",x"23180e",x"23180d",x"261d13",x"241d17",x"36291e",x"604833",x"473626",x"453525",x"473525",x"493524",x"433120",x"422f1e",x"3f2c1c",x"3c291a",x"372617",x"2f1e10",x"392718",x"3a291a",x"372718",x"3d2b1b",x"402d1d",x"3a291a",x"3f2d1e",x"3d2b1c",x"39281a",x"3d2b1c",x"342517",x"3c2b1b",x"352516",x"352416",x"392819",x"3a291a",x"3b291a",x"3b2a1a",x"3a291a",x"382819",x"3a291a",x"39291a",x"362617",x"362618",x"332417",x"362618",x"312316",x"2d2013",x"2c1e12",x"26190f",x"25190e",x"1e130a",x"22170d",x"22170d",x"21170c",x"20160c",x"21160d",x"20160c",x"21170d",x"21170e",x"21170f",x"20170d",x"21180f",x"21180f",x"20170e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2018",x"2a2018",x"2f2218",x"312318",x"322318",x"321d10",x"321d10",x"150e07",x"150e07",x"150e07",x"170f07",x"1f1209",x"1c1108",x"391f0d",x"351f0e",x"351f0f",x"36200f",x"361f0f",x"39200f",x"351e0e",x"3b2310",x"37200f",x"2e1b0c",x"2f1b0c",x"36200e",x"38210f",x"37200f",x"38200f",x"341e0e",x"331d0d",x"361e0e",x"321c0d",x"371f0e",x"371f0e",x"3a210f",x"3a210f",x"361f0e",x"341d0d",x"301b0c",x"351e0d",x"331d0d",x"311c0c",x"311c0c",x"321c0c",x"341d0d",x"341d0d",x"351e0d",x"351e0d",x"341d0d",x"371f0e",x"361f0e",x"37200e",x"321c0d",x"371f0e",x"3a2210",x"3a2210",x"3c2311",x"382110",x"38210f",x"3a2210",x"392210",x"3c2411",x"39210f",x"3d2310",x"3c2310",x"38210f",x"37200f",x"3a2210",x"3a2110",x"3d2411",x"191008",x"29180a",x"2a180b",x"2c1a0d",x"23160b",x"26170b",x"3f2411",x"331d0e",x"2d190b",x"27160a",x"311b0c",x"3c2210",x"38200e",x"351f0e",x"351e0d",x"221409",x"27170b",x"241509",x"19120b",x"19120c",x"171009",x"19110a",x"150e07",x"1a1008",x"28160a",x"2a170a",x"29170a",x"2b180a",x"2e190b",x"301b0b",x"2e190b",x"2e190a",x"2d180a",x"2e190a",x"2e1a0b",x"331c0c",x"351d0d",x"351f0e",x"3d2310",x"3a2210",x"3e2411",x"3a210f",x"38200e",x"351d0d",x"351d0d",x"311b0c",x"341d0d",x"351e0e",x"3a2210",x"38200f",x"39200f",x"39200f",x"38200f",x"392110",x"381f0e",x"3d2310",x"3b2210",x"402512",x"3e2511",x"3e2411",x"3a220f",x"361f0e",x"361f0e",x"381f0e",x"3c210f",x"3c2310",x"38200f",x"3b2210",x"3d2310",x"38200f",x"3c220f",x"3e230f",x"3a200e",x"361e0d",x"331c0c",x"321c0c",x"371e0d",x"351d0d",x"381f0e",x"160e07",x"25160a",x"2c1b0f",x"311f12",x"291a10",x"25190f",x"412510",x"381f0e",x"381f0e",x"3a210f",x"3f2310",x"371f0e",x"311b0b",x"38200e",x"321c0c",x"361f0e",x"361f0d",x"39200f",x"160e07",x"1a1008",x"3c291d",x"2f231b",x"18110a",x"27160a",x"28160a",x"3e2716",x"292019",x"241509",x"231409",x"29180b",x"3a200e",x"4b382a",x"4b382a"),
(x"5b4b3c",x"5b4b3c",x"514336",x"504133",x"513f31",x"503d2e",x"54402f",x"533f2e",x"503d2c",x"4f3b29",x"53402e",x"56412f",x"564332",x"55412f",x"534131",x"564331",x"564130",x"5f4936",x"614b38",x"634d39",x"604b37",x"69523d",x"664f3a",x"624b38",x"644d39",x"644d39",x"664e3a",x"614a36",x"624b37",x"644d3a",x"654d39",x"614b37",x"634d39",x"614b38",x"614b38",x"624a35",x"664d38",x"684e37",x"674e39",x"644c36",x"634932",x"664d34",x"624932",x"614832",x"5f4731",x"684d35",x"614831",x"644a32",x"644a31",x"604831",x"664b32",x"684c33",x"674c35",x"664c33",x"654b33",x"674d35",x"634a34",x"664d36",x"624a35",x"5f4936",x"5f4936",x"5e4836",x"614a38",x"5d4836",x"604a37",x"604a36",x"5e4936",x"5d4835",x"604a36",x"5e4935",x"594534",x"594633",x"564333",x"584533",x"544131",x"524031",x"53402e",x"523f2e",x"4d3d2d",x"4e3d2f",x"514032",x"514030",x"4f3f33",x"4f3f33",x"150e07",x"4f3925",x"402d1d",x"3c2a1a",x"3a291a",x"372618",x"3b2a1b",x"201811",x"573f2a",x"453323",x"3d2d1f",x"3c2c1e",x"39291b",x"342416",x"3a2819",x"352517",x"382719",x"352617",x"3a2a1a",x"3d2b1c",x"342515",x"312214",x"362618",x"342416",x"352517",x"332315",x"342416",x"392819",x"342416",x"382719",x"362618",x"322315",x"3a2919",x"382819",x"332416",x"322215",x"312215",x"2d1f12",x"322315",x"2f2013",x"2e2013",x"2b1e11",x"2c1e12",x"2a1d11",x"2d1f12",x"2a1d11",x"261a0f",x"2a1d11",x"2a1d11",x"291d11",x"2a1d11",x"2a1d11",x"261a0e",x"291c10",x"20150c",x"21160c",x"21170d",x"22170d",x"271c13",x"211b14",x"35281d",x"59422e",x"493627",x"463324",x"493625",x"473423",x"44301f",x"412d1c",x"3f2d1c",x"3d2b1b",x"3f2c1c",x"3f2c1c",x"3a291a",x"3f2d1c",x"3c2a1b",x"3b291a",x"412e1d",x"3b291a",x"3c2b1b",x"392819",x"3d2b1b",x"3d2b1c",x"3f2d1d",x"3d2c1c",x"332315",x"3a2818",x"392819",x"372618",x"382719",x"392819",x"332415",x"362618",x"342416",x"312215",x"342416",x"362517",x"312315",x"2f2114",x"2e2013",x"322215",x"2b1e11",x"291c11",x"2a1d11",x"271b10",x"23180d",x"22170d",x"23180d",x"1f150b",x"1f150c",x"1f150b",x"1e150c",x"20170d",x"1f160d",x"20160d",x"241a11",x"241a11",x"20170e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b2119",x"2b2119",x"2f2319",x"332319",x"332218",x"311f11",x"311f11",x"150e07",x"150e07",x"150e07",x"180f07",x"241509",x"221409",x"351d0b",x"341e0e",x"321d0d",x"361f0f",x"351f0f",x"361f0e",x"351e0d",x"321d0e",x"351e0e",x"331d0d",x"2c190c",x"392110",x"37200f",x"37200e",x"2e1a0b",x"301c0c",x"371f0e",x"341e0d",x"2d1a0c",x"301b0c",x"321d0d",x"392110",x"38200f",x"351e0d",x"3a210f",x"331d0d",x"3d2310",x"361f0e",x"371f0e",x"39200f",x"3a2110",x"3b2210",x"38200f",x"39210f",x"3b2310",x"3c2311",x"3e2511",x"37200f",x"3a2210",x"3c2311",x"3f2512",x"412613",x"402612",x"3d2511",x"3f2512",x"412612",x"3a2210",x"3b2311",x"3b2311",x"3c2311",x"3f2511",x"3e2412",x"402613",x"402612",x"371f0e",x"38200e",x"351d0d",x"1d1208",x"2c1a0c",x"321e0e",x"321e0f",x"2d1c0e",x"2b1a0d",x"432712",x"321c0e",x"2a170a",x"251509",x"331c0c",x"3b220f",x"38200e",x"3e2411",x"361f0e",x"221409",x"27170b",x"231409",x"19120b",x"19120b",x"17110a",x"1d130b",x"1e1208",x"1e1108",x"29170a",x"2a170a",x"2b180a",x"2d190a",x"311b0c",x"351d0d",x"331d0d",x"331d0d",x"301a0b",x"2d180a",x"2b170a",x"321b0b",x"361f0e",x"361f0e",x"361f0e",x"3b2210",x"3c2311",x"3c2311",x"37200f",x"37200f",x"38200e",x"311c0c",x"351e0e",x"39210f",x"351e0e",x"3b2210",x"321d0e",x"351e0e",x"36200f",x"311c0d",x"3b2210",x"3c2311",x"3b2310",x"39200f",x"3a220f",x"39200e",x"3a210f",x"38200e",x"371f0e",x"39200f",x"39200f",x"3b2210",x"3d2411",x"3e2511",x"3e2310",x"3d2310",x"3f2411",x"3e2411",x"3d2310",x"3a210f",x"3a210f",x"38200e",x"3c2311",x"3a2210",x"38200e",x"170f07",x"301c0d",x"311f11",x"372213",x"2d1d11",x"2b1c11",x"422511",x"38200f",x"39200e",x"3b220f",x"3b220f",x"381f0e",x"331c0c",x"371f0e",x"311b0b",x"36200e",x"38200f",x"3c220f",x"160e07",x"1b1108",x"412e21",x"33261e",x"1a140d",x"27160a",x"27160a",x"3b2415",x"262019",x"231509",x"25150a",x"29180b",x"3a200e",x"483224",x"483224"),
(x"5c4c3e",x"5c4c3e",x"58493b",x"544638",x"534233",x"544232",x"4e3c2d",x"564230",x"55412f",x"58422e",x"5f4a35",x"5e4836",x"604c3a",x"5f4c3a",x"5d4734",x"5c4735",x"5e4835",x"614c37",x"664f3b",x"654d37",x"654e38",x"67503b",x"644c37",x"67503b",x"6b523d",x"674e3a",x"664f3a",x"664f3b",x"6a513c",x"67503b",x"69523c",x"654f3b",x"69513b",x"6d563f",x"69533d",x"68543d",x"6e553e",x"70573f",x"6b513b",x"6c533b",x"6a513b",x"6a5138",x"6e563c",x"6d523a",x"694f39",x"6a5038",x"634a33",x"664c35",x"6c5038",x"6a4f36",x"664b34",x"604831",x"654a32",x"6a5138",x"664b35",x"674d35",x"684e37",x"664d37",x"674d36",x"644c36",x"654e38",x"634c38",x"654e3a",x"644d39",x"614b38",x"664f3c",x"66513d",x"624f3b",x"654e3a",x"614a36",x"5e4735",x"5e4937",x"5e4836",x"5e4837",x"5c4937",x"584534",x"5a4634",x"594533",x"544030",x"523f2f",x"544233",x"574535",x"493c2f",x"493c2f",x"150e07",x"4c3825",x"412f1e",x"3f2d1d",x"3f2d1c",x"3c2a1b",x"3c2b1c",x"221a11",x"59422c",x"4a3625",x"423021",x"3c2c1d",x"3d2c1c",x"3f2e1e",x"3c2c1d",x"3c2e1e",x"362719",x"402e1e",x"3d2b1c",x"412f1f",x"3c2b1c",x"3d2b1c",x"38291a",x"3c2b1c",x"3f2d1d",x"3a291a",x"382718",x"3a2819",x"3b2a1b",x"3a2a1a",x"342416",x"342415",x"382718",x"3a2a1a",x"342516",x"362618",x"342416",x"352517",x"2f2013",x"2f2114",x"322316",x"332416",x"352517",x"2d1f13",x"2e2013",x"302215",x"2d2114",x"2f2316",x"2f2215",x"2c1f13",x"2c1f12",x"2d2014",x"271b10",x"261a10",x"251a0f",x"24190f",x"24190f",x"23180e",x"271c12",x"211a14",x"382b1f",x"5d4530",x"413023",x"413121",x"443221",x"433121",x"402e1d",x"422f1e",x"45311f",x"422f1e",x"422f1d",x"473221",x"463220",x"412f1e",x"4a3522",x"3f2d1c",x"422f1e",x"453221",x"433221",x"453624",x"493624",x"453221",x"3f2d1d",x"453221",x"412f1f",x"382819",x"413020",x"402e1e",x"3f2d1d",x"3d2b1b",x"3a2819",x"372718",x"3b2a1b",x"392819",x"322316",x"2d2012",x"322315",x"342618",x"2f2114",x"302214",x"2b1e12",x"291c11",x"291c10",x"261a0f",x"2a1d11",x"21170d",x"2a1d11",x"20160c",x"21170d",x"23190f",x"231a10",x"231a0f",x"251b10",x"251b12",x"241a11",x"251b12",x"231910",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b211a",x"2b211a",x"2e2118",x"33241a",x"352419",x"341f10",x"341f10",x"150e07",x"150e07",x"150e07",x"1d1108",x"23150a",x"25160a",x"3d220e",x"341e0d",x"341d0d",x"321c0d",x"2d1a0b",x"2e1b0c",x"321d0d",x"341e0e",x"321d0e",x"37200f",x"3e2411",x"351f0f",x"351f0f",x"321e0e",x"351f0f",x"3d2411",x"3f2512",x"351f0f",x"3d2411",x"38200f",x"3e2512",x"3d2411",x"392110",x"3d2411",x"3d2411",x"3d2411",x"392110",x"361f0f",x"361f0e",x"39210f",x"3d2410",x"38200f",x"361e0e",x"311c0c",x"38200e",x"351e0d",x"39210f",x"3c2310",x"3a2110",x"3c2310",x"3a2210",x"3a210f",x"371e0d",x"361f0e",x"381f0e",x"371f0e",x"351e0d",x"37200f",x"402511",x"3d2411",x"402512",x"3e2411",x"3e2411",x"3f2512",x"3a210f",x"341d0d",x"39200e",x"180f08",x"2a180b",x"26160a",x"301d0e",x"2a190d",x"2a1a0d",x"472a15",x"371f0f",x"2e190b",x"2b180b",x"331c0c",x"3c2310",x"3f2410",x"3a210f",x"3f2511",x"24150a",x"28170b",x"231409",x"19120c",x"17110a",x"18110a",x"1e1208",x"231409",x"231409",x"2b170a",x"271609",x"2c180a",x"2d190b",x"321c0c",x"311c0c",x"311c0c",x"311b0c",x"321c0c",x"321c0c",x"331c0d",x"321c0c",x"311b0c",x"361e0d",x"311c0c",x"321c0c",x"321c0c",x"351d0d",x"39200f",x"3a2210",x"3e2411",x"3a210f",x"3c220f",x"39200f",x"351e0e",x"381f0e",x"3a210f",x"3a2110",x"39200f",x"3b2311",x"3f2512",x"3f2511",x"3e2511",x"412712",x"422712",x"3f2512",x"3d2411",x"442813",x"3f2512",x"3f2512",x"3d2411",x"402512",x"3f2512",x"36200f",x"3c2311",x"3e2411",x"3e2511",x"3c2310",x"3e2411",x"3a220f",x"3a210f",x"3c2310",x"39200f",x"37200f",x"3b210f",x"170f07",x"28180c",x"342011",x"352012",x"2c1d11",x"26190f",x"462712",x"39200e",x"331d0d",x"38200e",x"381f0e",x"37200e",x"341d0d",x"381f0e",x"321b0b",x"3c2310",x"3e2411",x"3f2511",x"160e07",x"1d1108",x"3f2b1e",x"32261d",x"19120b",x"26160a",x"27160a",x"3c2415",x"272019",x"25150a",x"26160a",x"2f1b0d",x"3d220e",x"462e1f",x"462e1f"),
(x"57483b",x"57483b",x"554638",x"544436",x"564435",x"524131",x"564231",x"523f2e",x"56402e",x"52402f",x"594432",x"564231",x"614c3a",x"5f4a37",x"5d4835",x"5e4a37",x"624c38",x"634c38",x"674d38",x"6c533d",x"694f39",x"644c38",x"634a34",x"674e39",x"654e39",x"644e39",x"644d38",x"684e38",x"6c533c",x"654c36",x"6b523d",x"6a513c",x"6d543e",x"6c533d",x"6c543f",x"674f3a",x"69513c",x"6a513a",x"6b523a",x"6b523b",x"634c35",x"674f39",x"674f38",x"694f38",x"69503a",x"67503b",x"684f39",x"6a513a",x"664d37",x"664d35",x"664c36",x"6a4f35",x"674d35",x"614831",x"644a33",x"674c35",x"614730",x"674d35",x"684e37",x"644b36",x"674e39",x"624b36",x"634c38",x"624a36",x"624c37",x"624b37",x"644c39",x"614a37",x"644d38",x"5d4733",x"614a36",x"5e4936",x"5b4835",x"604c3a",x"594734",x"564333",x"5a4636",x"564332",x"564231",x"554231",x"554333",x"564435",x"4b3d31",x"4b3d31",x"150e07",x"45311f",x"3e2b1b",x"3a2919",x"3e2c1c",x"3c2a1b",x"3b2a1b",x"1b150e",x"624931",x"453222",x"3d2d1e",x"38281b",x"42301f",x"3f2d1d",x"3e2d1d",x"322316",x"3d2c1d",x"3a2819",x"3f2d1d",x"3f2d1e",x"3a2a1b",x"3f2f1f",x"3d2b1c",x"3b2a1b",x"3e2c1d",x"3d2c1c",x"3d2c1c",x"3d2c1d",x"3b2a1a",x"3f2d1d",x"3b2a1a",x"3c2b1b",x"39281a",x"342416",x"362517",x"362617",x"342416",x"332416",x"362517",x"2e2013",x"302215",x"2d1f12",x"322316",x"2f2114",x"2e2013",x"302214",x"2a1e12",x"2d2013",x"2b1e12",x"2a1d11",x"2a1d11",x"261b10",x"2a1e12",x"261b10",x"23190e",x"23180e",x"24190f",x"24190e",x"271c12",x"201912",x"35291e",x"5b442f",x"493727",x"4d3a29",x"463424",x"422f1d",x"3c2a1b",x"3e2b1b",x"412e1d",x"3f2c1c",x"432f1e",x"3f2c1c",x"453220",x"402d1c",x"43301f",x"412e1d",x"453220",x"422f1e",x"412f1f",x"43301f",x"443120",x"3f2c1c",x"453220",x"443120",x"3d2c1c",x"3f2e1e",x"3b2a1b",x"3d2b1c",x"3d2b1c",x"3c2b1b",x"3d2c1c",x"3b2a1b",x"3b2a1a",x"342517",x"352617",x"362718",x"352617",x"302214",x"302114",x"312214",x"2c1f12",x"2a1d11",x"281b10",x"2a1d11",x"2a1d11",x"25190e",x"261a0f",x"21160c",x"21170d",x"23190f",x"23190f",x"23180f",x"251a11",x"23190f",x"241a10",x"241a11",x"211910",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291f17",x"291f17",x"2f2117",x"302117",x"342418",x"331f11",x"331f11",x"160e07",x"150e07",x"150e07",x"1d1208",x"25150a",x"1e1209",x"3b210f",x"37200f",x"361f0e",x"311c0c",x"361e0d",x"371f0e",x"361f0f",x"36200f",x"2b190c",x"37200f",x"37200f",x"361e0e",x"29180b",x"36200f",x"3b2310",x"392110",x"38200f",x"331e0e",x"3a2110",x"37200f",x"3d2411",x"3e2411",x"3e2512",x"402612",x"3d2311",x"3c2311",x"3f2512",x"3a2210",x"3c2311",x"3a2210",x"39210f",x"351d0d",x"351e0d",x"3c2311",x"3e2411",x"3f2411",x"38200f",x"39210f",x"38200f",x"3e2411",x"3f2411",x"3e2411",x"402612",x"3d2411",x"3c2210",x"402612",x"3b2210",x"3a2210",x"3d2311",x"402512",x"402511",x"3f2411",x"3d2410",x"3e2411",x"351e0d",x"3a2210",x"3b2211",x"180f08",x"26170a",x"2e1a0c",x"331d0f",x"25170b",x"29180c",x"472a14",x"311c0c",x"2d190b",x"29170a",x"3a220f",x"38200f",x"3d2310",x"3b210f",x"3b2210",x"26160a",x"2b190b",x"241409",x"1a130c",x"171009",x"171009",x"201309",x"28170a",x"231509",x"321d0d",x"2f1b0c",x"2c190b",x"321c0d",x"361f0e",x"361f0e",x"361f0e",x"37200f",x"361f0e",x"321c0c",x"331c0c",x"341d0c",x"301a0b",x"351e0d",x"38200f",x"3f2411",x"392110",x"39210f",x"3c2311",x"3b2210",x"3d2310",x"3d2411",x"3d2411",x"3b2210",x"361e0d",x"391f0e",x"3a210f",x"3d2311",x"402612",x"3f2411",x"3c2310",x"39210f",x"3a210f",x"3c2310",x"3e2411",x"3f2512",x"3e2512",x"3e2411",x"3b2210",x"3e2511",x"3c2311",x"3c2311",x"3d2311",x"412713",x"3d2411",x"412612",x"3a2210",x"3d2311",x"422713",x"422712",x"3e2411",x"402512",x"3a200f",x"331c0c",x"402512",x"170f07",x"2f1d0e",x"311e10",x"342011",x"2e1d11",x"2b1c10",x"482a15",x"371f0e",x"39200f",x"361e0d",x"3a210f",x"38200f",x"341d0d",x"39200e",x"311b0b",x"3a210f",x"38210f",x"3c210f",x"170f07",x"1e1209",x"3d2a1d",x"2f231a",x"19120b",x"241509",x"25150a",x"351f10",x"1e1811",x"251509",x"27160a",x"2c1a0c",x"3b210e",x"452f21",x"452f21"),
(x"58493c",x"58493c",x"5a493a",x"564435",x"4e3d2d",x"524031",x"523f2f",x"58422f",x"4f3c2c",x"594330",x"5c4633",x"604a38",x"654f3a",x"604b38",x"614b37",x"624b38",x"664e39",x"664e3a",x"654e38",x"6a523b",x"69503b",x"674f39",x"654d38",x"695039",x"684e38",x"6a513b",x"6a5037",x"6e543b",x"70543c",x"72573f",x"6c513b",x"694f38",x"69513c",x"674f39",x"6c533e",x"6a513b",x"694f3a",x"6b523c",x"674e39",x"6d523c",x"6c5139",x"6d543b",x"6a5039",x"684f38",x"6f543d",x"674e35",x"624c36",x"664c35",x"654d37",x"674e36",x"634b35",x"6a5037",x"694e36",x"684e36",x"664c35",x"674c35",x"684e36",x"674e37",x"664c36",x"664d38",x"664d37",x"6a503a",x"644c37",x"634a36",x"664e39",x"604936",x"644d39",x"604a37",x"5e4834",x"604a36",x"5a4432",x"5d4935",x"5f4836",x"5d4936",x"5b4836",x"594534",x"594432",x"584432",x"584433",x"584332",x"554332",x"594636",x"4a3d30",x"4a3d30",x"150e07",x"473320",x"3f2d1c",x"3e2c1b",x"3d2a1b",x"3d2b1b",x"3d2b1c",x"1b150e",x"604731",x"4c3827",x"3b2b1c",x"3c2c1d",x"422f1f",x"3b2a1b",x"3f2d1d",x"39281a",x"422f1e",x"3a2a1b",x"382718",x"402e1e",x"3c2a1b",x"3f2d1d",x"402f1e",x"3c2a1b",x"3d2c1c",x"3c2a1b",x"3b2a1a",x"3a281a",x"3a291a",x"412f1e",x"3b2a1b",x"3c2b1b",x"3b2a1a",x"3a291a",x"382718",x"342416",x"342416",x"362617",x"362618",x"372719",x"362719",x"352618",x"312215",x"2e2013",x"322316",x"2d2013",x"2d2014",x"2b1e12",x"251a0f",x"2c1f13",x"271b10",x"2a1d12",x"2a1d11",x"2d2013",x"24190f",x"24190f",x"24190f",x"24190e",x"23180f",x"1e1811",x"372a1d",x"59422e",x"473526",x"4b3827",x"473423",x"3d2b1c",x"44301e",x"412e1d",x"45301f",x"402e1d",x"422f1e",x"453220",x"42301f",x"4b3724",x"46311f",x"44311f",x"412e1e",x"412f1e",x"443120",x"412e1e",x"45311f",x"42301f",x"3d2b1b",x"412f1f",x"412f1e",x"453221",x"42301f",x"3b2a1b",x"3b2a1b",x"3d2b1c",x"3d2b1b",x"3a281a",x"392819",x"392819",x"3a291a",x"3a2a1a",x"362617",x"332416",x"322315",x"312214",x"2c1f12",x"2c1e12",x"2c1f12",x"2a1e12",x"24190e",x"2c1f13",x"251a0f",x"21170d",x"241a10",x"241910",x"271c11",x"241911",x"231910",x"271c12",x"221910",x"241a11",x"21180f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a2018",x"2a2018",x"2f2218",x"312318",x"342217",x"361f10",x"361f10",x"160e07",x"150e07",x"150e07",x"150e07",x"1f1209",x"231509",x"3c220f",x"321d0d",x"331d0d",x"321c0c",x"36200e",x"311c0c",x"301b0c",x"2d1a0b",x"2f1b0c",x"341e0d",x"37200f",x"37200f",x"37200f",x"3c2310",x"341e0e",x"331d0d",x"38200f",x"3a2210",x"3b2311",x"3c2411",x"392110",x"2d190b",x"351e0e",x"3b2310",x"392110",x"351f0e",x"3f2511",x"3a220f",x"38200f",x"351d0d",x"351d0d",x"371f0e",x"351d0d",x"381f0e",x"381f0e",x"391f0e",x"3a200e",x"3b220f",x"3a210f",x"3b210f",x"371f0e",x"361e0d",x"361e0d",x"38200f",x"39210f",x"371f0e",x"331c0c",x"341d0c",x"331c0d",x"3a220f",x"3a210f",x"39210f",x"3a220f",x"3b2210",x"3d2310",x"392110",x"3a210f",x"191008",x"26160a",x"2c1a0d",x"2f1c0d",x"2c1b0d",x"291a0d",x"3d2211",x"351d0e",x"301b0c",x"2c190b",x"361f0e",x"361f0e",x"3a210f",x"412612",x"3a210f",x"26160a",x"2c1a0c",x"251509",x"17110a",x"171009",x"150e07",x"211309",x"24150a",x"231509",x"321c0c",x"2d190b",x"2a170a",x"27160a",x"2e190b",x"311b0c",x"341d0d",x"351e0d",x"341d0d",x"37200f",x"36200f",x"3d2411",x"3a210f",x"39210f",x"3c2310",x"39210f",x"38200e",x"361f0d",x"361e0d",x"341d0d",x"361e0d",x"38200e",x"3a210f",x"371f0e",x"38200e",x"3b2210",x"38200f",x"39200f",x"321c0d",x"3a200f",x"38200f",x"38200f",x"3b2210",x"3d2310",x"3c2310",x"3b2210",x"3b2210",x"3c2310",x"3e2511",x"3f2512",x"3f2512",x"3d2411",x"361e0e",x"321b0c",x"3a2210",x"3d2411",x"3b2210",x"3e2411",x"3a2210",x"3a210f",x"381f0e",x"361e0d",x"321c0c",x"3a200e",x"39200e",x"160f07",x"29170a",x"2e1b0d",x"311d0f",x"2c1b0f",x"28190f",x"492a15",x"3a210f",x"361e0d",x"3d2310",x"38200e",x"351d0d",x"311c0c",x"2c190b",x"351d0d",x"371f0e",x"371f0f",x"371e0d",x"180f08",x"1e1209",x"3e2c1f",x"261c13",x"171009",x"231409",x"24150a",x"382110",x"231c15",x"25150a",x"27170a",x"2e1b0d",x"3d220f",x"4b3426",x"4b3426"),
(x"584839",x"584839",x"5c4b3b",x"524031",x"554131",x"544232",x"564232",x"56412e",x"58422f",x"594332",x"574331",x"5c4633",x"614b37",x"624d3a",x"5e4835",x"604a37",x"634d39",x"614b37",x"684f3c",x"624b37",x"6a513a",x"69503a",x"634c36",x"644c36",x"644d38",x"674e38",x"674e38",x"6d523a",x"6a5036",x"6e543c",x"6d533c",x"6c513a",x"6a513a",x"6b523b",x"6c533e",x"6b513b",x"6e543b",x"69503a",x"72563e",x"6d523a",x"6d523a",x"71543b",x"6e523b",x"6a4f37",x"6c523a",x"6a513a",x"644d39",x"684f38",x"695038",x"634b34",x"634833",x"644b35",x"684d36",x"664c35",x"604732",x"614933",x"614833",x"684e36",x"634a34",x"674d38",x"634b36",x"664d38",x"644b36",x"624a35",x"684f39",x"654d39",x"674f3a",x"634b37",x"644c38",x"634c38",x"644c36",x"5c4632",x"5f4a36",x"5e4835",x"594331",x"594534",x"5a4534",x"584332",x"534130",x"544031",x"554332",x"5a4736",x"4d3f33",x"4d3f33",x"150e07",x"402d1c",x"372718",x"382718",x"392819",x"3a2819",x"382819",x"1c150e",x"59402b",x"473523",x"3d2d1e",x"3e2d1e",x"402e1e",x"463221",x"42301f",x"3c2b1c",x"3d2c1c",x"3f2d1d",x"3f2d1d",x"412f1e",x"3f2d1d",x"423020",x"402d1d",x"3d2b1c",x"3d2b1c",x"3e2d1d",x"3e2c1c",x"3e2c1c",x"3d2b1c",x"3a2919",x"3a2919",x"3c2a1a",x"382718",x"382718",x"352516",x"332315",x"312214",x"352517",x"322315",x"322316",x"332416",x"2f2114",x"342517",x"2f2114",x"302215",x"302215",x"2f2115",x"2c1f13",x"2e2014",x"2d2014",x"2e2014",x"261a0f",x"2b1e12",x"2b1e12",x"23180e",x"24190e",x"24190e",x"271b10",x"241a10",x"1d160f",x"36291c",x"563f2c",x"463324",x"443222",x"433121",x"412e1e",x"3f2d1c",x"402d1b",x"3f2d1c",x"422f1e",x"3d2b1b",x"402e1d",x"3f2c1c",x"453220",x"44311f",x"432f1f",x"42301f",x"463221",x"483422",x"473322",x"453220",x"463221",x"473422",x"43301f",x"433120",x"433120",x"402e1d",x"3d2b1c",x"3a291a",x"3d2c1c",x"3c2b1b",x"3c2a1a",x"3a291a",x"392818",x"392818",x"372617",x"332315",x"312215",x"2f2114",x"2f2013",x"2e2013",x"2b1e12",x"2a1d11",x"2a1d11",x"251a0f",x"23180e",x"261a0f",x"261a0f",x"261b10",x"261b11",x"251b11",x"271c13",x"241a11",x"251a11",x"251b11",x"21180f",x"221910",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281e16",x"281e16",x"302219",x"302117",x"332216",x"351e0e",x"351e0e",x"160e07",x"150e07",x"150e07",x"1d1108",x"1c1108",x"170f07",x"381f0d",x"2f1b0c",x"321c0d",x"2f1b0c",x"321d0d",x"321d0d",x"2d1a0b",x"2f1b0c",x"301b0c",x"321c0d",x"38200f",x"351e0d",x"341d0d",x"351e0e",x"351e0d",x"331d0d",x"37200f",x"361f0e",x"38200f",x"38200e",x"3a2210",x"382110",x"36200f",x"39210f",x"3a2210",x"38200f",x"38200f",x"3a210f",x"39200f",x"3d2311",x"3d2310",x"341d0d",x"301a0b",x"2d190a",x"311a0b",x"381f0e",x"3c2310",x"38200e",x"351e0d",x"361e0d",x"331c0c",x"311b0b",x"341d0c",x"351d0d",x"331c0d",x"371f0e",x"381f0e",x"3a210f",x"38200f",x"361f0e",x"371f0e",x"371f0e",x"3b220f",x"3b2210",x"3d2310",x"3c220f",x"3a200f",x"150e07",x"26160a",x"2c1a0d",x"2e1b0d",x"28180c",x"26170b",x"3e2311",x"341c0e",x"2e1a0b",x"2c190b",x"341d0d",x"311c0c",x"38200f",x"3e2511",x"361e0e",x"27170a",x"2d1a0c",x"261609",x"171009",x"17100a",x"150e07",x"1d1208",x"241509",x"231409",x"2d190a",x"321c0c",x"321c0c",x"301c0d",x"311d0d",x"331d0d",x"341e0d",x"341d0d",x"341d0d",x"361f0e",x"39200e",x"3a210f",x"371f0e",x"321c0c",x"331c0c",x"3a210f",x"39210f",x"3d2411",x"3b2210",x"351e0e",x"341d0d",x"311b0c",x"321c0c",x"3a210f",x"3c2310",x"39200f",x"3e2410",x"3a2210",x"38200e",x"37200e",x"3a210f",x"39210f",x"39200e",x"39200f",x"371f0e",x"371f0e",x"39200f",x"3a220f",x"39200f",x"3a2210",x"371f0e",x"361f0e",x"392110",x"3a2210",x"3b2310",x"38210f",x"3a2210",x"3a210f",x"38200e",x"3a210f",x"3b220f",x"3d2311",x"39200e",x"321b0b",x"331b0c",x"160e07",x"26160a",x"321d0f",x"2f1d0f",x"291a0f",x"26180e",x"482a15",x"382010",x"3a210f",x"39200e",x"39210f",x"351d0d",x"361e0d",x"30190b",x"321c0c",x"331d0d",x"351e0d",x"3b210f",x"180f08",x"1f1308",x"3c271a",x"251a11",x"171009",x"231509",x"24150a",x"37200f",x"28221b",x"27170a",x"28170b",x"321d0e",x"3a1f0d",x"483122",x"483122"),
(x"5d4b3c",x"5d4b3c",x"534334",x"514030",x"4a3a2d",x"4f3e2e",x"503d2d",x"56412f",x"57412e",x"594431",x"574230",x"604936",x"5f4a37",x"5e4836",x"634d39",x"614c39",x"664f3b",x"644e3b",x"634c37",x"674f3a",x"6c513a",x"6a503b",x"6b5139",x"6e543d",x"6b5039",x"6f533a",x"6d5139",x"6f553d",x"6d5139",x"6e523a",x"6c5139",x"684f38",x"6b5138",x"6b5038",x"664d38",x"654c36",x"5e4532",x"654c36",x"6a4f37",x"6d5138",x"6a4f37",x"6c4f37",x"6d5139",x"6d5139",x"6c5138",x"6b5038",x"6a4f39",x"664c36",x"674e38",x"644c36",x"664b35",x"614933",x"674e37",x"674d37",x"694d37",x"6d533a",x"634a34",x"634a35",x"694f38",x"694f38",x"654c36",x"624a34",x"644b35",x"654c36",x"644d38",x"634b36",x"5d4735",x"604935",x"57412f",x"5d4834",x"5f4732",x"614934",x"5c4532",x"5e4834",x"574230",x"56412f",x"523f2e",x"534130",x"564331",x"554030",x"544232",x"5c4838",x"504135",x"504135",x"150e07",x"422e1d",x"3c2a1b",x"3f2e1e",x"3b291a",x"3c2a1a",x"3d2c1c",x"1b150e",x"5c432e",x"453323",x"412f20",x"3f2e1e",x"3c2b1b",x"43301f",x"3f2c1c",x"3f2c1c",x"362517",x"362617",x"3c2a1b",x"3f2d1c",x"3a291a",x"3c2a1b",x"402e1e",x"3b2919",x"322316",x"3d2b1b",x"3e2c1c",x"3e2b1c",x"3b2a1b",x"3d2c1c",x"3d2b1b",x"392819",x"3b2a1a",x"382718",x"342416",x"3b2a1b",x"382718",x"362517",x"382719",x"3d2c1c",x"342416",x"342517",x"322316",x"332416",x"332416",x"322316",x"2e1f13",x"2b1d11",x"26190f",x"2a1d11",x"281b10",x"2c1f12",x"25190f",x"251a0f",x"251a0f",x"23180d",x"25190f",x"22170d",x"241a0f",x"1d160f",x"33271c",x"57402c",x"463323",x"423021",x"453322",x"3d2b1c",x"453220",x"402e1e",x"422e1d",x"473220",x"453220",x"42301f",x"412e1d",x"443120",x"442f1e",x"3d2b1c",x"44311f",x"493422",x"44301f",x"422f1d",x"3a2819",x"3f2d1c",x"412d1d",x"432f1e",x"3f2c1c",x"422f1f",x"422f1f",x"412e1d",x"382718",x"382718",x"3b291a",x"3b2a1b",x"3a291a",x"372718",x"382718",x"352517",x"372718",x"342416",x"342416",x"322416",x"312215",x"2c1e12",x"2b1e12",x"2d2013",x"23180e",x"251a0f",x"23180d",x"23180e",x"23180d",x"241a10",x"24190f",x"22180f",x"20180f",x"221910",x"251b12",x"241b11",x"221a11",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"271d15",x"271d15",x"2e2016",x"2f2015",x"362215",x"361f0f",x"361f0f",x"160e07",x"150e07",x"150e07",x"1a1008",x"1a1008",x"180f07",x"3f230f",x"301b0c",x"361e0d",x"331d0d",x"331d0d",x"311b0c",x"311c0c",x"311c0c",x"321c0c",x"351e0d",x"371f0e",x"371f0e",x"39200f",x"351e0d",x"351e0e",x"341d0d",x"351d0d",x"331d0d",x"321c0d",x"381f0e",x"351e0d",x"28170a",x"371f0f",x"3a2210",x"3a2210",x"39200f",x"361f0e",x"3d2311",x"371f0d",x"3c2310",x"39210f",x"351e0e",x"39210f",x"38200f",x"321c0c",x"3a210f",x"361e0d",x"341d0c",x"321b0b",x"2f190b",x"311b0b",x"351d0d",x"341c0c",x"341d0d",x"331c0c",x"331c0c",x"331c0c",x"381f0e",x"3d2310",x"361f0e",x"38200e",x"39200e",x"361e0d",x"331b0b",x"341c0c",x"361d0d",x"321b0b",x"160e07",x"251509",x"29170c",x"28180d",x"26170d",x"28190d",x"3d2413",x"21130b",x"2e1b0d",x"311c0c",x"361e0d",x"301b0c",x"3b2210",x"3d2310",x"38200f",x"28170a",x"2e1b0c",x"28160a",x"171009",x"18110a",x"150e07",x"180f07",x"211309",x"231409",x"2c190b",x"331d0d",x"2e190b",x"341d0d",x"2c180b",x"2f1a0b",x"2e1a0b",x"341e0d",x"331d0d",x"301b0c",x"311c0c",x"321c0d",x"341e0d",x"38200f",x"341e0d",x"3a210f",x"341d0d",x"361e0d",x"3b210f",x"39200e",x"311b0c",x"311c0c",x"311c0c",x"381f0e",x"381f0e",x"38200e",x"3b210f",x"3b210f",x"381f0e",x"371f0e",x"371f0e",x"3b210f",x"3b220f",x"38200e",x"361e0d",x"341d0d",x"351e0d",x"351d0d",x"3b210f",x"371f0e",x"321c0c",x"361e0d",x"341d0d",x"351e0e",x"36200f",x"382110",x"37200f",x"341e0d",x"38200f",x"402511",x"3f2411",x"3c2310",x"3a210f",x"3e2411",x"3a2210",x"150e07",x"27160a",x"2d1b0d",x"2e1b0f",x"26180e",x"25170d",x"472915",x"382010",x"361e0d",x"351d0d",x"3b2210",x"381f0e",x"381f0e",x"2d170a",x"321c0c",x"311b0c",x"371f0e",x"39200f",x"180f08",x"1f1208",x"3d2517",x"2b1e14",x"1a130c",x"241509",x"25160a",x"331c0d",x"2a241d",x"27170a",x"28170b",x"311d0d",x"321a09",x"4a3220",x"4a3220"),
(x"644f3d",x"644f3d",x"524132",x"4b3c2e",x"524132",x"513e2e",x"4e3c2c",x"513d2d",x"58412e",x"59432e",x"584432",x"5e4734",x"614d3b",x"67503d",x"66503d",x"644e3a",x"6a523e",x"664f3b",x"664f3c",x"6d543f",x"6e553f",x"70563f",x"70563f",x"6b513a",x"71543c",x"6f533a",x"74563c",x"6f533a",x"70543a",x"71543a",x"6b5037",x"6d523a",x"6f533b",x"6f523b",x"664b35",x"614833",x"674c36",x"684d37",x"684c36",x"6b5037",x"6e5138",x"6c5036",x"684e36",x"6e5238",x"71543a",x"71553b",x"71563e",x"6e533a",x"6c5139",x"664d36",x"6b5139",x"694e37",x"6b5139",x"73563d",x"6e543a",x"6c5039",x"634a34",x"664d38",x"694f39",x"644c36",x"6a5038",x"654c36",x"684e37",x"634a36",x"674d37",x"654c37",x"5c4532",x"5b4431",x"5f4631",x"614835",x"5d4530",x"5f4832",x"59432f",x"58422f",x"584330",x"594533",x"5b4633",x"574330",x"594534",x"5a4534",x"554231",x"5d4938",x"524336",x"524336",x"150e07",x"463321",x"433020",x"3f2d1d",x"3c2a1b",x"3f2d1d",x"3e2c1d",x"1b140d",x"5d452e",x"453322",x"3f2e1f",x"3c2c1d",x"402d1d",x"3c2a1b",x"382618",x"372617",x"3f2d1c",x"3e2b1c",x"3a2919",x"3c2a1b",x"3b2a1a",x"3c2a1b",x"3e2c1c",x"412f1e",x"3c2b1b",x"3f2d1d",x"3e2c1d",x"402d1d",x"3c2b1b",x"3b2a1b",x"3d2b1c",x"3d2b1c",x"3e2c1d",x"412f1f",x"3e2c1d",x"3a291a",x"382718",x"3c2b1b",x"382719",x"342516",x"342517",x"332416",x"302214",x"2d1f13",x"312215",x"312215",x"2b1d11",x"261a0f",x"2b1e11",x"291c11",x"2a1d11",x"2a1d11",x"271b10",x"25190e",x"271b10",x"261a0f",x"24190e",x"24190e",x"251b11",x"1e1811",x"34271b",x"543e2b",x"483625",x"463424",x"493625",x"4b3725",x"4c3725",x"4a3522",x"483321",x"483422",x"463220",x"3f2c1c",x"3f2d1d",x"453220",x"3f2c1c",x"3d2b1b",x"45311f",x"463220",x"3c2a19",x"3e2a1a",x"402d1d",x"402d1c",x"3f2d1c",x"432f1e",x"402d1c",x"422e1d",x"3d2b1b",x"402e1d",x"443220",x"42301f",x"3e2c1d",x"3c2b1b",x"3e2c1c",x"3b2a1b",x"382819",x"362718",x"39291a",x"3c2b1c",x"342517",x"352517",x"2f2114",x"2e2014",x"2f2114",x"291c11",x"261a0f",x"291c11",x"20160c",x"22170d",x"23180d",x"21170e",x"20160d",x"21180f",x"221910",x"241a11",x"231a11",x"251b12",x"221911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"271d15",x"271d15",x"2d1f15",x"2c1d14",x"352114",x"38200f",x"38200f",x"160e07",x"150e07",x"150e07",x"150e07",x"191008",x"201309",x"371e0d",x"331e0e",x"36200e",x"351e0d",x"361e0e",x"37200f",x"37200f",x"341d0d",x"341e0d",x"3b2210",x"37200f",x"361f0e",x"371f0e",x"3a210f",x"321c0d",x"341d0d",x"321c0c",x"351e0d",x"311c0d",x"39210f",x"38200f",x"301c0d",x"39210f",x"351f0e",x"39210f",x"39210f",x"37200f",x"3c2310",x"39210f",x"39200f",x"3a210f",x"331d0d",x"311c0c",x"361e0e",x"371f0e",x"351e0d",x"351d0d",x"351d0d",x"371f0e",x"331c0c",x"341c0c",x"321b0c",x"331c0c",x"331c0c",x"381f0e",x"371e0d",x"371e0d",x"371f0d",x"371e0d",x"351e0d",x"351e0d",x"3a210f",x"3d230f",x"39200e",x"3a210e",x"3c220f",x"39200e",x"1d1208",x"28170a",x"2b1a0c",x"28190e",x"26180e",x"26170d",x"412716",x"2a170b",x"351e0f",x"2c190b",x"381f0e",x"321c0d",x"36200f",x"3d2311",x"39210f",x"29180b",x"2c1a0c",x"28170a",x"171009",x"17110a",x"150e07",x"150e07",x"1e1208",x"231409",x"2f1a0b",x"2d190b",x"321c0c",x"311b0c",x"341d0d",x"311c0c",x"321c0d",x"341e0d",x"321c0d",x"311c0c",x"331d0d",x"2e1a0b",x"331d0d",x"39200f",x"37200f",x"361e0d",x"2f1a0b",x"351e0d",x"3a210f",x"371f0e",x"351e0d",x"361f0e",x"36200f",x"3d2411",x"402511",x"351e0d",x"3a210f",x"3b2310",x"381f0e",x"38200e",x"3e2411",x"38200f",x"38210f",x"361f0e",x"341d0d",x"331c0d",x"331d0d",x"371f0e",x"341d0d",x"361e0d",x"39200e",x"39200f",x"361f0e",x"38200f",x"37200e",x"38200f",x"37200f",x"39210f",x"37200f",x"361f0f",x"39210f",x"371f0e",x"351f0e",x"351d0d",x"351d0d",x"150e07",x"28170a",x"2a190c",x"2b1a0c",x"25180e",x"24170d",x"482a15",x"3a2211",x"38200e",x"3a210f",x"3a210f",x"3b220f",x"371f0d",x"2c180a",x"311c0c",x"311b0c",x"3a2210",x"3a200e",x"180f08",x"201309",x"3b2619",x"31251c",x"19130c",x"24150a",x"26160a",x"321d0f",x"282019",x"211309",x"2e1b0c",x"331e0e",x"361d0a",x"493221",x"493221"),
(x"6f5744",x"6f5744",x"574535",x"574535",x"544132",x"523f2e",x"55402f",x"54402f",x"57412f",x"5b4532",x"5b4533",x"5b4735",x"604b38",x"66503b",x"654f3b",x"66503a",x"69513d",x"6c5440",x"6d5642",x"745a43",x"705640",x"715740",x"705640",x"745a43",x"765941",x"775a40",x"6e543b",x"70543c",x"70543b",x"6e5237",x"6b5037",x"6c5138",x"6e523a",x"70543b",x"70533a",x"6b4f37",x"6f533b",x"6b5038",x"6d5138",x"6c5037",x"694e34",x"77573a",x"725439",x"70533a",x"6f533a",x"71543b",x"71553c",x"6f533a",x"694f38",x"6d543b",x"6d533b",x"6f553c",x"75583f",x"71563e",x"72563d",x"72563c",x"6d523a",x"6d533b",x"644b36",x"624a33",x"674d36",x"684c34",x"634b33",x"624932",x"684d36",x"684f39",x"654d37",x"614a34",x"624935",x"644a34",x"624832",x"5e4731",x"5a432d",x"5f4734",x"5e4834",x"5a4432",x"564231",x"5d4836",x"5d4836",x"5a4533",x"584432",x"624e3c",x"5a493a",x"5a493a",x"150e07",x"473322",x"433020",x"433121",x"422f1f",x"3f2d1d",x"3e2d1d",x"19130c",x"5d432e",x"473422",x"3d2c1c",x"3f2d1c",x"43301e",x"402d1c",x"3c2a1b",x"3d2b1b",x"412e1e",x"3f2d1c",x"412e1d",x"3e2c1b",x"372618",x"402d1d",x"43311f",x"3d2b1c",x"39281a",x"412e1f",x"3e2c1d",x"3f2d1d",x"3e2c1d",x"423020",x"402f1f",x"453221",x"423020",x"3f2d1d",x"3f2e1e",x"3d2d1e",x"422f1f",x"382819",x"3e2d1d",x"342416",x"332416",x"2d1f12",x"2e2013",x"2d1f12",x"312215",x"2f2114",x"2f2114",x"332416",x"2f2114",x"2a1d11",x"2a1d11",x"291c10",x"271b10",x"291d11",x"261a0f",x"23180e",x"21160d",x"271b10",x"281d12",x"1d160f",x"33271b",x"58412e",x"4d3b29",x"4e3b29",x"4e3a28",x"493624",x"493523",x"4e3927",x"4f3a26",x"483423",x"453221",x"402d1d",x"3d2b1b",x"402d1c",x"3f2d1b",x"422e1d",x"46311f",x"453220",x"483321",x"443120",x"453120",x"412e1d",x"412e1d",x"412d1c",x"3d2b1b",x"493422",x"473221",x"422f1e",x"412e1e",x"433120",x"433020",x"3f2d1d",x"3d2b1c",x"402e1e",x"3f2d1e",x"3c2b1d",x"3c2c1d",x"362618",x"38281a",x"37281a",x"352518",x"2f2115",x"2f2115",x"2b1e12",x"291c10",x"271b0f",x"23180d",x"24180e",x"23180e",x"23180e",x"23180e",x"231910",x"241911",x"241b11",x"241a11",x"231a11",x"221911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"261b12",x"261b12",x"271b12",x"2a1b10",x"311f11",x"371f0e",x"371f0e",x"160e07",x"150e07",x"150e07",x"150e07",x"1f1209",x"1c1108",x"3f230f",x"321c0d",x"361f0e",x"301b0c",x"392110",x"37200f",x"39210f",x"351e0e",x"341e0d",x"361f0e",x"38200f",x"301b0c",x"331c0d",x"351e0d",x"341d0d",x"361f0e",x"3c2311",x"331d0e",x"38200f",x"3d2311",x"39210f",x"2f1b0c",x"341d0d",x"331d0d",x"321c0d",x"341d0d",x"351e0d",x"3a210f",x"341d0d",x"361e0d",x"361f0e",x"38200e",x"361f0e",x"38210f",x"331d0d",x"361e0e",x"3a2210",x"392210",x"3b2310",x"39210f",x"3d2411",x"3b2210",x"3d2311",x"402512",x"402511",x"412512",x"3e2411",x"3d2411",x"3c2311",x"3a2210",x"3d2311",x"3d2311",x"39200f",x"351e0d",x"3d220f",x"381f0e",x"3c210f",x"1c1108",x"29180b",x"311d0f",x"2e1b0e",x"27190e",x"26180c",x"3d2515",x"2c190e",x"392111",x"2b180a",x"311b0b",x"2d190b",x"321d0d",x"3b2210",x"392110",x"29180b",x"2a170b",x"27160a",x"17110a",x"17110a",x"150e07",x"170f07",x"1d1208",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"2a180b",x"2d1c0e",x"2e1c0e",x"23160b",x"1e140b",x"472916",x"372010",x"39200f",x"341d0d",x"412611",x"371f0e",x"321c0c",x"38200f",x"331c0c",x"331d0d",x"38200f",x"371e0c",x"180f07",x"221409",x"3f291b",x"35271e",x"19120b",x"24150a",x"27160a",x"341f10",x"251c15",x"372f27",x"2b180b",x"482a14",x"391f0a",x"5a4434",x"5a4434"),
(x"715a45",x"715a45",x"5a483a",x"554334",x"544234",x"544030",x"533f2e",x"54402f",x"513e2d",x"5b442f",x"594330",x"5a4532",x"5e4837",x"644d38",x"5c4736",x"654e3b",x"674f39",x"6c543f",x"654d38",x"70563f",x"6e533c",x"71563f",x"6e543e",x"6e543d",x"71573f",x"71553d",x"72573e",x"6a5038",x"71543a",x"72553a",x"73563c",x"72553b",x"6e543b",x"6f543b",x"72563b",x"71543a",x"6c5136",x"6c5039",x"6b5038",x"6a4f37",x"674c35",x"6d5136",x"6f5238",x"6c5036",x"6c4f36",x"6f5239",x"684e38",x"6d5036",x"6d5037",x"71543c",x"694f36",x"684d36",x"6b5038",x"705338",x"70523a",x"6b5037",x"694d35",x"664c35",x"695037",x"634a32",x"654b33",x"6e5137",x"674b33",x"664c35",x"684f37",x"6b5139",x"654d36",x"644b36",x"644c36",x"674d37",x"654b35",x"5b442f",x"5a422d",x"5a442f",x"574330",x"574230",x"574230",x"594432",x"564230",x"554130",x"594433",x"5f4a39",x"604e3e",x"604e3e",x"150e07",x"473220",x"3f2c1c",x"3f2c1c",x"3f2d1d",x"3c2b1b",x"3a2a1a",x"19120c",x"60472f",x"473423",x"402e1e",x"463222",x"3f2c1c",x"43301f",x"3b2a1b",x"3c2a1b",x"3d2b1b",x"3b291a",x"3d2b1b",x"3b2919",x"392718",x"3a2819",x"3a2819",x"3a291a",x"3e2c1c",x"3e2c1c",x"382718",x"3c2a1a",x"3f2c1c",x"3f2d1d",x"3c2a1b",x"3c2a1b",x"3e2c1c",x"3e2c1c",x"382718",x"3d2b1c",x"3f2d1d",x"382718",x"362718",x"342415",x"372718",x"332416",x"2f2013",x"2f2114",x"312215",x"362618",x"342516",x"312215",x"2c1e12",x"291c11",x"2c1e12",x"2b1e11",x"271a0f",x"281c10",x"281c10",x"24190e",x"22170d",x"23180d",x"251a11",x"1d160f",x"412f20",x"563f2c",x"463423",x"453221",x"433120",x"4a3522",x"483221",x"453120",x"473321",x"4a3422",x"483422",x"412d1c",x"3f2d1c",x"402d1c",x"43301e",x"43301f",x"422f1e",x"43301f",x"45311f",x"45301f",x"412d1c",x"412e1d",x"402d1c",x"3a2819",x"3c2919",x"3f2d1c",x"402d1c",x"402d1d",x"402d1d",x"412e1d",x"3e2c1c",x"3f2c1c",x"3e2b1b",x"3d2b1c",x"3a2919",x"3a2919",x"3a2919",x"342416",x"312215",x"2d1f13",x"322316",x"2f2114",x"2e2014",x"281c10",x"2b1e12",x"291c10",x"291c10",x"23180e",x"23180e",x"23180e",x"21180e",x"20180f",x"241910",x"241a12",x"241b11",x"211810",x"211810",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"241a12",x"241a12",x"271a11",x"2a1a0f",x"2d1b0e",x"361f0e",x"2d1a0b",x"160e07",x"150e07",x"150e07",x"150e07",x"211409",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"2c190c",x"2c190b",x"2f1c0e",x"27180c",x"21150b",x"21150b",x"402716",x"311d0f",x"331f0f",x"2d1a0d",x"341c0c",x"331c0c",x"301b0c",x"361f0e",x"38210f",x"28180b",x"29170a",x"261609",x"17100a",x"18110a",x"150e07",x"150e07",x"150e07",x"1f1309",x"180f08",x"1b1108",x"150e07",x"1c1108",x"1c1108",x"1d1108",x"170f07",x"190f07",x"170f07",x"180f08",x"150e07",x"1d1108",x"1d1208",x"1a1008",x"150e07",x"150e07",x"191008",x"1e1209",x"201309",x"1b1008",x"211409",x"28170b",x"201309",x"211409",x"26160a",x"26160a",x"1b1108",x"180f08",x"1f1309",x"26160a",x"1e1208",x"1b1008",x"1c1108",x"1d1108",x"231409",x"1d1108",x"25150a",x"201309",x"1e1208",x"1d1208",x"150e07",x"1b1108",x"211409",x"191008",x"1f1309",x"25160a",x"201309",x"1d1208",x"23150a",x"1d1208",x"211409",x"1f1309",x"1b1108",x"1c1108",x"221409",x"2c1a0c",x"2d1b0d",x"2d1b0c",x"23160c",x"1f130a",x"1c120a",x"462814",x"361f0f",x"361f0e",x"331d0d",x"351e0e",x"39210f",x"361f0e",x"3a2210",x"37200f",x"321c0c",x"3c2311",x"341d0d",x"191008",x"231509",x"3e281a",x"31261d",x"1a130c",x"24160a",x"26160a",x"492f1d",x"241a11",x"372f28",x"54341d",x"331d0e",x"502f17",x"482914",x"4a3325"),
(x"6e5743",x"6e5743",x"584638",x"5a4738",x"574535",x"554231",x"584432",x"584331",x"56412f",x"5e4732",x"5d4531",x"634c38",x"5d4734",x"634c38",x"644e39",x"644c39",x"6a503b",x"69513b",x"674e39",x"725740",x"725741",x"6e553f",x"6e543e",x"735942",x"735941",x"75593f",x"72563e",x"71543c",x"705338",x"70523a",x"694f37",x"6f5238",x"72543a",x"73563c",x"795a3e",x"74573c",x"72553b",x"73553b",x"73563b",x"72553a",x"694e37",x"74563d",x"71543a",x"74563a",x"74563c",x"6c5138",x"674d36",x"6e5239",x"694e36",x"6e5138",x"664c35",x"6d5137",x"6e5137",x"71543b",x"70543c",x"6e533a",x"6a4f36",x"6c5036",x"674d37",x"664b33",x"684d35",x"674b31",x"694e35",x"664b32",x"694e37",x"694e36",x"6b513a",x"684e37",x"6b513a",x"694f38",x"694f3a",x"644a33",x"614833",x"5f4833",x"5e4734",x"5c4633",x"574332",x"543f2d",x"594332",x"56412f",x"55412f",x"5b4837",x"614e3e",x"614e3e",x"150e07",x"43301f",x"3e2d1d",x"412f1f",x"402e1e",x"3d2c1c",x"3a291a",x"19120b",x"644931",x"453322",x"3c2b1d",x"38281b",x"3a2819",x"3d2b1b",x"463220",x"412e1e",x"402e1d",x"43301f",x"473321",x"43301f",x"3c2a1b",x"3c2b1b",x"3e2c1d",x"3c2a1b",x"3d2c1c",x"3e2c1c",x"412e1d",x"3d2b1b",x"3b2a1b",x"3e2b1b",x"3b291a",x"3a291a",x"3e2b1c",x"3f2d1d",x"3d2c1d",x"423020",x"3a2a1b",x"3a2a1a",x"3a291a",x"382719",x"342517",x"302215",x"302114",x"2d2013",x"322215",x"322315",x"322316",x"342417",x"2d2013",x"2d2013",x"2e2013",x"2b1e12",x"291c11",x"251a0f",x"261a0f",x"23180e",x"23180e",x"25190f",x"251a10",x"1b150e",x"453322",x"513a28",x"463222",x"4a3725",x"453121",x"443120",x"453221",x"493524",x"4b3724",x"483422",x"483321",x"422f1e",x"412e1d",x"422e1e",x"392719",x"3e2b1b",x"3e2c1c",x"45301f",x"473221",x"473221",x"473321",x"463220",x"463320",x"422f1e",x"3f2d1d",x"43301f",x"443120",x"422f1f",x"443120",x"44301f",x"402d1d",x"3d2b1c",x"3d2b1c",x"3a2919",x"362618",x"3a291a",x"3a2819",x"3a291a",x"372719",x"372819",x"332417",x"302215",x"2e2014",x"2c1e12",x"271b10",x"291c11",x"271b10",x"21160c",x"21170d",x"241a0f",x"241a10",x"241911",x"241a11",x"251b12",x"231a11",x"231a11",x"221911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231810",x"231810",x"2a1a10",x"28180d",x"331f0f",x"2c190b",x"26160a",x"160e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"191008",x"1f1309",x"1f1309",x"191008",x"191008",x"1d1208",x"23150a",x"1e1209",x"1b1108",x"180f08",x"180f08",x"22150a",x"24150a",x"1e1209",x"1e1209",x"24160a",x"26170b",x"28170b",x"1e1208",x"170f07",x"1a1008",x"180f07",x"1e1208",x"1d1108",x"211409",x"201309",x"201309",x"1b1008",x"201309",x"201309",x"211409",x"23150a",x"24150a",x"25150a",x"201309",x"24150a",x"27170b",x"2a190c",x"28180b",x"25160a",x"23150a",x"25160a",x"25160a",x"27170b",x"27170b",x"27170a",x"27170a",x"241509",x"231409",x"27170a",x"29180b",x"221409",x"26160a",x"25150a",x"211309",x"27160a",x"28170a",x"26160a",x"2c190b",x"29170b",x"27170a",x"2b1a0d",x"21150b",x"20150b",x"432a18",x"331e10",x"351f0f",x"2d1b0d",x"351e0d",x"341d0c",x"3a200e",x"39210f",x"351f0e",x"26160a",x"27160a",x"261609",x"17110a",x"17110a",x"150e07",x"150e07",x"170f07",x"1a1008",x"1c1108",x"201308",x"191007",x"1c1108",x"1f1208",x"201208",x"201208",x"1f1208",x"221409",x"1d1108",x"1b1108",x"1d1208",x"231509",x"221409",x"211409",x"211409",x"1e1209",x"1d1208",x"201309",x"26160a",x"2a180b",x"29180b",x"2c190c",x"25160a",x"29180b",x"26160a",x"28170b",x"211409",x"25160a",x"221409",x"28180b",x"2a190b",x"2c1a0c",x"26170b",x"23150a",x"29180b",x"23150a",x"23150a",x"28170b",x"211409",x"251509",x"201309",x"1e1208",x"29180a",x"28170a",x"25160a",x"25150a",x"27170a",x"231509",x"24150a",x"27170a",x"26160a",x"28170b",x"28170b",x"1d1108",x"25150a",x"22150a",x"27170b",x"23150a",x"181009",x"181009",x"3a2110",x"341d0e",x"38200e",x"351d0d",x"3a2110",x"3a210f",x"361f0e",x"38200f",x"38200f",x"331d0d",x"38210f",x"39210f",x"1a1008",x"26160a",x"3f2817",x"2f241b",x"18120b",x"23150a",x"26160a",x"331e10",x"211912",x"351f0f",x"452b18",x"311c0d",x"3a200d",x"452f22",x"452f22"),
(x"6f5845",x"6f5845",x"5a493a",x"5a4737",x"554332",x"574433",x"594533",x"55402e",x"57422f",x"5a4431",x"574331",x"614a35",x"614b38",x"634c37",x"69503c",x"664e39",x"6e553e",x"67503b",x"6e543e",x"765b42",x"71583f",x"735940",x"7a5e46",x"795d45",x"7c6149",x"785c44",x"765941",x"785a42",x"76593f",x"73573d",x"74563b",x"76583d",x"785a3f",x"7a5b3f",x"7a5b3f",x"795a3f",x"74583e",x"75583e",x"76583d",x"705339",x"74563a",x"73563c",x"72543a",x"75583c",x"6f523a",x"72543a",x"74573d",x"71543b",x"71543c",x"70553c",x"70533a",x"6d5239",x"72563c",x"705339",x"77593e",x"72563c",x"795b3f",x"70543b",x"6d5239",x"6e5139",x"6c5036",x"6e5137",x"6f5237",x"6f5238",x"73563b",x"71563c",x"74573e",x"74573f",x"6f543d",x"6f533c",x"6a5038",x"644b34",x"644b34",x"5f4733",x"5d4734",x"5c4532",x"5b4532",x"5b4533",x"5b4633",x"574332",x"554332",x"5f4c3b",x"685443",x"685443",x"150e07",x"43301f",x"433120",x"402e1e",x"423020",x"3e2d1d",x"3c2b1c",x"1d150e",x"6f5238",x"493423",x"402e1f",x"453121",x"42301f",x"453221",x"453221",x"402e1e",x"42301f",x"453221",x"433120",x"432f1e",x"3f2d1c",x"3f2c1c",x"3f2d1c",x"402e1d",x"402d1d",x"422f1f",x"3d2c1c",x"3e2c1c",x"402e1e",x"43301f",x"453220",x"42301f",x"412f1f",x"3e2c1c",x"402e1e",x"402e1e",x"443221",x"412f1f",x"412f1f",x"39291a",x"362718",x"392819",x"362618",x"362618",x"39291a",x"332517",x"342517",x"352518",x"302215",x"2f2115",x"2f2115",x"2a1d11",x"2a1d11",x"2b1d12",x"23180e",x"23180e",x"23180e",x"24190e",x"24190e",x"19130c",x"453222",x"58402d",x"473523",x"4d3927",x"473423",x"483422",x"4e3926",x"4d3825",x"4f3a28",x"443221",x"493524",x"483423",x"473321",x"44301f",x"45311f",x"422f1e",x"473322",x"4b3725",x"483422",x"4e3926",x"4a3523",x"4b3625",x"4b3624",x"422f1e",x"44301f",x"443120",x"453220",x"43301f",x"43301f",x"422f1f",x"443120",x"402d1d",x"402e1e",x"3e2c1d",x"3f2d1d",x"3b2a1b",x"3a2a1b",x"3a2a1a",x"39281a",x"372719",x"38291b",x"362719",x"2d1f13",x"2a1d12",x"2c1f13",x"291c11",x"25190f",x"24180e",x"24190f",x"251b11",x"21180f",x"251b12",x"241a11",x"231a11",x"251c12",x"241b11",x"231911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"22170f",x"22170f",x"27170d",x"2a190e",x"2f1c0d",x"2d1a0c",x"241509",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f07",x"1a1008",x"1a1008",x"1c1108",x"1e1209",x"24150a",x"191008",x"211409",x"1d1208",x"27170a",x"231409",x"1c1108",x"1e1208",x"1e1208",x"241509",x"211309",x"1b1108",x"1b1008",x"1d1108",x"170f07",x"1c1108",x"190f07",x"160e07",x"1c1108",x"1d1108",x"1b1008",x"1f1208",x"1b1008",x"1b1008",x"1b1008",x"1d1108",x"201208",x"1e1208",x"211309",x"26160a",x"221409",x"221409",x"27160a",x"29170b",x"26160a",x"25160a",x"201309",x"29180b",x"27170a",x"25160a",x"25150a",x"27160a",x"231409",x"211309",x"1e1208",x"1c1108",x"201309",x"26160a",x"241509",x"231409",x"25150a",x"241509",x"28170a",x"221409",x"221409",x"191008",x"191008",x"4e2f18",x"311d0f",x"351f0f",x"26180c",x"331c0c",x"351d0d",x"341d0d",x"3a2110",x"361e0d",x"24150a",x"251509",x"2c190b",x"211308",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"160e07",x"150e07",x"1a1008",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"150e07",x"150e07",x"4a2b16",x"361f0f",x"321c0c",x"311b0c",x"331d0d",x"361f0e",x"39210f",x"341d0d",x"3a2210",x"3a2110",x"341d0d",x"3e2411",x"3b210f",x"1b1108",x"26150a",x"372110",x"2d231b",x"1b140e",x"211409",x"25160a",x"50392a",x"231d16",x"3b2312",x"362113",x"2e1b0c",x"361e0d",x"4c3627",x"4c3627"),
(x"665241",x"665241",x"564638",x"554536",x"544233",x"54412f",x"584432",x"584432",x"5b4533",x"5d4734",x"554331",x"614a36",x"634b37",x"664e3a",x"654d37",x"654c37",x"684f38",x"6f533c",x"6f5540",x"745942",x"755b43",x"735943",x"785c43",x"775c44",x"745941",x"735840",x"70563f",x"6d543b",x"6f533b",x"6f5239",x"6e5139",x"6c4f35",x"715439",x"72533a",x"715339",x"76583f",x"795c41",x"72553a",x"77593e",x"77593e",x"785940",x"75583f",x"7b5d42",x"785a40",x"795b41",x"71533a",x"72553a",x"6d5138",x"70543a",x"76583d",x"73563c",x"78593e",x"775a3e",x"75573f",x"795a40",x"7a5b3f",x"6f5137",x"6c5038",x"6b4f35",x"6c5035",x"6b5036",x"674c33",x"684b31",x"6b4d33",x"6b5035",x"684d35",x"6d5239",x"6f543b",x"6c523a",x"6d533c",x"6a503a",x"6b533b",x"695039",x"674e39",x"614a36",x"604936",x"5c4633",x"594331",x"54402f",x"544131",x"574232",x"604c3b",x"655140",x"655140",x"150e07",x"433120",x"423020",x"3d2c1d",x"382718",x"382818",x"362617",x"1e160f",x"674c33",x"443121",x"402f1f",x"382819",x"3f2d1c",x"3d2a1a",x"3f2d1c",x"412f1e",x"412f1f",x"3f2d1d",x"443120",x"453221",x"463221",x"42301f",x"412f1f",x"402e1e",x"4c3725",x"422f1e",x"3c2a1a",x"3e2c1c",x"3e2b1b",x"43301f",x"43301f",x"412f1f",x"3e2d1d",x"453221",x"423020",x"453220",x"392819",x"372718",x"352517",x"332415",x"372718",x"332315",x"312214",x"2d1e12",x"312214",x"2f2013",x"2e2013",x"2f2114",x"302215",x"2f2114",x"302215",x"2e2114",x"2c1f13",x"271b10",x"271b10",x"271b10",x"24190f",x"23180e",x"22170d",x"171009",x"402d1e",x"543d2a",x"473524",x"4d3927",x"4a3624",x"453221",x"4a3623",x"4a3523",x"473220",x"463220",x"432f1e",x"3f2d1c",x"473220",x"402c1b",x"3d2a1a",x"402c1b",x"432f1e",x"432e1d",x"412e1d",x"4a3522",x"473322",x"4a3523",x"483422",x"463221",x"483423",x"473322",x"473322",x"463221",x"4b3624",x"43301f",x"412e1d",x"402d1c",x"3d2a1b",x"412e1e",x"3c2b1c",x"3f2e1e",x"3c2b1c",x"3c2a1b",x"3b2a1b",x"3c2a1b",x"352517",x"322315",x"2d1f12",x"2a1d11",x"281c10",x"25190e",x"25190e",x"20160c",x"23190e",x"22180f",x"241a11",x"261b11",x"241a11",x"241b12",x"221910",x"221a11",x"271d14",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"21160d",x"21160d",x"26180e",x"26170b",x"29180c",x"2b190c",x"201309",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"1d1108",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"150e07",x"1d1208",x"150e07",x"1d1208",x"180f08",x"1e1208",x"150e07",x"150e07",x"180f08",x"170f07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"160e07",x"1c1108",x"180f07",x"180f07",x"190f08",x"191008",x"1a1008",x"191008",x"3e2311",x"301d0f",x"361f10",x"311c0c",x"341d0d",x"341c0d",x"39200e",x"3c2310",x"361e0d",x"211309",x"25150a",x"2c190b",x"1f1208",x"19130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4b2b15",x"331d0e",x"38210f",x"351d0d",x"3c2311",x"38200e",x"392110",x"351d0d",x"3a2110",x"3c2311",x"39200e",x"3a2110",x"3a200e",x"1c1108",x"201309",x"634c3b",x"30251c",x"1c160f",x"1e1208",x"1f1309",x"3a291d",x"201912",x"452a17",x"372112",x"311d0d",x"3e220e",x"3b210f",x"3b210f"),
(x"7f634b",x"7f634b",x"594739",x"594637",x"5a4635",x"584432",x"574331",x"544130",x"5d4735",x"5b4533",x"604a36",x"664f3b",x"674f3a",x"68503b",x"6d533b",x"6b513a",x"71573f",x"70543d",x"73583f",x"785c44",x"775c44",x"7a5d44",x"795e45",x"7a5e46",x"785c45",x"745a42",x"765a41",x"6d533c",x"74563c",x"6f533a",x"74573d",x"7b5c3f",x"775a3f",x"74583f",x"735439",x"78593e",x"7a5c42",x"7b5c42",x"77583e",x"795b3f",x"785a3f",x"785b40",x"795c42",x"7f6145",x"806245",x"7a5c3f",x"7a5d43",x"7a5b3f",x"775a41",x"7b5d44",x"75593f",x"7b5c40",x"7d5f43",x"76593e",x"795c40",x"7a5b3f",x"71543b",x"6d5238",x"705339",x"674b34",x"6a4d34",x"674b32",x"70543a",x"71543a",x"705339",x"74583d",x"70533b",x"75583f",x"75583f",x"72563e",x"6e533c",x"6c513a",x"684f3a",x"654c36",x"674f39",x"67503a",x"684e37",x"5e4734",x"5c4733",x"5f4936",x"5e4936",x"634f3d",x"695544",x"695544",x"150e07",x"493523",x"433120",x"402e1e",x"3d2b1b",x"3a2819",x"392819",x"1d160e",x"644930",x"473422",x"412f20",x"493424",x"402e1d",x"422f1e",x"432f1e",x"412f1e",x"433020",x"3b2a1b",x"453120",x"43301f",x"3e2c1d",x"412f1e",x"443221",x"473423",x"503a27",x"4b3724",x"463321",x"483422",x"493523",x"493523",x"453321",x"433120",x"473422",x"423120",x"433120",x"423020",x"3f2d1c",x"3b291a",x"3d2b1b",x"342415",x"342415",x"332314",x"312214",x"3a281a",x"322316",x"302214",x"322315",x"332416",x"312316",x"2e2014",x"2f2114",x"2c1f13",x"2f2114",x"2a1d11",x"281c11",x"281d11",x"281c11",x"251a0f",x"251a0f",x"171009",x"423020",x"523c2a",x"4c3827",x"4d3927",x"4b3724",x"4b3724",x"4a3624",x"493523",x"4a3522",x"493421",x"483321",x"422d1c",x"422f1c",x"422e1c",x"473220",x"483422",x"45311f",x"473320",x"45301f",x"4b3623",x"4d3826",x"4c3624",x"473221",x"4b3724",x"493423",x"483422",x"4a3624",x"4d3926",x"523c28",x"4d3926",x"4c3725",x"473321",x"4c3724",x"473322",x"443120",x"3f2d1d",x"3d2c1c",x"3b2b1c",x"3c2b1c",x"3d2c1c",x"362617",x"332316",x"322316",x"2a1c11",x"261a0e",x"261a0e",x"281c10",x"21160d",x"241a0f",x"271c11",x"231910",x"271c12",x"251a11",x"251b12",x"231a11",x"231a12",x"231a11",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"20150c",x"20150c",x"25160c",x"29190c",x"2a180c",x"2d190b",x"26160a",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f07",x"180f08",x"180f07",x"180f08",x"180f08",x"180f08",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f08",x"180f08",x"180f08",x"422513",x"2d1b0f",x"351f0f",x"2e1a0c",x"38200e",x"381f0e",x"38200f",x"3b2210",x"361e0e",x"1d1108",x"24150a",x"29180b",x"1e1208",x"1a120c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f07",x"190f08",x"190f08",x"180f08",x"191008",x"180f08",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"4d2c16",x"331e0f",x"3e2411",x"38200f",x"39210f",x"381f0e",x"3d2311",x"371e0e",x"3f2411",x"3f2512",x"361e0d",x"371f0e",x"432712",x"1e1209",x"221409",x"594333",x"2c231b",x"1d160f",x"1b1108",x"1b1108",x"3c2d22",x"211a13",x"432816",x"3a2413",x"321d0e",x"3f230f",x"432b1c",x"432b1c"),
(x"7c614a",x"7c614a",x"564536",x"594839",x"524031",x"544131",x"5b4533",x"594534",x"5b4532",x"614a36",x"604935",x"5e4734",x"624934",x"69513b",x"6a5139",x"694f38",x"6e533d",x"694f39",x"684e38",x"6c523b",x"72563e",x"755942",x"755a43",x"745942",x"6f553e",x"6f5640",x"745941",x"755a41",x"6b513a",x"6d503a",x"74573c",x"6f533a",x"74573d",x"75583e",x"795a41",x"7a5b3f",x"73563d",x"76593f",x"7a5c41",x"785b41",x"785a3f",x"795b3f",x"785a40",x"7a5c41",x"75573c",x"795d43",x"7d5e44",x"74583e",x"785a40",x"70543c",x"70543b",x"71553c",x"76593e",x"775b41",x"75563c",x"71543b",x"6d5137",x"6a4f35",x"6f5238",x"6f5239",x"6b5037",x"694c34",x"6d5139",x"6c5138",x"6c5138",x"72553c",x"6f523a",x"75583f",x"6e523a",x"71563f",x"6f543c",x"6f543d",x"6c523d",x"654d37",x"654c37",x"5f4934",x"5e4834",x"5e4835",x"5c4734",x"594533",x"5f4a37",x"5a4635",x"625141",x"625141",x"150e07",x"412f1e",x"402d1c",x"3a2819",x"372718",x"372617",x"362617",x"1b140e",x"64482f",x"473221",x"473423",x"402e1e",x"3d2b1b",x"402e1d",x"422e1d",x"443120",x"432f1e",x"422f1e",x"483422",x"43301f",x"402e1e",x"443120",x"453220",x"473321",x"412e1d",x"453221",x"412f1f",x"42301f",x"3f2d1d",x"3c2a1b",x"3a2919",x"402d1d",x"453220",x"433120",x"3e2c1c",x"3d2b1b",x"3c2a1a",x"3a2819",x"382718",x"372718",x"352516",x"352416",x"342416",x"372718",x"312215",x"332416",x"302114",x"352517",x"312316",x"2e2013",x"312316",x"2d1f13",x"2a1d12",x"2c1f13",x"2a1d11",x"24180e",x"251a0f",x"271b10",x"271b10",x"171009",x"413120",x"4e3826",x"422f1f",x"453222",x"4b3624",x"493523",x"483321",x"422f1e",x"422f1d",x"402d1c",x"45301f",x"473220",x"412e1d",x"442f1d",x"422e1d",x"422f1d",x"473220",x"4a3422",x"4c3622",x"493522",x"4d3724",x"4c3623",x"4e3926",x"4b3624",x"463221",x"483422",x"4a3522",x"4c3623",x"45311f",x"473322",x"463221",x"463221",x"4d3826",x"412d1d",x"3c2a1a",x"3f2c1c",x"3e2d1d",x"3f2d1d",x"392819",x"332315",x"352516",x"312214",x"302114",x"2e1f13",x"261a0f",x"271a0f",x"271b0f",x"21170d",x"21160e",x"241a11",x"251a11",x"271c12",x"251c12",x"251b12",x"261c13",x"231a11",x"231a11",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f140b",x"1f140b",x"27180c",x"29180d",x"281609",x"2b180a",x"27160a",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"190f08",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"190f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"180f07",x"190f08",x"190f08",x"190f08",x"190f08",x"190f08",x"180f07",x"190f07",x"190f08",x"180f07",x"180f07",x"180f08",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"452813",x"2b1a0d",x"321d0e",x"2b180b",x"39200e",x"38200e",x"3a210f",x"3b2210",x"38200e",x"1c1108",x"211309",x"29180b",x"1d1108",x"311b0c",x"311b0c",x"301b0b",x"351d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f07",x"190f08",x"190f08",x"180f08",x"191008",x"180f08",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e220f",x"452812",x"442611",x"462814",x"4b2a13",x"3a210f",x"3d2310",x"381f0e",x"39210f",x"39200e",x"3e2411",x"39200f",x"3c220f",x"3d2411",x"341d0d",x"39200f",x"3f2410",x"1f1309",x"221409",x"553d2c",x"2f261e",x"1e1711",x"180f08",x"191008",x"3e2d22",x"211a13",x"3f2514",x"372111",x"321d0e",x"412410",x"452b1c",x"452b1c"),
(x"785e47",x"785e47",x"5c4b3d",x"5a493b",x"554333",x"544233",x"594432",x"594432",x"604a36",x"634b37",x"664e39",x"634c37",x"674e38",x"6d533a",x"6e5136",x"6f543c",x"6d5239",x"71573f",x"775a40",x"755a41",x"6f553c",x"745840",x"735941",x"755942",x"785c43",x"735740",x"72553c",x"7c5d44",x"77593e",x"7a5e43",x"795d43",x"6b4f36",x"72563a",x"78593e",x"74573d",x"765a40",x"71543c",x"74573e",x"785a40",x"785940",x"816144",x"7a5c42",x"806146",x"7c5d42",x"75573d",x"785b40",x"775a3f",x"74583d",x"7b5e43",x"765941",x"785b42",x"73583f",x"74583e",x"795a40",x"74583e",x"77583d",x"72563b",x"72533a",x"6d5138",x"77583e",x"72553b",x"755a3f",x"795b41",x"654b32",x"6e5339",x"70543a",x"71553c",x"72563e",x"70543b",x"6f543c",x"6e543d",x"6d543d",x"70543e",x"69503b",x"6c523c",x"684e39",x"624a35",x"614a35",x"5f4935",x"5b4634",x"5e4937",x"634e3d",x"625142",x"625142",x"150e07",x"422f1f",x"402e1d",x"3f2c1c",x"3d2b1c",x"3a2919",x"362517",x"1b130b",x"705238",x"4e3a28",x"4a3625",x"3e2b1a",x"3f2d1b",x"442f1d",x"473322",x"42301f",x"422f1e",x"453120",x"4a3523",x"473221",x"473322",x"433120",x"443221",x"473422",x"43301e",x"473320",x"473321",x"473322",x"493523",x"3f2d1d",x"463221",x"493523",x"412e1e",x"473221",x"422f1e",x"3d2b1b",x"3d2b1c",x"3c2a1b",x"3c2a1a",x"3f2d1d",x"402e1d",x"3e2c1d",x"3f2d1d",x"322314",x"352516",x"322315",x"352517",x"332417",x"352517",x"2e2014",x"2e2014",x"2b1e12",x"2d2014",x"2a1e12",x"281c11",x"25190f",x"23180e",x"261b0f",x"261a0f",x"171009",x"4f3b28",x"58412d",x"4e3a27",x"4b3726",x"4b3623",x"493423",x"4d3724",x"463220",x"473321",x"432f1e",x"412e1c",x"473321",x"493422",x"473322",x"4f3926",x"422f1c",x"432f1d",x"493320",x"4c3624",x"4d3825",x"483321",x"483422",x"4f3a26",x"4c3623",x"503a27",x"4e3926",x"4f3b27",x"4a3523",x"453220",x"4b3623",x"4b3623",x"463221",x"4a3624",x"4a3524",x"493423",x"443221",x"412e1d",x"402e1e",x"3b2a1b",x"382819",x"342517",x"332416",x"312215",x"2b1e12",x"2b1e12",x"2c1f13",x"271b10",x"1f150b",x"23190e",x"24190f",x"271c11",x"241a11",x"241a11",x"241b11",x"231a11",x"221910",x"221a11",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"20140b",x"20140b",x"29190c",x"29170a",x"271509",x"2c180a",x"331c0c",x"361e0c",x"341d0c",x"331c0c",x"422612",x"341d0d",x"3b210f",x"3e230f",x"452712",x"422611",x"412511",x"422510",x"3e220f",x"3f2410",x"3f2511",x"452813",x"412511",x"462712",x"402411",x"3d220f",x"2f1709",x"3d220e",x"422611",x"432712",x"3d230f",x"3e220f",x"3f2410",x"442712",x"412611",x"482a14",x"482a14",x"472914",x"4f2f18",x"442813",x"422611",x"472914",x"402512",x"472914",x"412511",x"3f2410",x"402410",x"3e230f",x"3e2310",x"402511",x"452813",x"432712",x"432712",x"432813",x"3d2411",x"412612",x"452914",x"452813",x"422611",x"432711",x"452812",x"412611",x"3c220f",x"3b210f",x"3a210f",x"3a200f",x"3d2310",x"3f2310",x"412510",x"3c220f",x"412611",x"3f2410",x"331c0c",x"331c0d",x"321c0d",x"361e0f",x"3e2412",x"2e1d0f",x"2f1d0e",x"29170b",x"341e0d",x"371f0e",x"3a210f",x"392110",x"3d2310",x"1c1008",x"211409",x"2a180b",x"2b180b",x"301b0b",x"2a170a",x"2a1709",x"381f0d",x"3c210f",x"341c0c",x"341c0d",x"381f0e",x"361e0d",x"381f0d",x"381f0e",x"3a210e",x"3c220f",x"3b210f",x"3a210f",x"3e2311",x"402611",x"3d2310",x"3d2310",x"38200e",x"3b210f",x"3b210f",x"3e2310",x"3b210f",x"3a200e",x"3c220f",x"39200f",x"432712",x"422611",x"402410",x"3f2410",x"412511",x"402410",x"3f2410",x"3c220f",x"3f2511",x"432712",x"442712",x"422612",x"3f2310",x"3c210f",x"3b200e",x"402311",x"412511",x"442712",x"432612",x"472914",x"432611",x"3b210f",x"3e230f",x"402411",x"3e2410",x"3c220f",x"38200e",x"3e220f",x"3c200e",x"3b200e",x"391f0d",x"391e0c",x"3a200e",x"412510",x"41240f",x"371e0d",x"3a200e",x"3e2311",x"412411",x"351e0d",x"3f2410",x"371e0d",x"3d2310",x"39200e",x"361f0e",x"3d2311",x"3a210f",x"381f0e",x"321b0b",x"3b220f",x"361c0c",x"211409",x"231509",x"523b2b",x"282018",x"1e1711",x"170f07",x"170f07",x"3a2b1f",x"2e271f",x"452915",x"3f2614",x"2f1b0c",x"402310",x"4b311f",x"4b311f"),
(x"6e5843",x"6e5843",x"5b4b3c",x"524234",x"524133",x"513e2e",x"533f2f",x"574331",x"5c4735",x"634b37",x"664d38",x"654d38",x"6a5038",x"6a4f38",x"6f5239",x"6e5339",x"6b5038",x"6e513a",x"6e533c",x"70553e",x"73563d",x"6e533c",x"6f553d",x"6f543d",x"76583f",x"75583f",x"75583f",x"73573e",x"74583f",x"7b5d44",x"6f5339",x"7a5b3f",x"6d5138",x"74553a",x"75573c",x"6c5138",x"6b5039",x"6c4f38",x"6a4f39",x"75583e",x"7b5e43",x"785a40",x"76593f",x"70543c",x"75593f",x"775a41",x"7b5d42",x"71553c",x"76593f",x"6f513a",x"70553d",x"73583f",x"6d543c",x"70543a",x"73563b",x"72553b",x"73553b",x"72563c",x"74563d",x"6f5338",x"73563c",x"73553b",x"6c4f37",x"6e5137",x"694d35",x"6a5036",x"6f5339",x"684d34",x"6d5239",x"6b5038",x"6b513b",x"6a513b",x"6d5640",x"674f3a",x"664c38",x"624a35",x"5d4733",x"5f4834",x"5b4533",x"5b4634",x"5a4736",x"624e3c",x"6e5846",x"6e5846",x"150e07",x"422f1d",x"3f2d1c",x"3b291a",x"3d2b1b",x"3c2a1b",x"362517",x"17110a",x"62482f",x"4f3a27",x"3f2d1b",x"45311f",x"3e2b1a",x"44301d",x"422e1d",x"3a2819",x"3c2a1a",x"3f2c1b",x"432f1e",x"463220",x"463222",x"412e1e",x"453120",x"44301f",x"493522",x"473221",x"483322",x"422f1e",x"43301e",x"412e1d",x"44311f",x"4a3523",x"463220",x"422f1d",x"432f1e",x"402d1c",x"3d2b1b",x"422f1e",x"3f2c1c",x"3f2c1c",x"3e2c1c",x"3c2a1b",x"372716",x"3a2818",x"302113",x"322314",x"322215",x"2d1f13",x"2d1f13",x"2d1f13",x"2d1f13",x"2d1f13",x"2c1f13",x"2b1e12",x"291d11",x"25190f",x"261a0f",x"261a0f",x"261a10",x"19130c",x"473322",x"4e3825",x"453321",x"483423",x"4a3523",x"422f1d",x"483321",x"473220",x"4c3623",x"463221",x"422f1e",x"473220",x"453120",x"473221",x"493320",x"4c3521",x"45311e",x"44301d",x"473220",x"442f1d",x"46311f",x"44311f",x"483321",x"4a3523",x"4c3825",x"4d3824",x"4a3523",x"45311f",x"4c3623",x"4b3623",x"4f3925",x"422f1e",x"44311f",x"432f1e",x"43301f",x"443120",x"402d1d",x"3a2919",x"3a2819",x"382818",x"342416",x"352517",x"322315",x"2c1e12",x"2a1d12",x"291c11",x"271b0f",x"25190e",x"1e140b",x"20170d",x"231910",x"241910",x"241a11",x"231a11",x"241c13",x"241b13",x"231b13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"21140b",x"21140b",x"29190d",x"29170a",x"271509",x"2c180a",x"261509",x"2e190a",x"2c180a",x"321c0c",x"351d0d",x"381f0e",x"3a200e",x"371f0e",x"3a200e",x"3a200e",x"3b200e",x"381f0d",x"38200e",x"3e220f",x"3c210f",x"3c220f",x"402410",x"3e220f",x"361e0d",x"321b0c",x"371f0e",x"39200e",x"3a210f",x"3c210f",x"39200e",x"371f0e",x"371e0d",x"3b210f",x"361e0d",x"361d0d",x"3c210f",x"371e0d",x"361e0d",x"351d0d",x"361e0d",x"391f0d",x"381e0d",x"351d0c",x"341c0c",x"30190b",x"321a0b",x"321b0b",x"351c0d",x"371e0d",x"3a200e",x"3d2210",x"402511",x"3d220f",x"3b200e",x"321a0b",x"3a200e",x"3f2410",x"3e230f",x"3d2411",x"3f2410",x"3b220f",x"3b210f",x"391f0d",x"371e0d",x"381e0d",x"371d0c",x"361d0c",x"371d0d",x"391f0d",x"341d0d",x"3a210e",x"361f0e",x"361f0f",x"382010",x"2f1c0f",x"372012",x"331f10",x"351f0f",x"28170b",x"331d0d",x"341d0d",x"331d0d",x"3d2411",x"3a210f",x"1c1008",x"231509",x"2a180b",x"201308",x"29170a",x"2e1a0c",x"301b0b",x"311b0b",x"321c0c",x"301a0a",x"321c0b",x"341d0c",x"331c0b",x"301a0a",x"371e0c",x"40230f",x"2f190a",x"3b210e",x"351d0c",x"3b210f",x"381f0d",x"361e0d",x"371e0c",x"341c0c",x"301a0b",x"351c0c",x"361e0d",x"361e0d",x"331c0d",x"331d0d",x"321c0d",x"361e0d",x"381f0e",x"3a200e",x"3a210f",x"3e2310",x"3d220f",x"3e2310",x"3f2310",x"3e220f",x"3e230f",x"3d2310",x"321b0c",x"361e0d",x"3c220f",x"39200e",x"3d220f",x"3a200e",x"3e2310",x"3b210f",x"3b210f",x"3c210f",x"391f0e",x"3a200e",x"3b210f",x"3c210e",x"391f0d",x"3c210e",x"3b200e",x"371d0c",x"321b0c",x"2e190b",x"311a0b",x"2e180a",x"2d180a",x"331b0c",x"341c0d",x"341d0d",x"39200e",x"3d2310",x"3b210f",x"3f2410",x"3a210f",x"3a210f",x"371f0e",x"39200f",x"3a2210",x"39200f",x"3a210f",x"291408",x"351e0e",x"402410",x"22150a",x"241509",x"503c2e",x"393129",x"1f1812",x"160e07",x"160e07",x"2b241d",x"2f2720",x"3e2311",x"372111",x"2f1c0d",x"391f0d",x"482d1a",x"482d1a"),
(x"765d48",x"765d48",x"5a493b",x"514234",x"4b3c2d",x"544130",x"5b4432",x"5b4532",x"604935",x"634b36",x"604833",x"604833",x"674d36",x"644a34",x"664c35",x"694e35",x"694e36",x"6c513b",x"6e523b",x"6c513a",x"70553e",x"6f543c",x"664d35",x"6d513a",x"6f553c",x"6e5137",x"6f533a",x"6b5038",x"74563c",x"71543b",x"715438",x"705238",x"6d5036",x"705138",x"74553c",x"6d4f37",x"6e5239",x"73553a",x"74553d",x"74563c",x"75583e",x"75583d",x"71543a",x"795a40",x"72553b",x"71543a",x"70523b",x"70533a",x"74563d",x"74563d",x"74553a",x"72563b",x"71553c",x"6b5038",x"6b5038",x"685037",x"71543b",x"6e5238",x"6e5035",x"6f5238",x"73563c",x"715339",x"6d5038",x"6c5038",x"6b5037",x"674d36",x"6f523b",x"6a4e37",x"6f5239",x"70543b",x"6b513c",x"6b513c",x"69513b",x"604a36",x"604935",x"644b36",x"5c4532",x"584330",x"57412f",x"564332",x"574435",x"614e3e",x"705a48",x"705a48",x"150e07",x"3e2c1c",x"382718",x"382718",x"3c2a1b",x"362617",x"332315",x"171009",x"644930",x"42301f",x"3d2c1b",x"3f2c1b",x"422d1c",x"3f2c1b",x"432f1e",x"402d1c",x"3c2a1a",x"45301f",x"473220",x"4a3522",x"43301f",x"3f2d1c",x"412d1d",x"473321",x"422f1e",x"422e1d",x"432f1e",x"3f2c1b",x"44301f",x"432f1e",x"45311f",x"422f1e",x"483422",x"43301e",x"3e2b1b",x"3c2a1a",x"3c2a1b",x"3c2a1a",x"3a2819",x"3b291a",x"3e2c1c",x"3d2b1b",x"342315",x"312214",x"322214",x"322314",x"342416",x"2e2013",x"2f2013",x"312214",x"2e1f13",x"2a1d11",x"2b1e12",x"2a1d11",x"24190e",x"251a0f",x"24190e",x"24180e",x"21170d",x"19120b",x"473422",x"4c3724",x"453121",x"483523",x"473322",x"463220",x"3c2a1a",x"432f1e",x"412d1c",x"402d1c",x"3f2c1b",x"402d1c",x"473220",x"473220",x"422e1c",x"45301d",x"45301d",x"45301d",x"483421",x"422e1d",x"46321f",x"493321",x"4a3421",x"483321",x"4a3522",x"473221",x"46321f",x"493421",x"45301f",x"44301e",x"442f1e",x"412d1c",x"453120",x"422e1d",x"45311f",x"422f1e",x"402e1e",x"3d2b1b",x"362617",x"312215",x"342416",x"342416",x"2d2013",x"2c1e12",x"2e1f13",x"281c10",x"20160c",x"20160c",x"20160c",x"20160d",x"23180f",x"22190f",x"221810",x"241a11",x"241b13",x"241b13",x"211a12",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"22150b",x"22150b",x"2a190d",x"2b1a0d",x"2b180a",x"2d190a",x"251509",x"28160a",x"2d190a",x"351d0d",x"381f0e",x"3a200f",x"3a210f",x"381f0e",x"3a200e",x"39200e",x"351d0d",x"381f0e",x"381f0e",x"371f0e",x"39200e",x"331c0c",x"331c0c",x"39200e",x"39200f",x"331c0c",x"321c0c",x"38200e",x"3a200e",x"3b210f",x"351f0e",x"351d0d",x"351d0d",x"351d0d",x"341d0d",x"311b0b",x"321b0c",x"321b0b",x"331c0c",x"311b0b",x"321b0b",x"2e180b",x"301a0b",x"331b0b",x"301a0b",x"2d1a0b",x"2d180b",x"2f1a0b",x"311b0c",x"371f0e",x"381f0e",x"3a200f",x"311c0c",x"311b0c",x"361e0d",x"331c0c",x"341c0c",x"361d0d",x"371f0d",x"381f0e",x"39200e",x"2e1a0b",x"351e0d",x"3b210f",x"3c210f",x"381f0d",x"3b220f",x"351d0c",x"3c210f",x"391f0e",x"371f0e",x"361e0e",x"371e0d",x"341d0e",x"311c0d",x"2e1b0e",x"2e1c0f",x"301d10",x"2c1b0e",x"26160a",x"321c0d",x"331d0d",x"371f0e",x"3b2311",x"3d2311",x"1e1208",x"25160a",x"2b190b",x"211309",x"241509",x"2c190b",x"2c190b",x"2f1a0b",x"2b180a",x"301b0b",x"321c0b",x"341d0c",x"351d0c",x"321c0b",x"2f1a0a",x"371e0d",x"301b0b",x"381f0e",x"30190b",x"371e0d",x"351d0d",x"361d0c",x"341d0c",x"311b0b",x"2c180a",x"2c180a",x"331c0c",x"341d0d",x"38200e",x"371f0e",x"331d0d",x"311b0c",x"361e0d",x"351d0d",x"331c0c",x"361e0d",x"381f0e",x"3a210f",x"381f0e",x"321b0c",x"341d0c",x"351e0d",x"311c0c",x"2f1a0b",x"381f0e",x"38200e",x"381f0e",x"3a210f",x"3a210f",x"381f0e",x"321c0c",x"3a200e",x"321b0b",x"2e190b",x"2d180b",x"2c190b",x"341c0c",x"301a0b",x"321b0b",x"301a0b",x"311b0b",x"301a0b",x"2e190b",x"2d190b",x"2e1a0b",x"301a0b",x"371f0d",x"381f0e",x"39200e",x"3b210f",x"3d2310",x"3f2411",x"3c220f",x"351e0d",x"371f0e",x"3b2310",x"3d2411",x"3a210f",x"3c2311",x"361e0d",x"3c2310",x"150e07",x"150e07",x"150e07",x"52483e",x"51483e",x"180f07",x"1a1008",x"1c1108",x"50463c",x"50463d",x"3d2211",x"362011",x"301c0d",x"391f0d",x"492c1a",x"492c1a"),
(x"84674f",x"84674f",x"5a4a3d",x"5a4838",x"524132",x"5c4735",x"5e4835",x"5b4532",x"5d4733",x"5f4834",x"614935",x"634a34",x"684e37",x"644b35",x"674c35",x"604732",x"6b503a",x"695039",x"6c5139",x"6f533c",x"6f533b",x"72563e",x"6e523a",x"73553d",x"73553c",x"72553c",x"7c5b40",x"725339",x"75563c",x"765639",x"7e5e42",x"73553a",x"75573c",x"77593f",x"77583e",x"72553c",x"70533b",x"79593f",x"7f5e42",x"795a3e",x"77583e",x"76573c",x"74563b",x"73563c",x"6f5237",x"6e5138",x"6a4e37",x"644b36",x"6f533a",x"6e5137",x"75563b",x"73543c",x"70543d",x"6b503a",x"6f533b",x"6c5139",x"74563d",x"795a3e",x"7a5b3f",x"735439",x"74553b",x"72553a",x"7b5d42",x"6d5138",x"73543c",x"74573e",x"71543a",x"78593d",x"6e5238",x"76593f",x"73573f",x"6c523a",x"6c523c",x"684f3b",x"614935",x"604834",x"5a4430",x"584331",x"55402f",x"554232",x"5b4837",x"604f3f",x"6c5746",x"6c5746",x"150e07",x"3f2c1c",x"3b291a",x"3e2c1b",x"3b2919",x"372718",x"382719",x"191109",x"644930",x"453120",x"453322",x"3c2a1a",x"463120",x"4a3422",x"493321",x"44311f",x"402d1c",x"44311f",x"4a3522",x"473220",x"43301f",x"422e1d",x"412e1d",x"412d1c",x"3f2d1c",x"3e2b1b",x"3c2919",x"402d1c",x"422f1e",x"3f2d1c",x"402d1c",x"422e1d",x"43301f",x"402d1d",x"3f2c1c",x"3e2c1c",x"3a2919",x"3f2c1c",x"3f2c1c",x"3d2a1a",x"3a2819",x"3b2919",x"433020",x"352517",x"3a2919",x"39281a",x"362617",x"372718",x"302114",x"332416",x"2e2013",x"2a1d11",x"2f2114",x"2a1d11",x"2a1d11",x"23180d",x"23180d",x"21160c",x"20160c",x"17110a",x"412f1e",x"4a3522",x"45311f",x"4a3522",x"443120",x"43301f",x"3f2c1c",x"473220",x"463220",x"3f2d1c",x"473221",x"422e1d",x"432f1e",x"46321f",x"523c28",x"422e1d",x"483321",x"4e3824",x"4b3522",x"493421",x"45301f",x"493522",x"513a26",x"493321",x"483321",x"463120",x"473320",x"432f1e",x"412d1c",x"422f1d",x"402c1c",x"412e1d",x"412e1d",x"3e2c1b",x"402d1c",x"422f1d",x"422f1e",x"3b2a1b",x"3a2919",x"342416",x"382718",x"362618",x"342416",x"302113",x"2c1e12",x"271a0f",x"271b10",x"21170d",x"22180e",x"23180f",x"23190f",x"241b11",x"211910",x"231b11",x"241b12",x"201811",x"201911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24160b",x"24160b",x"29190c",x"2c1a0c",x"321c0c",x"301a0b",x"2c190b",x"2d190b",x"2e190b",x"321c0c",x"331c0c",x"321c0c",x"321b0c",x"341c0c",x"3a200f",x"3a210f",x"381f0e",x"361e0d",x"341c0c",x"331b0b",x"30190b",x"2f1a0b",x"371e0d",x"3c220f",x"3c210f",x"351e0d",x"341d0d",x"321c0d",x"3b210f",x"371f0e",x"341d0d",x"311b0c",x"2e190b",x"331c0b",x"301a0b",x"311b0c",x"331c0c",x"341d0c",x"371f0d",x"341d0c",x"341c0c",x"321b0c",x"351d0d",x"361e0d",x"361f0e",x"361e0d",x"2c190b",x"311b0c",x"341d0d",x"351d0d",x"371f0e",x"3a210f",x"381f0e",x"321c0c",x"3b200e",x"361d0d",x"381f0e",x"3c220f",x"381f0e",x"3a210f",x"3a2210",x"37200e",x"3a210f",x"391f0e",x"39200e",x"3e2310",x"3f2410",x"3a200e",x"39200e",x"371e0e",x"3b2210",x"3d2310",x"3c2310",x"3c2211",x"321d0f",x"331d0f",x"301d10",x"321f10",x"331e10",x"24150a",x"351e0d",x"361f0e",x"341d0d",x"412612",x"402511",x"221409",x"26170a",x"29170a",x"27170a",x"2d1a0c",x"27160a",x"261509",x"38200e",x"351e0e",x"331c0c",x"321c0b",x"341c0c",x"371e0d",x"341d0c",x"321c0c",x"39200e",x"351e0d",x"39200e",x"331c0c",x"3a200e",x"3b210e",x"341c0c",x"321b0b",x"351d0c",x"321c0c",x"341d0c",x"341d0c",x"371f0d",x"321c0c",x"2f1a0b",x"301a0b",x"331c0c",x"3a210f",x"371f0e",x"361e0d",x"331c0c",x"341c0c",x"2d180a",x"321b0b",x"311b0c",x"371f0e",x"301b0c",x"341d0d",x"351d0d",x"371f0d",x"381f0e",x"361e0d",x"381f0d",x"341d0d",x"341c0c",x"311a0b",x"301a0b",x"371e0d",x"331d0c",x"321b0c",x"341d0c",x"341d0c",x"361d0c",x"321b0b",x"371e0d",x"391f0e",x"39200f",x"3c220f",x"38200e",x"311b0c",x"361e0d",x"39200e",x"3c210f",x"3b210f",x"3b220f",x"351e0d",x"462814",x"39200f",x"351d0d",x"381f0e",x"38210f",x"3f2411",x"3f2512",x"3d2411",x"361e0d",x"3a2110",x"160e07",x"180f08",x"180f07",x"4d3d31",x"423a31",x"170f07",x"191008",x"1c1108",x"373028",x"4e453b",x"452713",x"382111",x"311d0e",x"361d0c",x"472b18",x"472b18"),
(x"7e624a",x"7e624a",x"58483b",x"584638",x"534131",x"584332",x"5b4534",x"5e4834",x"5f4936",x"624c39",x"644d38",x"634d38",x"6f523a",x"695037",x"6d533c",x"71563d",x"785b40",x"745940",x"6c513a",x"6f523b",x"6f533b",x"71543c",x"73573f",x"77593f",x"75573c",x"76573c",x"78593f",x"78593d",x"7b5c40",x"7a5b3f",x"76573a",x"78593d",x"75563a",x"73543a",x"715238",x"78593e",x"715338",x"705237",x"77593f",x"78593d",x"7c5d42",x"765a3f",x"795b40",x"785c41",x"795c40",x"72563c",x"70533b",x"73573d",x"7f5f43",x"74563c",x"76573d",x"73553c",x"6b5138",x"6f5238",x"72553d",x"76593e",x"74563c",x"77593e",x"7b5b3f",x"7b5c3f",x"795c40",x"7d5e42",x"75563b",x"73563c",x"715339",x"694f38",x"6a4e37",x"71543b",x"6f5239",x"6e523a",x"71553e",x"6a513b",x"705740",x"69513b",x"664f3b",x"5e4a36",x"614a36",x"5d4734",x"5d4836",x"5f4937",x"604c3a",x"62503f",x"6a5747",x"6a5747",x"150e07",x"3e2b1b",x"3c2b1b",x"3c2a1b",x"3a2919",x"342416",x"362617",x"1b130b",x"6a4e34",x"4b3826",x"412e1f",x"463220",x"44301e",x"3f2c1b",x"3e2b1a",x"412e1d",x"3e2b1b",x"432f1e",x"453120",x"473321",x"483422",x"41301f",x"453320",x"443321",x"473322",x"443220",x"43301f",x"463220",x"4a3623",x"453220",x"422f1e",x"3d2b1b",x"402d1c",x"412e1d",x"43301f",x"422f1e",x"432f1e",x"412e1d",x"402d1d",x"3f2d1d",x"412f1d",x"422f1f",x"392819",x"3a2819",x"392718",x"352516",x"342315",x"362617",x"2b1e11",x"2c1e12",x"2e2014",x"2e2013",x"2f2115",x"281d11",x"261a10",x"23190e",x"24190f",x"24190f",x"23180e",x"150e07",x"453220",x"4b3523",x"412f1e",x"45311f",x"412e1c",x"432f1d",x"453220",x"46311f",x"473320",x"45311f",x"473221",x"493422",x"4c3724",x"4d3825",x"483321",x"493321",x"45311e",x"422f1d",x"432e1d",x"493421",x"44301e",x"422f1d",x"453120",x"473321",x"4c3725",x"473523",x"4a3623",x"483523",x"4b3624",x"463221",x"473320",x"4a3523",x"4c3623",x"463220",x"432f1e",x"3f2d1c",x"3d2b1a",x"3b2919",x"3e2c1c",x"3b2a1a",x"3b2a1a",x"362618",x"342416",x"2d2013",x"2e2014",x"2e2114",x"23180d",x"23180d",x"23190f",x"20170d",x"1f160e",x"221a12",x"211911",x"231a12",x"201912",x"201911",x"201911",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24160b",x"24160b",x"2c1a0d",x"2d1b0c",x"321c0e",x"341c0c",x"2d1a0b",x"2b180a",x"321c0c",x"361e0d",x"3a210f",x"38200f",x"381f0e",x"371f0e",x"3b210f",x"341d0d",x"371f0e",x"3e2310",x"3b210f",x"38200e",x"38200e",x"3c220f",x"3c230f",x"381f0e",x"351d0d",x"39200e",x"331d0d",x"381f0e",x"3b210f",x"39200e",x"351d0d",x"331c0c",x"311b0b",x"301a0b",x"301a0b",x"2e190b",x"311b0b",x"321b0c",x"311b0b",x"311b0b",x"311b0b",x"2f190b",x"321b0b",x"331c0c",x"331d0c",x"331c0c",x"351d0d",x"371f0e",x"341d0d",x"2f1a0b",x"31190b",x"331b0b",x"2f1a0b",x"301a0b",x"311a0b",x"301a0b",x"351e0d",x"3b200e",x"381f0e",x"331c0c",x"381f0e",x"3a210e",x"3a200f",x"3a210f",x"3a210f",x"3b210f",x"381f0d",x"361e0d",x"381f0e",x"321c0c",x"371f0e",x"361e0d",x"361f0e",x"3a210f",x"371f0f",x"331d0e",x"332011",x"2f1b0e",x"2d1c0d",x"2c190b",x"341d0d",x"3c2310",x"39200f",x"3d2411",x"3a2110",x"23150a",x"241509",x"211208",x"221409",x"29170a",x"311c0d",x"311d0d",x"311c0d",x"2d190b",x"2e190b",x"2c170a",x"2c180a",x"321c0c",x"38200e",x"341d0d",x"371e0d",x"39200e",x"412511",x"39200e",x"3b200e",x"3c230f",x"3a210f",x"38200e",x"3e2310",x"361d0d",x"321b0b",x"381f0e",x"3b220f",x"351e0e",x"351e0e",x"381f0e",x"361f0d",x"3b2210",x"391f0e",x"3a210f",x"371f0e",x"38200e",x"3a210f",x"381f0e",x"341d0d",x"331c0d",x"301b0c",x"311c0c",x"381f0e",x"361e0d",x"371f0e",x"361f0e",x"371f0e",x"351d0d",x"321c0b",x"321b0c",x"2f1a0b",x"301a0b",x"321b0b",x"2f1a0b",x"2f1a0b",x"311a0b",x"2f1a0b",x"2e190b",x"321b0c",x"361d0d",x"331c0c",x"341d0c",x"311c0c",x"351e0d",x"371f0d",x"351d0d",x"321b0b",x"331b0b",x"321b0b",x"3d2310",x"422712",x"371e0d",x"371f0d",x"3b220f",x"3f2411",x"412512",x"3c2310",x"39210f",x"351d0d",x"3c2310",x"160f07",x"1d1108",x"1b1008",x"443123",x"3e362d",x"180f07",x"1a1008",x"1c1108",x"322821",x"4d443a",x"442713",x"311d0f",x"2e1b0d",x"391f0d",x"472d1b",x"472d1b"),
(x"84664d",x"84664d",x"5c4c3e",x"5d4b3c",x"594637",x"594433",x"604a35",x"624c38",x"664e3b",x"664e39",x"684f3a",x"6a513b",x"674e39",x"695039",x"75583f",x"72563d",x"765940",x"765941",x"785b40",x"73563f",x"71533c",x"73563e",x"74573e",x"785a3f",x"73563c",x"795a3e",x"75573c",x"71543a",x"7a5b3d",x"78583c",x"7a5a3e",x"78583d",x"7b5c40",x"7a5b3f",x"76573a",x"7a5a3d",x"7c5b3e",x"78593d",x"7d5d40",x"7d5e43",x"7e5e43",x"826244",x"785b40",x"785a3f",x"76573d",x"71543a",x"73563a",x"70523a",x"7b5b3e",x"795b40",x"785a3e",x"77583d",x"74563d",x"70543b",x"72543a",x"76583d",x"73563c",x"7a5a3f",x"785a3e",x"76573c",x"7a5c3f",x"785a3e",x"77583c",x"7c5b3f",x"785a3f",x"75583e",x"77573d",x"75573c",x"76583e",x"73573c",x"75583f",x"745942",x"745942",x"6c533b",x"6c523b",x"664e39",x"614935",x"5b4533",x"5d4734",x"574332",x"5d4a39",x"625243",x"6f5b49",x"6f5b49",x"150e07",x"3c2a1a",x"3a2819",x"392818",x"372618",x"382718",x"332416",x"19120b",x"644a32",x"473423",x"453121",x"44311f",x"493321",x"473220",x"483320",x"422e1d",x"43301e",x"46321f",x"453220",x"4c3825",x"483422",x"4b3724",x"473321",x"473321",x"453120",x"412e1d",x"43301f",x"422f1d",x"402d1d",x"432f1e",x"453120",x"402d1c",x"402d1c",x"3d2b1b",x"402d1c",x"402d1c",x"3b291a",x"432f1e",x"3e2b1c",x"362617",x"3c2b1b",x"402d1c",x"3c2a1a",x"3d2b1b",x"3c2a1b",x"3a2819",x"342416",x"332315",x"332416",x"2f2113",x"2a1d11",x"2d2014",x"2d2014",x"2b1e12",x"271b10",x"24190e",x"23180e",x"23180d",x"23180e",x"150e07",x"3e2b1c",x"463220",x"433120",x"463220",x"45311f",x"46311f",x"422f1e",x"45311f",x"43301e",x"483321",x"453120",x"46311f",x"4a3523",x"483320",x"473220",x"483320",x"483321",x"473220",x"483320",x"45301e",x"45311f",x"45311f",x"483422",x"493624",x"4e3926",x"4c3825",x"493523",x"4a3623",x"483321",x"493321",x"493422",x"432f1e",x"483321",x"473220",x"3f2d1c",x"3e2c1b",x"402d1c",x"3b291a",x"3d2b1b",x"3b291a",x"382818",x"382718",x"342416",x"2d1f13",x"2c1f13",x"261a0f",x"281b10",x"23180d",x"241910",x"261b11",x"231910",x"221810",x"231911",x"201811",x"201911",x"201911",x"201811",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24160b",x"24160b",x"2a180c",x"2d1a0d",x"321d0e",x"331c0e",x"2c1a0c",x"321d0d",x"38200f",x"36200f",x"3c2310",x"3b2210",x"3f2411",x"3a2210",x"381f0e",x"381f0d",x"331c0c",x"351e0d",x"371f0d",x"351e0d",x"3d230f",x"361e0d",x"3a200e",x"39200e",x"3f2410",x"381f0e",x"371f0d",x"3b210e",x"3b200e",x"3a200e",x"361e0e",x"381f0e",x"39200f",x"381f0e",x"351d0c",x"361e0d",x"341d0d",x"341c0c",x"371e0d",x"351d0d",x"371f0d",x"361e0d",x"331d0c",x"321b0c",x"321b0c",x"321c0c",x"321c0c",x"381f0e",x"351e0d",x"2e1a0b",x"331c0c",x"331c0c",x"331c0c",x"361e0d",x"351d0c",x"341d0c",x"311b0c",x"331c0c",x"351d0d",x"361f0e",x"311c0c",x"321c0c",x"3a210f",x"3a210f",x"381f0e",x"39200e",x"351e0d",x"321b0c",x"371e0d",x"371e0e",x"361e0d",x"361f0d",x"341d0d",x"381f0e",x"382010",x"361f0f",x"361f0f",x"321d0f",x"2d1a0d",x"2b180b",x"341d0d",x"37200f",x"371f0e",x"3f2512",x"38200f",x"25160a",x"28170b",x"2a180b",x"1e1208",x"211308",x"261509",x"29170a",x"2c190b",x"301b0c",x"361f0e",x"361f0e",x"39210f",x"361e0e",x"38200e",x"38200e",x"39200e",x"39200e",x"3b210e",x"381e0d",x"331c0c",x"331c0c",x"371e0d",x"371f0e",x"3e2310",x"3d2310",x"3b2210",x"3c2311",x"3c2311",x"3b2210",x"341d0d",x"3a2210",x"3a210f",x"3a200e",x"391f0d",x"371e0d",x"39200e",x"38200e",x"381f0e",x"39200e",x"351d0d",x"381f0e",x"371f0e",x"371f0e",x"341d0c",x"371f0e",x"381f0e",x"331d0d",x"351d0d",x"381f0e",x"3a210f",x"39200e",x"341d0d",x"351d0d",x"361e0d",x"331d0c",x"361d0d",x"351d0d",x"301a0b",x"351d0d",x"351e0d",x"321c0c",x"361e0d",x"321c0c",x"371f0d",x"341d0d",x"381f0e",x"381f0e",x"3a200e",x"361e0d",x"351d0c",x"3d230f",x"3e2411",x"351d0d",x"3a210f",x"3c2310",x"3a210f",x"3c2310",x"3e2411",x"3e2411",x"331c0c",x"39210f",x"170f07",x"211309",x"1f1208",x"412d21",x"383129",x"180f08",x"1a1008",x"1c1108",x"32271f",x"4d443b",x"3e2311",x"311c0d",x"29180b",x"381f0d",x"472f1f",x"472f1f"),
(x"82664e",x"82664e",x"594a3c",x"5a4b3d",x"534234",x"524031",x"5b4735",x"624b37",x"614a36",x"6c533c",x"69513b",x"6a503b",x"70553e",x"73573f",x"765941",x"785d45",x"7d6047",x"71543d",x"74573f",x"74583f",x"76593f",x"785a40",x"775a3f",x"74573e",x"74573c",x"72553b",x"76573d",x"785a3e",x"75583d",x"7c5b3f",x"79593d",x"77573c",x"7c5d3f",x"7b5a3e",x"7d5b3f",x"74573a",x"715137",x"735439",x"745439",x"7c5c3f",x"7b5b40",x"7e5e41",x"7b5c41",x"74563c",x"785b40",x"785b3f",x"79593d",x"78593f",x"806044",x"78583c",x"75563a",x"77583d",x"79593f",x"7a5b3f",x"77583e",x"74553c",x"73553b",x"76593f",x"78593e",x"7b5c40",x"78593f",x"795a3f",x"78593f",x"78593f",x"72553a",x"73563d",x"75573e",x"6f5439",x"674c36",x"6e513a",x"6d523c",x"755940",x"755942",x"725941",x"715640",x"634b36",x"674f3a",x"5c4532",x"614b37",x"5e4936",x"5e4b3b",x"605040",x"735e4c",x"735e4c",x"150e07",x"3b2a1b",x"3a2819",x"362617",x"342416",x"352517",x"312215",x"1a130c",x"5d422d",x"493423",x"412e1f",x"443120",x"43301e",x"412e1d",x"402d1d",x"402d1c",x"382617",x"3a2819",x"422e1d",x"44311f",x"3f2c1c",x"473322",x"412f1f",x"3d2b1b",x"422f1f",x"43301f",x"44311f",x"43311f",x"483423",x"402d1c",x"3c2a1a",x"3e2c1c",x"3d2b1b",x"3f2d1c",x"3f2d1c",x"3f2d1c",x"3c2a1a",x"3c2a1a",x"392819",x"3a2819",x"3b2919",x"3d2a1b",x"3e2b1b",x"392818",x"3a2919",x"382718",x"352517",x"302114",x"2b1d11",x"2d1f12",x"2b1d11",x"2f2114",x"261a0f",x"2f2115",x"271b10",x"22170d",x"21170d",x"21160d",x"21170d",x"150e07",x"433120",x"463220",x"432f1e",x"483322",x"402d1c",x"43301f",x"412e1d",x"3f2c1c",x"402d1c",x"402d1d",x"422e1d",x"412e1d",x"412e1d",x"473220",x"422e1d",x"44301e",x"45311f",x"412e1d",x"432f1e",x"3f2d1b",x"342315",x"3d2a1a",x"3d2b1a",x"453220",x"412e1e",x"433120",x"43301f",x"412e1d",x"453220",x"493422",x"473320",x"43311f",x"443221",x"3f2c1c",x"3d2b1b",x"3c2a1b",x"3b2a1a",x"3f2d1c",x"3a2819",x"362517",x"362517",x"332315",x"302114",x"2e2013",x"281c10",x"281c10",x"25190e",x"22170d",x"20160c",x"20170f",x"211911",x"1e160f",x"1d160f",x"1f1810",x"201811",x"1f1811",x"201912",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25170b",x"25170b",x"2b190c",x"2f1b0d",x"341d0e",x"351e0e",x"27160a",x"2e1a0b",x"2f1b0c",x"341d0e",x"321c0d",x"351d0d",x"351d0d",x"371e0d",x"331c0c",x"341c0c",x"381f0e",x"3a210f",x"39200e",x"3c220f",x"3a210f",x"3c220f",x"3a210f",x"39200e",x"3a200e",x"351d0d",x"351e0d",x"3c2210",x"3f2410",x"3b2310",x"37200f",x"38200f",x"351d0d",x"341c0c",x"331c0c",x"381f0e",x"38200e",x"39200f",x"381f0e",x"3a200f",x"38200e",x"341d0d",x"351d0d",x"381f0e",x"381f0e",x"3c220f",x"3a210f",x"3a210f",x"351e0e",x"38200e",x"361f0d",x"39200e",x"371f0e",x"371f0e",x"3c210f",x"351d0c",x"311b0b",x"2f1a0b",x"2f180b",x"321c0c",x"38200e",x"39200e",x"351d0d",x"38200e",x"3a220f",x"361f0e",x"301a0b",x"38200e",x"371f0e",x"351d0c",x"361e0d",x"371e0d",x"351e0d",x"381f0e",x"361f0f",x"371f0f",x"351f0f",x"2f1b0e",x"301b0c",x"2b180b",x"341d0d",x"351f0e",x"321c0c",x"3d2310",x"3b220f",x"24150a",x"2a190b",x"2b190b",x"1e1108",x"231409",x"271609",x"281609",x"2d190b",x"321c0c",x"341d0d",x"311b0c",x"311b0c",x"371f0d",x"381f0e",x"3d230f",x"3c230f",x"3b210f",x"3a210f",x"3a210f",x"3a210f",x"381f0e",x"39200e",x"412511",x"3b210f",x"3a200e",x"3c220f",x"3c2310",x"39200f",x"351d0d",x"311b0c",x"311c0c",x"341d0c",x"351d0c",x"3a200e",x"3f2410",x"3b210f",x"39200e",x"3a210f",x"3b220f",x"3d230f",x"3b210f",x"3b210f",x"311b0c",x"341d0d",x"361f0e",x"3a210f",x"3a210f",x"341e0e",x"3a210f",x"351d0d",x"311b0c",x"2c180b",x"351d0d",x"381f0e",x"3a210f",x"3a210f",x"381f0e",x"371f0e",x"371f0d",x"321c0c",x"361e0d",x"38200e",x"3d2310",x"38200f",x"39200e",x"3a210f",x"39200f",x"39200e",x"381f0e",x"381f0e",x"3a2210",x"3a210f",x"331c0c",x"3a210f",x"361e0d",x"3e2310",x"3d2310",x"3b2210",x"3c2310",x"341d0d",x"3a2110",x"181008",x"25150a",x"231409",x"402f23",x"332b24",x"180f07",x"1a1008",x"1c1108",x"36281f",x"453c33",x"3b2110",x"321d0d",x"2e1b0c",x"3e2310",x"4c311f",x"4c311f"),
(x"806750",x"806750",x"5e4e41",x"625142",x"5e4c3c",x"614d3b",x"644e3b",x"674f3b",x"6e543e",x"6e543e",x"6c533e",x"70543d",x"6a503b",x"68503b",x"6c5440",x"745944",x"785d45",x"795d44",x"765b42",x"775b43",x"7b5e44",x"795c43",x"765a41",x"775b42",x"75583f",x"775a3f",x"7c5d42",x"7b5c41",x"7c5d41",x"7c5e41",x"7e5f43",x"806045",x"7f5f43",x"806043",x"816145",x"826144",x"816042",x"7f5e41",x"7c5d41",x"805f43",x"7d5e41",x"7f5e40",x"7a5a3f",x"77583c",x"705238",x"715439",x"705338",x"75563b",x"75583d",x"7e5d41",x"7d5d42",x"7b5b3f",x"7c5d42",x"7d5d40",x"7d5d42",x"7d5d40",x"7a5a3f",x"78593f",x"7c5d42",x"7f5f43",x"7c5e42",x"7d5f45",x"7f6045",x"806045",x"7f6045",x"7d5e43",x"7e5f44",x"765840",x"785a41",x"76593f",x"7b5d42",x"775a42",x"785c43",x"735943",x"785b42",x"6b523b",x"604936",x"5c4632",x"604937",x"5c4737",x"5b493a",x"5c4b3c",x"735e4c",x"735e4c",x"150e07",x"3b2a1a",x"382718",x"382818",x"322315",x"322214",x"312215",x"21180e",x"5c432c",x"402f20",x"3f2f1f",x"443120",x"3e2c1c",x"412f1e",x"463221",x"412f1f",x"3f2c1c",x"3f2c1c",x"422f1f",x"3c2a1b",x"3d2c1c",x"3e2d1d",x"3d2b1c",x"3a2919",x"342416",x"382718",x"382718",x"3b2a1a",x"3d2b1b",x"3a291a",x"392819",x"3a2819",x"3a2819",x"3b2a1a",x"3c2a1b",x"382818",x"362617",x"352516",x"3a291a",x"39281a",x"382819",x"39281a",x"3b2a1b",x"3b2a1b",x"362718",x"362718",x"3a291a",x"352517",x"322316",x"291c10",x"2f2114",x"2c1f13",x"2a1d11",x"24190f",x"21170d",x"23180d",x"1f150b",x"1d130a",x"20150c",x"150e07",x"493422",x"3e2d1d",x"382819",x"3a2819",x"3f2c1c",x"382819",x"3a2919",x"3b291a",x"392819",x"3a2819",x"3d2b1c",x"432f1f",x"3d2b1b",x"3c2b1c",x"3a291a",x"412f1e",x"43301f",x"412f1e",x"412f1f",x"422f1f",x"3f2c1c",x"3a2919",x"412e1e",x"3d2c1c",x"3c2b1b",x"402e1d",x"3c2a1b",x"3a2919",x"3b2919",x"3b2919",x"3c2a1a",x"382718",x"3b2a1a",x"382818",x"392819",x"382818",x"372618",x"3a291a",x"362617",x"312215",x"322315",x"2f2013",x"2e2014",x"2b1e12",x"2b1e12",x"261b10",x"24190f",x"21170d",x"21170d",x"21180f",x"241a12",x"1f160f",x"201911",x"211912",x"1f1812",x"201912",x"1f1811",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"27180c",x"27180c",x"2d1a0d",x"311c0d",x"381f0f",x"351e0e",x"251509",x"28160a",x"28170a",x"2d190b",x"331d0d",x"361f0e",x"37200e",x"39210f",x"3e2411",x"3e2411",x"3b2210",x"39200e",x"341c0c",x"331c0c",x"361e0d",x"361d0d",x"341e0d",x"3d2612",x"3f2612",x"3d2411",x"3b2411",x"422813",x"412713",x"3f2713",x"3f2712",x"3a2411",x"3c2411",x"3c2210",x"3c2310",x"3b2210",x"3d2310",x"3e2410",x"381f0e",x"321c0c",x"321c0c",x"331c0c",x"361f0e",x"3b2210",x"412612",x"3b2210",x"3d2410",x"3c2310",x"3b220f",x"3a220f",x"3b210f",x"3a210f",x"3c2310",x"3a210f",x"3b210f",x"381f0d",x"361d0d",x"331d0c",x"321b0b",x"301a0b",x"341c0c",x"341d0c",x"361e0d",x"301a0b",x"341d0d",x"371f0e",x"371f0e",x"311b0c",x"341d0d",x"371f0e",x"38200e",x"38200e",x"351e0d",x"361f0e",x"3b220f",x"301c0e",x"341f0f",x"2f1b0e",x"2d1a0b",x"2d190b",x"341d0c",x"412511",x"341d0d",x"301c0c",x"301c0c",x"231509",x"29180b",x"2d1a0c",x"201309",x"26160a",x"2c180b",x"2c190b",x"2f1b0c",x"301b0c",x"2f1a0b",x"2e1a0b",x"311b0c",x"331c0c",x"381f0d",x"381f0d",x"331c0c",x"351c0c",x"341c0c",x"301a0b",x"321b0c",x"321b0b",x"341c0c",x"341c0c",x"331b0b",x"2f1a0b",x"301a0b",x"351d0d",x"361e0d",x"361f0e",x"351e0d",x"3a210f",x"402511",x"3e2411",x"412511",x"402410",x"391f0e",x"331c0c",x"371e0d",x"361d0c",x"351e0d",x"3b2310",x"3e2612",x"3d2411",x"3b2311",x"382210",x"412613",x"412713",x"402713",x"402713",x"3c2411",x"37200f",x"38200f",x"38210f",x"3c2310",x"38200f",x"3a200f",x"341d0d",x"321d0d",x"351c0c",x"361f0e",x"3c2210",x"3c2310",x"3e2411",x"3c2310",x"3b2210",x"39200f",x"3d2310",x"3a210f",x"3b220f",x"3e2310",x"361e0d",x"3a200f",x"351d0d",x"3a210f",x"361e0d",x"38200f",x"331c0d",x"371f0e",x"3a210f",x"341d0d",x"3d2310",x"191008",x"27160a",x"27170a",x"433023",x"322a23",x"180f08",x"1b1108",x"231409",x"402b1c",x"433b32",x"3e2110",x"321d0d",x"2c1a0c",x"3f230f",x"4b3120",x"4b3120"),
(x"7e644d",x"7e644d",x"5c4e42",x"5d4d3f",x"5d4c3c",x"5d4b3b",x"644f3d",x"674f3b",x"6a513c",x"6b523c",x"6d543e",x"634c38",x"705844",x"715945",x"705944",x"775c46",x"70563f",x"745a44",x"6f553f",x"755a43",x"735840",x"765a43",x"765941",x"7a5d43",x"7c5e41",x"7f5f44",x"7e5f45",x"785b41",x"7b5e43",x"7c5f44",x"7b5d42",x"7f5f43",x"7a5c41",x"7d5d40",x"7e5d41",x"785a3f",x"7a5a3e",x"73543a",x"77583d",x"79593e",x"79583d",x"7a5a3f",x"705339",x"6c5037",x"73563c",x"6f5138",x"725439",x"74553a",x"6f543a",x"795a3f",x"79583d",x"7b5b3f",x"75573a",x"75573c",x"73553c",x"7b5b3f",x"7b5d42",x"795b41",x"7c5c41",x"7e5e43",x"806043",x"826247",x"7a5b40",x"7c5d43",x"785b40",x"76593f",x"775a40",x"745740",x"6e533e",x"6b523b",x"71563f",x"755942",x"775b45",x"715843",x"6d5541",x"69523f",x"68523f",x"624c3b",x"5c4939",x"5b4838",x"57483b",x"5b4c3e",x"6d5948",x"6d5948",x"150e07",x"332315",x"332415",x"2b1d11",x"302114",x"302114",x"312215",x"251a0f",x"4d3723",x"372719",x"312215",x"2f2114",x"342517",x"312214",x"342416",x"302114",x"2f2014",x"2d1f13",x"2c1e12",x"2e1f13",x"2e1f13",x"322215",x"302114",x"2f2113",x"2f2114",x"2f2013",x"2e2013",x"2d1f12",x"2f2114",x"2c1e12",x"2a1d11",x"2a1d11",x"281b0f",x"2b1e11",x"2c1e12",x"2f2114",x"2c1e12",x"291d11",x"2a1d11",x"2b1d11",x"2b1d11",x"2e2013",x"2d1f13",x"2b1e12",x"302214",x"2a1d11",x"2a1d11",x"24190e",x"291c11",x"261a0f",x"24190e",x"20160c",x"20160c",x"20150c",x"1f150b",x"181008",x"191109",x"1c130a",x"181008",x"150e07",x"3f2d1c",x"312215",x"2e1f14",x"312214",x"2b1d11",x"2d2013",x"2a1d11",x"2f2114",x"2d1f13",x"312215",x"2e2013",x"2e2013",x"312315",x"302214",x"2f2014",x"2f2114",x"322416",x"322315",x"322316",x"302114",x"312215",x"2b1d11",x"302114",x"312214",x"302114",x"302114",x"2c1e12",x"2e2013",x"312215",x"2d1f12",x"2a1d11",x"2d1f12",x"2c1e12",x"2c1e12",x"291c10",x"2a1d11",x"291c11",x"2a1d11",x"2a1d11",x"2b1e11",x"281b10",x"2b1e11",x"251a0f",x"23180d",x"251a0f",x"21170d",x"1e140b",x"191109",x"1b130b",x"1c150d",x"1e160f",x"1c150e",x"1d1710",x"1d1610",x"1f1912",x"1f1811",x"1f1811",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b1a0d",x"2b1a0d",x"311c0d",x"341d0d",x"371e0f",x"392010",x"201309",x"2e1a0b",x"2c190b",x"301b0c",x"331d0d",x"331c0c",x"351d0d",x"2c190b",x"331c0c",x"341d0d",x"331c0c",x"2d180b",x"2d180a",x"211107",x"261207",x"371e0d",x"351c0c",x"341d0c",x"39200e",x"39200f",x"3a220f",x"3a210f",x"371f0e",x"38200e",x"3a210f",x"3a210f",x"3a210f",x"3b220f",x"3f2411",x"3e2411",x"3b2310",x"3a2310",x"402511",x"3a210f",x"39210f",x"351e0e",x"3b2210",x"39200f",x"38200e",x"3d2310",x"39200e",x"3b2210",x"3b2210",x"341d0d",x"3d2310",x"351f0e",x"3c2310",x"3b220f",x"3d220f",x"3a210f",x"3d2310",x"39210f",x"38200f",x"3b2210",x"3a2210",x"361f0e",x"371f0e",x"371f0e",x"321c0c",x"331d0d",x"311c0c",x"351d0d",x"371f0e",x"361f0e",x"331c0c",x"351d0d",x"371f0d",x"3b210f",x"331d0d",x"372010",x"351f0f",x"311d0e",x"321c0d",x"2a170a",x"331c0c",x"341e0e",x"341d0d",x"331d0d",x"331d0d",x"231409",x"2a190b",x"2d1a0c",x"1c1108",x"201309",x"2c190b",x"25160a",x"2e1a0b",x"2f1a0c",x"321c0c",x"321c0c",x"331d0d",x"361e0d",x"361e0d",x"351d0d",x"371e0d",x"361e0d",x"371e0d",x"371e0d",x"351d0c",x"341c0c",x"361e0d",x"361e0d",x"371e0d",x"381f0d",x"381f0e",x"371f0d",x"341d0d",x"301b0c",x"381f0e",x"381f0d",x"341d0d",x"301b0c",x"361e0d",x"321b0b",x"311a0b",x"271408",x"251107",x"341c0c",x"351d0c",x"331b0c",x"341d0d",x"3a210f",x"3b2210",x"38200f",x"38200e",x"3c2310",x"3a210f",x"3b2210",x"3d2310",x"3c220f",x"3e2310",x"3c2310",x"3e2311",x"3b2210",x"3d2411",x"39200f",x"38200f",x"38200e",x"3a210f",x"361f0e",x"351e0e",x"3a210f",x"3e2310",x"3b2210",x"412512",x"3c2310",x"3a210f",x"3a210f",x"402511",x"39200f",x"3b220f",x"351e0d",x"381f0e",x"3a210f",x"3a2210",x"3a2210",x"38210f",x"3e2511",x"351d0d",x"3d2411",x"1a1008",x"2b190b",x"2d1a0c",x"341d0c",x"372f26",x"180f08",x"1c1108",x"231409",x"503320",x"413830",x"3d2210",x"311c0c",x"301c0e",x"3b200e",x"4a301f",x"4a301f"),
(x"755d4a",x"755d4a",x"5a4e43",x"5c4f43",x"645243",x"695543",x"675240",x"68523e",x"6a5542",x"6f5642",x"725946",x"705844",x"745c48",x"79614d",x"80654f",x"785f4b",x"775e48",x"775d46",x"765c45",x"795d46",x"7d6047",x"765c45",x"7b5f45",x"795d43",x"795b42",x"7c6046",x"795c43",x"7a5d45",x"7b6049",x"7a5e46",x"7c5f45",x"7b5d44",x"795b40",x"72563e",x"816043",x"7f5f45",x"805e43",x"785a3f",x"72553a",x"75573d",x"76583c",x"7b5b41",x"77593d",x"7c5c40",x"78593e",x"7d5c41",x"7e5e41",x"77583e",x"77583d",x"795a3f",x"795b3f",x"785a3f",x"795c40",x"74573d",x"7a5c41",x"77593f",x"78593e",x"785a3f",x"7b5b41",x"7e6043",x"826348",x"7f6147",x"7c5e43",x"7e6148",x"7a5e45",x"785c44",x"7a5c44",x"7a5d46",x"755943",x"785b44",x"745a43",x"775c45",x"755a45",x"715844",x"6e5744",x"705a47",x"6e5846",x"715b48",x"6a5543",x"5e4d3d",x"56493c",x"574b40",x"645445",x"645445",x"150e07",x"26190e",x"281c10",x"261a0e",x"261a0f",x"23180d",x"25190e",x"20160c",x"3d2b1b",x"191109",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191109",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2c1b",x"181008",x"181008",x"191008",x"1c130a",x"181008",x"181008",x"181008",x"150e07",x"181008",x"191109",x"191109",x"191109",x"150e07",x"191109",x"1e140b",x"20160c",x"191109",x"1d140b",x"191109",x"1e140b",x"20160c",x"1c130a",x"1c130a",x"1f150b",x"1d130b",x"1f150b",x"1d140b",x"1c130a",x"191109",x"191109",x"1f150b",x"181008",x"181008",x"181008",x"191008",x"181008",x"181008",x"181008",x"181008",x"181008",x"181008",x"191109",x"191109",x"191109",x"191109",x"191109",x"150e07",x"17110a",x"19130c",x"1b150e",x"1c150e",x"1d1710",x"1e1711",x"1e1711",x"201912",x"1f1812",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1c0d",x"2f1c0d",x"331d0d",x"361e0e",x"3d2210",x"3c2211",x"231409",x"261409",x"2a1709",x"2d190b",x"351d0d",x"2e190b",x"3a200e",x"331c0c",x"341d0c",x"2f1a0b",x"2f1a0c",x"351d0d",x"351d0d",x"381f0e",x"361e0d",x"39200e",x"391f0e",x"38200e",x"3d2310",x"3b2210",x"3a210f",x"3d2310",x"3a220f",x"3c2310",x"36200e",x"3b210f",x"371f0e",x"371e0d",x"361e0e",x"371e0d",x"39200e",x"39200e",x"39200e",x"38200f",x"3c2310",x"38200e",x"3d2310",x"39200f",x"3d2310",x"3b220f",x"3c220f",x"3a200e",x"38200e",x"39210f",x"3a210f",x"321d0d",x"361f0e",x"3b2210",x"3c2310",x"39200e",x"3a210f",x"361e0d",x"331d0c",x"391f0e",x"341d0d",x"371f0e",x"341d0d",x"381f0e",x"341c0c",x"331c0c",x"351d0d",x"331c0c",x"331c0c",x"321c0c",x"371f0e",x"351e0e",x"371f0d",x"381f0e",x"3c220f",x"351e0f",x"3e2413",x"311d0e",x"311c0c",x"29170a",x"321b0c",x"3b210f",x"381f0e",x"38200f",x"361f0e",x"231509",x"28170b",x"2a180b",x"1d1108",x"201208",x"28160a",x"2a170a",x"27160a",x"2c190b",x"2c180a",x"2e190a",x"2d180a",x"2e190b",x"2f190b",x"2e180a",x"2c170a",x"2f190a",x"2d180a",x"251207",x"2c1609",x"2d180a",x"311b0b",x"2e180a",x"331b0b",x"2f190a",x"2f190a",x"361d0c",x"2f1a0b",x"2f1a0b",x"351d0d",x"301b0b",x"321c0c",x"351d0d",x"371f0e",x"371f0d",x"39200e",x"391f0e",x"361e0d",x"39200e",x"3a200e",x"381f0e",x"3a210f",x"39200f",x"3b2210",x"39200f",x"3e2410",x"3e2411",x"402511",x"3e2310",x"3a200e",x"371f0d",x"361e0d",x"381f0e",x"3d220f",x"361e0d",x"3c210f",x"38200f",x"3b2210",x"351e0e",x"38200e",x"39200f",x"311c0d",x"3b220f",x"3b220f",x"381f0e",x"3c220f",x"3a210f",x"3e2310",x"3e2310",x"412611",x"3f2411",x"3b2210",x"371f0e",x"39210f",x"39200f",x"3f2512",x"3d2411",x"38200f",x"3c2311",x"381f0e",x"3d2411",x"1a1008",x"2a180b",x"301b0d",x"493224",x"362d25",x"180f07",x"1c1108",x"211409",x"362111",x"3e352c",x"3f2311",x"311d0d",x"2b190c",x"3b200e",x"482f1e",x"482f1e"),
(x"7c6450",x"7c6450",x"876b54",x"896c54",x"83674f",x"83654d",x"85674e",x"85674e",x"836750",x"8f6e53",x"917155",x"8b6b50",x"8d6f54",x"917157",x"8d6e53",x"937356",x"937254",x"8d6d51",x"937255",x"89694c",x"8d6c50",x"8e6c50",x"8f6c4d",x"8e6c50",x"8b694d",x"8b6a4d",x"86664a",x"826148",x"836147",x"8c6a4d",x"8f6d4f",x"947254",x"8e6b4b",x"8e6b4d",x"8f6b4d",x"8f6b4d",x"896648",x"8a6649",x"896648",x"876446",x"876546",x"926d4e",x"916d4e",x"8d6849",x"8d6947",x"886548",x"856244",x"8a6749",x"8b6849",x"846144",x"896747",x"7f5f40",x"866347",x"876345",x"8a6648",x"866447",x"866549",x"866548",x"856447",x"816045",x"836147",x"8f6d51",x"8f6e51",x"937152",x"8f6d50",x"906e52",x"906f51",x"8f6d51",x"89684d",x"8a674c",x"86664c",x"896a4f",x"88694e",x"917155",x"937358",x"896b53",x"8f6f55",x"8b6d54",x"84674f",x"8f7054",x"8b6e54",x"856a54",x"745e4c",x"745e4c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"362618",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"19130c",x"1b140d",x"1b150e",x"1d1710",x"1d1610",x"1f1811",x"1f1811",x"211a13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0e",x"311c0e",x"351e0e",x"3b2110",x"3f2311",x"3b200e",x"27160a",x"2a170a",x"2d190a",x"321c0c",x"29170a",x"351d0d",x"361e0d",x"371f0e",x"2e1a0b",x"39200e",x"351e0e",x"341e0e",x"3b2210",x"39210f",x"3a210f",x"3a210f",x"3a210f",x"3c210f",x"3b220f",x"3a210f",x"3a210f",x"38200f",x"391f0e",x"3a210f",x"3a2110",x"39200e",x"371f0e",x"38200e",x"3b2210",x"3d2310",x"351e0d",x"3d2310",x"3a2210",x"3c2310",x"3b2210",x"3d2310",x"3c230f",x"3c220f",x"3a210f",x"3b220f",x"3c2310",x"3b220f",x"3c230f",x"3a200f",x"3a210f",x"38200e",x"341d0d",x"361e0e",x"321c0c",x"361f0d",x"39200e",x"361e0d",x"2e1a0b",x"301b0b",x"301b0b",x"331c0c",x"311c0c",x"361e0d",x"351e0d",x"351d0c",x"301a0b",x"2b180a",x"2a170a",x"311b0b",x"2f1a0b",x"331c0c",x"361e0d",x"351e0d",x"331c0c",x"361f10",x"351f10",x"341e0f",x"2a180b",x"28160a",x"331c0c",x"3d2311",x"3d2310",x"3b2210",x"38200e",x"24150a",x"27170a",x"2b180b",x"1d1208",x"221409",x"251509",x"27160a",x"2f1a0b",x"2d180a",x"2a160a",x"2e190b",x"371f0d",x"341d0d",x"351d0d",x"301b0c",x"341d0d",x"381f0e",x"38200e",x"371f0d",x"371f0d",x"371e0d",x"351d0d",x"351d0c",x"381f0d",x"391f0d",x"361d0d",x"361e0c",x"351d0d",x"341d0d",x"3a210f",x"3a210e",x"3b210f",x"3c230f",x"3a210f",x"3f2411",x"3f2410",x"3f2411",x"3b220f",x"3b210f",x"39200e",x"3a200f",x"371f0e",x"3b210f",x"3b2210",x"3b2210",x"371f0e",x"38200f",x"402511",x"3f2410",x"39200e",x"371f0e",x"38200e",x"3a2210",x"301b0c",x"3c2210",x"3e2410",x"3e2411",x"402511",x"3b220f",x"39200f",x"39200e",x"38200e",x"3a210f",x"3c2310",x"3b220f",x"3d2310",x"3d230f",x"3c220f",x"3b220f",x"38200e",x"3c2310",x"3a210f",x"371f0e",x"39200f",x"38200f",x"3c2311",x"351f0f",x"39210f",x"3d220f",x"341d0d",x"3f2411",x"191008",x"2a180b",x"311d0d",x"3c2515",x"352920",x"180f08",x"1c1108",x"211409",x"342011",x"362d25",x"432612",x"341f10",x"2c1a0c",x"3c210f",x"4a3020",x"4a3020"),
(x"705338",x"705338",x"6b4e35",x"735439",x"6f5137",x"674c34",x"71533a",x"73553a",x"705238",x"6e4f34",x"6e4f35",x"735438",x"77563a",x"765639",x"78583a",x"7d5c3e",x"7a593c",x"7b5a3c",x"7f5d3e",x"7d5b3d",x"7e5c3d",x"805c3e",x"7b593b",x"765638",x"765638",x"7d5a3d",x"7e5d40",x"866244",x"7f5d42",x"856345",x"846244",x"856345",x"856345",x"835f41",x"815e3f",x"7b593b",x"7d5b3e",x"7c5a3d",x"7e5d3f",x"79583b",x"836042",x"876344",x"815e41",x"815f41",x"7b5a3d",x"815f41",x"805e3f",x"7d5c3f",x"77573b",x"75553a",x"79583d",x"7a5a3e",x"7d5c3e",x"7c5b3e",x"856343",x"805e41",x"805e40",x"805f41",x"805d3f",x"7d5b3d",x"7a593a",x"795739",x"7f5c3d",x"805d3f",x"805c3d",x"7a5839",x"815d3f",x"7f5d40",x"7a593d",x"7d5d3e",x"75573b",x"79593d",x"7a593d",x"745539",x"705136",x"6b4d33",x"6c4e35",x"654931",x"5d432c",x"6d5037",x"6f5138",x"715338",x"705238",x"705238",x"201911",x"201911",x"1e160f",x"1e160f",x"1d160e",x"1e170f",x"1f1710",x"1f1710",x"1c150d",x"1e150c",x"1c130a",x"181008",x"1b1108",x"191008",x"181008",x"1f150c",x"22170d",x"23180d",x"22170d",x"23180d",x"24190e",x"291c11",x"251a0f",x"2a1d11",x"2a1d11",x"2a1d11",x"2a1d11",x"2c1e12",x"2b1e12",x"2b1e11",x"322215",x"2f2113",x"372617",x"322316",x"2d1f13",x"2f2114",x"362516",x"362517",x"342416",x"332315",x"322214",x"342415",x"332315",x"2e1f12",x"26180b",x"28190a",x"362617",x"372718",x"372618",x"362618",x"382718",x"3b291a",x"402d1e",x"413021",x"402f21",x"3f2f20",x"4c3826",x"19130c",x"191109",x"191109",x"1e140b",x"191108",x"1d140b",x"1c130a",x"23180d",x"20160c",x"23180d",x"1f150b",x"21170c",x"25190e",x"23170d",x"24190e",x"21160c",x"22170d",x"20160c",x"22170c",x"1c1208",x"201409",x"21160c",x"291c11",x"24190e",x"281c10",x"271b0f",x"281c10",x"291c11",x"2b1e12",x"2b1e12",x"2c1f12",x"302214",x"2c1f13",x"302215",x"302114",x"2b1e12",x"2d1f12",x"2d1f13",x"2c1e11",x"312214",x"2a1d11",x"2d1f13",x"2a1d11",x"2a1d11",x"2e1f13",x"2c1e12",x"322315",x"2f2013",x"2f2013",x"322214",x"2e1f12",x"2d1c0d",x"412910",x"150e07",x"2b1e11",x"2c1e12",x"2c1f12",x"2d1f12",x"2c1e12",x"26160a",x"150e07",x"19130c",x"19130c",x"171009",x"171009",x"17110a",x"17110a",x"171009",x"19130c",x"1a130c",x"1c150f",x"1b140e",x"1d160f",x"1d1710",x"1d1710",x"1c160f",x"1e1811",x"1e1811",x"1e1811",x"1d1710",x"1d1610",x"1d160f",x"1d160f",x"1c160f",x"1d1710",x"1c150f",x"1d160f",x"1d160f",x"1c150f",x"1c150e",x"1b150e",x"1b150e",x"1c150e",x"1b150e",x"1b150e",x"1b150e",x"1c150e",x"1b150e",x"1b150e",x"1c150e",x"1b150d",x"1b150e",x"1b150e",x"1b150e",x"1b140d",x"1b140e",x"1c150e",x"1c150e",x"1c150e",x"1b150e",x"1b140e",x"1c150e",x"1b140e",x"1d1710",x"1d1710",x"1e1710",x"1f1912",x"201912",x"201913",x"221b15",x"221b15",x"241d16",x"231c16",x"231c15",x"241d16",x"241d16",x"241d16",x"221b14",x"211a14",x"201a14",x"201913",x"1e1711",x"1e1710",x"1d1610",x"1d1610",x"1d1710",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341d0f",x"341d0f",x"331c0d",x"3a210f",x"402410",x"3b210e",x"29170a",x"2f1b0b",x"2f1b0b",x"331d0d",x"311b0c",x"381f0e",x"3a210f",x"3b220f",x"39200e",x"361e0d",x"3a200e",x"3d2310",x"422612",x"462813",x"432712",x"452813",x"432712",x"432712",x"412411",x"3f2411",x"3f2410",x"3f2310",x"3e2310",x"3e230f",x"3c220f",x"3c220f",x"3a210f",x"3d220f",x"3b210f",x"371e0d",x"391f0e",x"3a200e",x"381f0e",x"39200e",x"3c210f",x"3c220f",x"3e220f",x"3c210f",x"371e0d",x"351d0c",x"391f0d",x"371e0d",x"381f0d",x"371e0d",x"361e0d",x"3b200e",x"361e0d",x"331c0c",x"371e0d",x"3b210f",x"3a210e",x"371f0d",x"371e0d",x"351d0d",x"371e0d",x"381f0d",x"3a200e",x"3c210f",x"3b210f",x"3b200e",x"371f0e",x"341d0d",x"331d0d",x"3f2410",x"3a210f",x"381f0e",x"39200e",x"341c0c",x"371f0f",x"39200f",x"3a2110",x"321e0e",x"2a180b",x"2a180b",x"311b0c",x"3c2310",x"3a210f",x"412612",x"39210f",x"231509",x"29170b",x"2d1a0b",x"1f1209",x"2c1a0b",x"2b190b",x"2b180b",x"2e1a0b",x"341d0d",x"361e0d",x"381f0e",x"3b220f",x"3f2411",x"3e2410",x"3d2310",x"3d2310",x"3f2410",x"3e230f",x"3e2310",x"3d230f",x"3b210f",x"3c220f",x"3e220f",x"40240f",x"3b210e",x"3e220f",x"3a200e",x"341d0d",x"3e220f",x"3f2410",x"432712",x"402410",x"3b200e",x"3a1f0e",x"432611",x"462913",x"442813",x"432712",x"3f2511",x"432712",x"422612",x"3d230f",x"3e2410",x"3e2310",x"3e230f",x"3f2410",x"3e230f",x"3d230f",x"412511",x"3b210e",x"3b210f",x"3a200e",x"361e0d",x"331c0c",x"371f0e",x"351d0d",x"381f0e",x"3b210f",x"3c220f",x"3b210f",x"371e0d",x"351d0c",x"361d0c",x"351d0c",x"391f0d",x"361e0d",x"381f0d",x"371e0d",x"371f0d",x"361e0d",x"3b2210",x"371f0e",x"3a200e",x"341e0d",x"311c0c",x"361f0f",x"37200f",x"351e0e",x"3a2110",x"331d0d",x"381f0e",x"191008",x"28170a",x"311c0d",x"3e2514",x"342920",x"180f08",x"1c1108",x"211409",x"321c0e",x"372f27",x"3d2312",x"352010",x"2a190c",x"3a200e",x"4c3221",x"4c3221"),
(x"8e7056",x"907259",x"907156",x"886c53",x"7a5f4a",x"5a4b3d",x"5e4d3f",x"625142",x"645343",x"685646",x"695748",x"6b594a",x"675545",x"675647",x"635141",x"645242",x"625141",x"625142",x"655444",x"655444",x"665445",x"6d5a4a",x"6b5949",x"6b5948",x"6c5b4b",x"6e5b4b",x"6a5748",x"6c5949",x"6e5b4b",x"6e5c4b",x"6c5948",x"6b5847",x"6d5a49",x"6e5b4a",x"6b5a4a",x"6e5b4b",x"675646",x"6b594a",x"695747",x"695747",x"6c5949",x"675546",x"655444",x"695645",x"6b5847",x"695646",x"685646",x"695645",x"655343",x"665343",x"6a5747",x"695644",x"6c5949",x"6c5948",x"6b5848",x"6b5847",x"685546",x"695645",x"675241",x"695442",x"675341",x"685442",x"675241",x"634f3d",x"63513f",x"655241",x"645140",x"635141",x"614f3f",x"604e3f",x"5f4d3d",x"604e3f",x"624f3f",x"605041",x"625142",x"665342",x"635141",x"614f40",x"615040",x"82664d",x"886a50",x"8a6a50",x"8c6d51",x"8c6c51",x"201911",x"201811",x"201911",x"201911",x"201811",x"1f1710",x"211910",x"1e170f",x"1d150d",x"1b130b",x"191008",x"181008",x"181008",x"23180e",x"1d140b",x"20150c",x"20160c",x"21170d",x"25190e",x"25190e",x"23180d",x"23180d",x"261a0f",x"2a1d11",x"2b1e12",x"302215",x"2c1f12",x"2e2013",x"312214",x"2e2013",x"2e2013",x"312214",x"312114",x"302214",x"332315",x"332315",x"382818",x"342416",x"382819",x"382818",x"382718",x"362618",x"322315",x"302013",x"352516",x"3b2a1a",x"362517",x"332316",x"392818",x"352517",x"3e2b1b",x"402f1e",x"3f2d1e",x"402f20",x"413122",x"433223",x"553f2b",x"1b140e",x"1e160d",x"1d140b",x"191109",x"1d140b",x"1c130a",x"20160c",x"20160c",x"21170d",x"22170d",x"20150c",x"20160c",x"23180d",x"20160c",x"23180d",x"23180d",x"25190f",x"21170d",x"25190e",x"271b0f",x"261a0f",x"22170d",x"281b10",x"281b10",x"2a1d11",x"2e2013",x"281c10",x"2b1d11",x"2b1d11",x"2b1e12",x"2d2013",x"2b1e12",x"302214",x"2c1f12",x"312214",x"2e2013",x"2e2013",x"2d1f13",x"2c1e12",x"2a1d11",x"2d1f12",x"312215",x"322215",x"2e2013",x"2e1f13",x"332416",x"312215",x"312214",x"322315",x"322215",x"322214",x"412e1c",x"5d442c",x"150e07",x"2c1e12",x"302114",x"2f2013",x"312214",x"2e2013",x"211309",x"19120b",x"19120b",x"1c150d",x"1b130b",x"1b130b",x"1f160d",x"1b130b",x"1b130b",x"211810",x"1f170e",x"221911",x"1e170f",x"231a12",x"231a12",x"221a11",x"261c13",x"241c14",x"251b13",x"241b13",x"251b12",x"231a11",x"1f1811",x"231a12",x"241b13",x"251b13",x"241b13",x"231b13",x"261c13",x"221911",x"221911",x"221a11",x"231a11",x"241b11",x"251b12",x"231911",x"231911",x"221a11",x"241b11",x"241b12",x"241a11",x"221911",x"231a11",x"241a11",x"251b12",x"241a11",x"211910",x"221911",x"221911",x"241b11",x"241b12",x"221911",x"241b12",x"241b11",x"251c12",x"241a12",x"251c14",x"251c14",x"271e15",x"261e16",x"271f17",x"271e16",x"2a2118",x"2b2219",x"282017",x"2b2219",x"292018",x"292018",x"281f17",x"292017",x"261d15",x"261e16",x"261d15",x"211a12",x"221a12",x"231b13",x"241b12",x"241b12",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1a0c",x"2f1a0c",x"3e2411",x"3a200e",x"412511",x"3a200e",x"211308",x"2a170a",x"2c180a",x"2f1a0b",x"3c210e",x"3c2310",x"39200f",x"3c2310",x"371f0e",x"3a210f",x"39210e",x"39210f",x"351e0d",x"361f0e",x"341d0d",x"38200e",x"381f0e",x"39200e",x"381f0f",x"331c0c",x"281408",x"331d0d",x"38200e",x"3a210f",x"3b210f",x"361e0d",x"39210f",x"3a220f",x"3b210f",x"3c2210",x"3e2411",x"402511",x"3f2411",x"3f2411",x"402511",x"3e230f",x"3b2210",x"3d2310",x"3a200e",x"3e2410",x"412612",x"3c2310",x"3a210f",x"371e0e",x"3b210f",x"3b220e",x"39200f",x"392210",x"381f0e",x"361e0d",x"3a210f",x"3b210f",x"3c220f",x"3d230f",x"3d220f",x"3d2310",x"361d0d",x"361d0d",x"381e0d",x"341c0c",x"3a200e",x"3a200e",x"39200d",x"3a200e",x"3c210f",x"381f0e",x"3b220f",x"361f0e",x"392010",x"3e2511",x"3c2311",x"311d0e",x"311c0d",x"2d1a0c",x"321b0c",x"3a2110",x"39210f",x"3e2411",x"38200e",x"221409",x"2a190b",x"2d1a0b",x"201309",x"2b190b",x"311c0d",x"351e0d",x"3c220f",x"3e2411",x"321d0d",x"2c190b",x"301b0c",x"361f0e",x"37200f",x"341f0e",x"36200f",x"3a2210",x"3a2110",x"351e0e",x"38200f",x"361f0e",x"3a210f",x"38200f",x"38200e",x"381f0e",x"361f0e",x"3b2210",x"3b220f",x"3a210f",x"38200e",x"3c2311",x"3d2310",x"3e2310",x"3d2210",x"3f2411",x"3c220f",x"3d2310",x"402511",x"3e2310",x"3b2210",x"39200e",x"3c210f",x"3b210f",x"3e2310",x"3b210f",x"371f0e",x"38200e",x"39200e",x"3d210e",x"3d220e",x"40230f",x"391f0d",x"391f0d",x"3b200e",x"3b200e",x"3d210f",x"391f0e",x"381f0d",x"3b200d",x"3b200d",x"3d220e",x"3f230f",x"432510",x"432611",x"371f0d",x"3c220f",x"361e0d",x"371f0d",x"361e0d",x"361e0c",x"38200f",x"3d2311",x"371f0e",x"341d0d",x"39200f",x"3b2210",x"351f0e",x"301c0c",x"3a2210",x"321c0c",x"351d0d",x"191008",x"26160a",x"301c0d",x"412816",x"33271e",x"180f08",x"1b1108",x"211409",x"341e10",x"372f27",x"412513",x"2e1c0e",x"2b190c",x"381e0d",x"473021",x"473021"),
(x"8e7056",x"907259",x"907156",x"886c53",x"7a5f4a",x"5a4b3d",x"5e4d3f",x"625142",x"645343",x"685646",x"695748",x"6b594a",x"675545",x"675647",x"635141",x"645242",x"625141",x"625142",x"655444",x"655444",x"665445",x"6d5a4a",x"6b5949",x"6b5948",x"6c5b4b",x"6e5b4b",x"6a5748",x"6c5949",x"6e5b4b",x"6e5c4b",x"6c5948",x"6b5847",x"6d5a49",x"6e5b4a",x"6b5a4a",x"6e5b4b",x"675646",x"6b594a",x"695747",x"695747",x"6c5949",x"675546",x"655444",x"695645",x"6b5847",x"695646",x"685646",x"695645",x"655343",x"665343",x"6a5747",x"695644",x"6c5949",x"6c5948",x"6b5848",x"6b5847",x"685546",x"695645",x"675241",x"695442",x"675341",x"685442",x"675241",x"634f3d",x"63513f",x"655241",x"645140",x"635141",x"614f3f",x"604e3f",x"5f4d3d",x"604e3f",x"624f3f",x"605041",x"625142",x"665342",x"635141",x"614f40",x"615040",x"82664d",x"886a50",x"8a6a50",x"8c6d51",x"8c6c51",x"201811",x"201911",x"201912",x"1f170f",x"201911",x"201911",x"1e170f",x"1f1710",x"1d150d",x"20160d",x"191109",x"191109",x"20160c",x"1e140b",x"20160c",x"21170c",x"23180d",x"23180d",x"261a0f",x"261a0f",x"2a1d11",x"281b10",x"281b10",x"2a1d11",x"291c10",x"2b1e11",x"2d1f13",x"322315",x"2d1f12",x"322315",x"362617",x"342416",x"342416",x"362617",x"372718",x"322315",x"332315",x"382718",x"3a2919",x"382718",x"372718",x"3b2a1a",x"382718",x"342416",x"372718",x"392818",x"342416",x"362617",x"3f2d1c",x"3a2919",x"3e2c1c",x"3d2c1d",x"3c2c1e",x"3f2e20",x"402f21",x"3d2d20",x"513b28",x"1b150e",x"1f160d",x"1e140b",x"191109",x"1e140b",x"191109",x"1d140b",x"21160c",x"21160d",x"23180d",x"21170d",x"22170d",x"23180e",x"251a0f",x"261a0f",x"20160c",x"24180e",x"23180d",x"25190e",x"291c10",x"251a0f",x"25190f",x"281c10",x"291c10",x"2c1f12",x"2d2013",x"2f2114",x"2a1d11",x"281b10",x"2d1f12",x"2e1f13",x"2b1d11",x"2f2114",x"2e1f13",x"342416",x"2f2013",x"2d2013",x"2d2013",x"322316",x"312315",x"362617",x"312215",x"2c1e12",x"2b1e12",x"2d2013",x"312215",x"352517",x"322416",x"362617",x"312214",x"332415",x"3f2c1c",x"5c422b",x"150e07",x"2e2013",x"312315",x"322315",x"342416",x"362617",x"170f07",x"19130c",x"19130c",x"1b130c",x"1b120a",x"1f150c",x"1b130c",x"20160d",x"1f160d",x"21180f",x"21170f",x"1e160f",x"1f1710",x"251b13",x"231b13",x"231a12",x"231b12",x"241b13",x"231b12",x"231a11",x"241b13",x"241a12",x"221a11",x"231a12",x"261c13",x"241b12",x"261d14",x"231910",x"241a11",x"221911",x"251a11",x"251a11",x"241b11",x"241a11",x"221911",x"241b11",x"221a11",x"221911",x"241b12",x"261c12",x"241b11",x"251a11",x"251a12",x"241b12",x"241b12",x"251b12",x"241b11",x"241a11",x"221911",x"261b13",x"251b12",x"231911",x"241b11",x"251b12",x"231b12",x"261d14",x"261d14",x"261c14",x"271d14",x"281e16",x"271d15",x"2a2018",x"2b2118",x"291f17",x"2b2219",x"282018",x"282017",x"271f17",x"281f17",x"261d15",x"261d15",x"251b13",x"241c13",x"241a11",x"241b12",x"241b13",x"231a11",x"231a11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"361f0f",x"361f0f",x"371e0f",x"381e0e",x"422611",x"371f0d",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"17110a",x"19120c",x"19130c",x"1c150e",x"1c150f",x"1a130c",x"321c0d",x"371f0e",x"4d2e15",x"3b2211",x"331d0e",x"27160a",x"341d0c",x"3d2310",x"3a210f",x"3a220f",x"361f0e",x"211309",x"29180b",x"301c0d",x"231409",x"19120b",x"160f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f08",x"180f08",x"180f07",x"180f07",x"170f07",x"180f07",x"180f07",x"180f08",x"180f07",x"180f07",x"180f08",x"180f08",x"180f08",x"181008",x"191109",x"1b130b",x"1c150e",x"1c150e",x"1c150e",x"492912",x"371e0e",x"402511",x"3a200e",x"3e2411",x"3b2210",x"3b2310",x"402612",x"36200f",x"36200f",x"311b0c",x"361f0e",x"180f07",x"261509",x"2e1b0d",x"3f2613",x"2e231a",x"191008",x"1b1108",x"23150b",x"321d0f",x"3d342c",x"4c433a",x"503929",x"2c1a0c",x"3b200e",x"493223",x"493223"),
(x"816853",x"8e7159",x"7f6752",x"7a614c",x"6e5743",x"52463b",x"4d4035",x"584b3f",x"584b3f",x"584a3d",x"594b3f",x"574b3e",x"514539",x"56473b",x"55473a",x"55483c",x"524539",x"534538",x"54473b",x"58493c",x"584a3e",x"5b4c3d",x"5d4f41",x"5c4e41",x"5d4d3e",x"5e5042",x"5a4b3f",x"5c4e40",x"5e4f42",x"615244",x"5d4e41",x"5a4a3b",x"5f5042",x"5b4d40",x"605145",x"605245",x"5e5042",x"5f5143",x"5f5143",x"5e4e40",x"5a4d41",x"554638",x"5a4a3b",x"564738",x"574738",x"5a4a3c",x"534336",x"5a4a3d",x"58493a",x"5b4c3e",x"5a4a3c",x"594a3c",x"5c4c3d",x"5b4b3c",x"5e4e3f",x"5a4b3d",x"5b4b3e",x"56483b",x"58493b",x"554638",x"55473b",x"544538",x"56473a",x"52463a",x"524538",x"544639",x"55473a",x"56493c",x"524439",x"544538",x"524537",x"514338",x"55483d",x"53473b",x"55473c",x"55473b",x"54463a",x"54473b",x"4f4235",x"795f48",x"83664b",x"8c6d53",x"6f5945",x"755d48",x"241b13",x"221a13",x"221a13",x"221a13",x"201911",x"201811",x"1e170f",x"1e170f",x"1d150d",x"1b130b",x"1d140b",x"23180d",x"20150c",x"24190e",x"21170c",x"21170c",x"20150b",x"20150b",x"271a0f",x"23180d",x"24180e",x"23180d",x"291c11",x"2b1e12",x"2e2013",x"2c1e12",x"2c1f12",x"312316",x"332416",x"342517",x"362618",x"342516",x"392819",x"3a291b",x"38281a",x"3b2a1c",x"3c2b1c",x"3a291a",x"3a291a",x"342416",x"342416",x"39281a",x"362618",x"382718",x"352416",x"352517",x"342415",x"352516",x"352516",x"392818",x"372719",x"3d2c1d",x"3d2d1f",x"413022",x"433223",x"423122",x"57402c",x"1c150f",x"20170d",x"22170d",x"1e150b",x"1f150c",x"1f150c",x"1e150b",x"1e150b",x"22170d",x"1f150c",x"1f150c",x"22170d",x"21170d",x"261a0f",x"25190f",x"23180d",x"261a0f",x"23180d",x"25190e",x"271b0f",x"24190e",x"261a0f",x"281c10",x"2d1f12",x"271b0f",x"281c10",x"2a1d11",x"271a0f",x"312114",x"312315",x"2c1e12",x"2c1e12",x"302214",x"2e2014",x"2f2115",x"2e2014",x"362619",x"312215",x"352517",x"352517",x"2f2115",x"372719",x"352618",x"342517",x"302214",x"362618",x"332316",x"322315",x"362617",x"382718",x"322315",x"402d1c",x"583f29",x"150e07",x"2e2013",x"332315",x"312214",x"312214",x"322315",x"150e07",x"19130c",x"19120c",x"1b130b",x"1b130b",x"191109",x"1e150b",x"23190f",x"1b130b",x"221810",x"211810",x"231a11",x"231a11",x"241b12",x"251c13",x"251b13",x"251c13",x"261d14",x"241a12",x"231a12",x"241b13",x"241b13",x"231b12",x"241b13",x"241a12",x"221a11",x"20180f",x"231a11",x"241911",x"221910",x"221911",x"221911",x"211810",x"251b12",x"231a11",x"251c12",x"261c13",x"261c13",x"251c12",x"251c12",x"251b12",x"231a11",x"231a12",x"251c12",x"261c13",x"261c12",x"261d13",x"261c12",x"251b12",x"231a11",x"261b13",x"251c12",x"241b12",x"251a12",x"251b12",x"261c13",x"251c13",x"271d14",x"261d14",x"271e15",x"281e16",x"291f17",x"281f16",x"271f17",x"271e16",x"292017",x"281f16",x"271e15",x"271e16",x"291f16",x"261d14",x"2a2017",x"201911",x"251b13",x"231a11",x"231a11",x"211910",x"211910",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"382011",x"382011",x"351d0d",x"301a0d",x"3f2310",x"3b220f",x"341d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"19120b",x"1b140e",x"1b140d",x"1c150e",x"1b140d",x"1b140d",x"573821",x"492c15",x"382110",x"311b0b",x"29180b",x"321c0c",x"3a210f",x"3b220f",x"3b210f",x"3a210f",x"231509",x"27170a",x"301c0d",x"1c150e",x"19120b",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"170f07",x"191109",x"1a130b",x"1c150d",x"1c150e",x"1c140d",x"4a2913",x"3a210f",x"3a210f",x"381f0e",x"39200e",x"402612",x"38200f",x"3e2511",x"3c2310",x"402612",x"351d0d",x"3e2411",x"180f07",x"26160a",x"2d1a0c",x"3d2412",x"2f251d",x"180f07",x"1c1108",x"23160b",x"2e1c0e",x"3e352d",x"51483e",x"513522",x"351f0e",x"492912",x"483020",x"483020"),
(x"735f4e",x"735f4d",x"5b4f43",x"53463b",x"4d4136",x"504439",x"4f4236",x"514539",x"52463b",x"52463a",x"4f4439",x"4a3e34",x"463b30",x"4d4033",x"4f4134",x"514337",x"4d3f32",x"504236",x"4f4135",x"514235",x"56483b",x"524437",x"524337",x"554537",x"524438",x"544539",x"524337",x"514235",x"504134",x"56483a",x"564739",x"554538",x"544537",x"57493c",x"584a3c",x"58483a",x"594a3d",x"5c4d40",x"594a3d",x"58493c",x"57483b",x"504235",x"4c3e32",x"473a2f",x"4d3f33",x"524133",x"524234",x"554434",x"524132",x"514133",x"4f3f32",x"534335",x"514133",x"544436",x"554538",x"524336",x"544538",x"544538",x"4f4135",x"504235",x"53463a",x"54473a",x"504236",x"534538",x"534539",x"4e3f31",x"504236",x"504336",x"4f4134",x"4c3f33",x"4e4034",x"4d3f34",x"4b3e32",x"4b3d32",x"463a30",x"44382f",x"483c31",x"493b30",x"504236",x"4c3f34",x"4b3d31",x"514336",x"4d4137",x"5d4c3d",x"211912",x"211912",x"231b14",x"211912",x"221a13",x"201811",x"201811",x"1e160f",x"1a120a",x"181008",x"191109",x"20150c",x"1f150c",x"22170d",x"1d130b",x"23180d",x"21160c",x"22170d",x"281c10",x"26190e",x"271a0f",x"261a0f",x"21150a",x"1f1409",x"291c10",x"2d1f12",x"2f2114",x"2f2114",x"312214",x"302114",x"2d1f12",x"382719",x"392919",x"362618",x"372719",x"392819",x"342517",x"382819",x"372617",x"352416",x"2e1f13",x"352517",x"392819",x"382718",x"352517",x"372718",x"3a291a",x"362616",x"372618",x"392819",x"3c2b1c",x"3a2a1c",x"3d2d20",x"3c2d1f",x"36261a",x"302318",x"4c3725",x"1d160f",x"20160d",x"1e140b",x"1d140b",x"1d140b",x"1d140b",x"21160d",x"21170d",x"21170d",x"23180e",x"20160c",x"23180e",x"20150c",x"23180e",x"23170d",x"20150c",x"23180e",x"24190e",x"281b10",x"271b10",x"22170d",x"2b1d11",x"261a0e",x"2b1e12",x"291c11",x"2a1d11",x"281b0f",x"302114",x"281b0f",x"22150a",x"1f1409",x"2b1d11",x"322215",x"342416",x"2d2013",x"2c1e12",x"2d1f13",x"302114",x"2d2013",x"392819",x"352517",x"2d2013",x"332416",x"312315",x"332316",x"2f2114",x"342315",x"2d1f12",x"342416",x"362618",x"332316",x"412e1e",x"59402a",x"150e07",x"2d1f13",x"312214",x"322315",x"312214",x"332214",x"150e07",x"19130c",x"19130c",x"19110a",x"1c130a",x"191109",x"191109",x"1b130b",x"1b130c",x"1f160d",x"20170f",x"1d150e",x"231a11",x"221a10",x"201911",x"241b13",x"231a12",x"231a12",x"251c13",x"231b13",x"221912",x"251c13",x"211910",x"221911",x"221911",x"241911",x"221910",x"211910",x"211810",x"211911",x"231a11",x"231910",x"22180f",x"21180f",x"1e150d",x"1d150c",x"241910",x"231910",x"241911",x"241911",x"231910",x"20180f",x"20170f",x"241910",x"241a11",x"241a11",x"23190f",x"231910",x"23190f",x"20180f",x"1f160e",x"221810",x"231911",x"231910",x"251a12",x"241a11",x"251b12",x"261c14",x"281f16",x"251c12",x"261e16",x"281e16",x"292018",x"291f17",x"271f17",x"251d15",x"251d15",x"231b14",x"251d14",x"251c15",x"261c14",x"251b13",x"231b13",x"221a11",x"221911",x"221810",x"1f160f",x"1f160f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"382111",x"382111",x"351d0e",x"251309",x"3e2310",x"351d0d",x"2e1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"1c1108",x"1f1208",x"231409",x"1f1309",x"231409",x"221409",x"1f1309",x"1f1208",x"1f1208",x"1c1108",x"1d1108",x"1c1108",x"1c1008",x"1b1008",x"191008",x"1a1008",x"1d1108",x"191008",x"1c1108",x"1d1208",x"150e07",x"1d1108",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"211309",x"1f1208",x"1d1108",x"150e07",x"201309",x"1e1208",x"1a1008",x"150e07",x"1a1008",x"1e1208",x"1c1108",x"1b1108",x"1b1008",x"1d1108",x"1c1108",x"1d1108",x"1e1108",x"1d1108",x"150e07",x"150e07",x"1c1108",x"23150b",x"19120b",x"21170e",x"1f160f",x"1c150e",x"1c150e",x"1c150e",x"533723",x"452913",x"351f0f",x"2e1a0b",x"27170a",x"351d0d",x"3a210f",x"3a210f",x"39200e",x"3b220f",x"23150a",x"27170a",x"2d1a0c",x"1d160f",x"1c150e",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"1a1008",x"180f08",x"150e07",x"150e07",x"1a1008",x"150e07",x"150e07",x"1a1008",x"180f08",x"150e07",x"1b1108",x"160e07",x"160e07",x"180f07",x"180f07",x"160f07",x"160e07",x"170f07",x"160e07",x"1a1007",x"180f07",x"191008",x"190f07",x"170f07",x"170f07",x"190f07",x"190f07",x"1c1108",x"170f07",x"1a1008",x"1c1108",x"191008",x"170f07",x"170f07",x"18110a",x"1e150d",x"1c150e",x"1e1610",x"1e1610",x"4d2c15",x"3a210f",x"39200f",x"321c0c",x"38200e",x"402612",x"422712",x"412612",x"39200f",x"402612",x"2f1a0b",x"39210f",x"180f08",x"26160a",x"2d1b0d",x"3e2412",x"30261e",x"191008",x"1c1108",x"23150b",x"2f1b0e",x"3e342c",x"51483e",x"221409",x"2f1b0d",x"4e2d15",x"482912",x"482912"),
(x"866b54",x"856951",x"574a3e",x"534639",x"52453a",x"514438",x"4d4034",x"514539",x"514438",x"4e4136",x"4a3e33",x"483b30",x"493e34",x"473b2f",x"483c31",x"4e4136",x"4e4034",x"4b3e32",x"4f4135",x"4e3f33",x"4c3d31",x"4e4034",x"4f4133",x"4f4134",x"4e3f32",x"4f4032",x"4e3d2f",x"4f3f31",x"4f3e30",x"544434",x"554334",x"534234",x"514133",x"544435",x"544336",x"534336",x"564538",x"534234",x"544537",x"504133",x"554535",x"504133",x"504133",x"4d3d30",x"47392c",x"4b3b2d",x"47382b",x"4d3c2e",x"4b3c2e",x"4e3e30",x"4e3e31",x"4e3e30",x"524133",x"4e3f31",x"503f31",x"4d3e31",x"4f3f32",x"4e3f31",x"4b3d31",x"4b3b2e",x"504133",x"4e3e30",x"4f3f32",x"544436",x"514235",x"4c3e31",x"4b3d30",x"4c3e31",x"4b3c30",x"4c3e32",x"4e3f31",x"483a2f",x"4b3d31",x"483b2e",x"43362a",x"44372c",x"46392e",x"473b2f",x"473b30",x"473a2f",x"483b30",x"4c3f32",x"58493b",x"56473a",x"261d16",x"271e16",x"231b14",x"221b14",x"261d15",x"221a13",x"201710",x"231911",x"20180f",x"1e150b",x"1e140b",x"1d140b",x"251a0f",x"20160c",x"24190e",x"23180d",x"22170d",x"22170d",x"24190e",x"24180e",x"2d2013",x"281c0f",x"271a0f",x"25190e",x"25190e",x"271a0f",x"281b0f",x"2a1c11",x"2b1d11",x"2e2013",x"302215",x"312215",x"322315",x"342416",x"372718",x"352517",x"382718",x"3b291a",x"372617",x"3f2d1c",x"3b291a",x"3d2b1c",x"3e2b1c",x"3d2b1c",x"342517",x"3a291a",x"392819",x"3e2b1b",x"3c2a1a",x"392a1b",x"3f2d1e",x"3b2b1e",x"443324",x"3d2e20",x"413122",x"403022",x"4b3624",x"1d160f",x"1d140c",x"1c130a",x"181008",x"1c130a",x"1d130b",x"1d130a",x"1d140b",x"24180e",x"22170d",x"20150c",x"20160c",x"25190f",x"22170d",x"291c11",x"23180d",x"2c1f13",x"291c11",x"291c11",x"251a0f",x"2b1e12",x"291d11",x"25190e",x"24190e",x"2d1f13",x"2c1e12",x"2b1d11",x"2f2114",x"291c10",x"2b1e11",x"2a1c11",x"25190e",x"281b0f",x"2c1e12",x"2e1f12",x"2b1e11",x"2f2114",x"2c1f12",x"302114",x"302114",x"2c1f12",x"2d1f13",x"302114",x"2d1f13",x"322316",x"352517",x"372718",x"382718",x"362718",x"372718",x"342517",x"43301f",x"5c422c",x"150e07",x"322315",x"332416",x"332416",x"362618",x"372618",x"150e07",x"17110a",x"17110a",x"181008",x"181008",x"181008",x"181008",x"181008",x"1e150c",x"1e150c",x"20160f",x"20160e",x"251b12",x"231a11",x"221911",x"1e170f",x"231b12",x"221911",x"211910",x"251b12",x"221911",x"221910",x"231911",x"221911",x"241b11",x"231910",x"23180f",x"231910",x"231910",x"231910",x"231910",x"221910",x"241a11",x"22190f",x"231910",x"21170f",x"20170e",x"1e160d",x"21170f",x"21170f",x"22190f",x"1f160d",x"221910",x"22180f",x"23190f",x"221810",x"23180f",x"231a10",x"21180f",x"231910",x"231810",x"231910",x"231910",x"241a10",x"251b12",x"241b11",x"241b12",x"251c13",x"251b12",x"271e15",x"241c14",x"241c14",x"261d15",x"271d16",x"271d15",x"261d16",x"271e16",x"231a12",x"231a12",x"221911",x"221911",x"211810",x"211910",x"1f170e",x"1c140d",x"20160e",x"20170e",x"20170e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351f10",x"351f10",x"371f10",x"251308",x"3f2412",x"361d0d",x"2b190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"150e07",x"180f07",x"221409",x"24150a",x"26160a",x"28180b",x"28180b",x"2a180b",x"29180b",x"2c1a0c",x"2a190b",x"2b190b",x"2a190b",x"27170b",x"27160a",x"241509",x"261509",x"29170a",x"241509",x"211309",x"231409",x"241509",x"24150a",x"1f1309",x"211309",x"231409",x"1d1108",x"1e1208",x"1f1208",x"25150a",x"25160a",x"241509",x"26160a",x"2b180b",x"241509",x"2c190b",x"26160a",x"2a180b",x"29170b",x"28170a",x"1b1108",x"27160a",x"26160a",x"27160a",x"211309",x"221409",x"27160a",x"221409",x"211409",x"231509",x"25160a",x"221409",x"1c1108",x"1f1309",x"231409",x"26170b",x"1b130c",x"21170e",x"1f160e",x"19130c",x"19130c",x"573e2c",x"40230e",x"361f0d",x"2e1a0c",x"2d1a0b",x"361e0d",x"381f0e",x"38200e",x"371e0d",x"38200f",x"221409",x"28180b",x"321d0e",x"1f1912",x"1c150e",x"171009",x"150e07",x"150e07",x"191008",x"221409",x"1c1108",x"241509",x"1a1008",x"150e07",x"1f1208",x"211309",x"1f1208",x"1f1208",x"1e1208",x"221409",x"231409",x"1d1108",x"1f1309",x"1b1108",x"1f1208",x"211309",x"1f1208",x"201309",x"26160a",x"25160a",x"29180b",x"24150a",x"27170a",x"231509",x"1e1208",x"1d1208",x"29180b",x"2a190b",x"25160a",x"29180b",x"29180b",x"29180b",x"22140a",x"28180b",x"22150a",x"221409",x"231409",x"1e1208",x"241509",x"221409",x"1f1208",x"221409",x"241509",x"211409",x"24150a",x"231409",x"211409",x"201309",x"231409",x"241509",x"241509",x"26160a",x"25150a",x"201309",x"26170d",x"291a0f",x"291b11",x"241911",x"1d160f",x"482913",x"3f2410",x"3d2410",x"361e0d",x"3a210f",x"442813",x"412612",x"432813",x"351d0d",x"3b2311",x"311a0b",x"3d2310",x"180f07",x"26160a",x"2b190b",x"3f2514",x"2c2119",x"191008",x"1c1108",x"23150b",x"2f1a0d",x"342b23",x"52483e",x"52483e",x"2f1b0d",x"4e2d15",x"482912",x"000000"),
(x"8b6f56",x"886b52",x"5a4d40",x"574b3e",x"51453a",x"504337",x"4b3e32",x"4d3f32",x"4a3d31",x"4a3d31",x"4c3e32",x"4b3d30",x"45372b",x"483a2d",x"514336",x"504235",x"504235",x"524336",x"504236",x"504032",x"534335",x"574739",x"514235",x"504134",x"4c3d2f",x"49392c",x"48382b",x"423327",x"48382b",x"4d3d2f",x"4c3c2d",x"514031",x"504032",x"503f31",x"4f3e30",x"4e3d2d",x"503f31",x"4e3e30",x"504031",x"4d3d2d",x"4c3c2d",x"493b2d",x"514031",x"503f30",x"544030",x"4d3d2e",x"544232",x"4d3d2f",x"544333",x"544233",x"4f3e30",x"514031",x"574535",x"514132",x"4e3e30",x"4b3b2d",x"483a2e",x"443629",x"44362a",x"403327",x"493a2e",x"4a3b2e",x"4a3a2d",x"4c3d30",x"4c3d2f",x"4c3d2f",x"4a3b2e",x"4d3e2f",x"4b3b2e",x"4f3f31",x"483a2d",x"4c3c2f",x"483a2e",x"46382d",x"4b3c2f",x"493c30",x"4d3f33",x"483b2e",x"4d3f33",x"4c3e31",x"4e4134",x"534538",x"604f41",x"5b4b3c",x"261d15",x"231c15",x"231c14",x"241c15",x"221b14",x"201911",x"1f1811",x"1d150e",x"1f160e",x"191009",x"1d130a",x"23180d",x"1e140b",x"23180e",x"24190e",x"20160d",x"23180e",x"24190f",x"2a1d12",x"2a1d12",x"281b0f",x"261a0f",x"2c1e12",x"2e2013",x"322316",x"312215",x"302214",x"322416",x"352618",x"352618",x"2f2114",x"352617",x"372719",x"3d2c1d",x"3c2b1c",x"382819",x"382718",x"332315",x"342416",x"2b1b0e",x"312214",x"382719",x"382718",x"3c2a1b",x"402d1d",x"3a291a",x"3a291a",x"3e2c1c",x"3f2d1d",x"433122",x"433123",x"453425",x"413222",x"3f3022",x"413123",x"463526",x"614832",x"1f1811",x"21190f",x"20170d",x"1e150c",x"21170d",x"1e140b",x"21160d",x"21170d",x"22170d",x"22170d",x"261a0f",x"24190e",x"261a0f",x"20160c",x"1d1309",x"20150c",x"291c11",x"271a0f",x"25190e",x"23180e",x"291c11",x"24180e",x"291d11",x"291c11",x"302215",x"2c1f13",x"2c1f13",x"2a1d11",x"2c1e11",x"312215",x"2d2013",x"2f2114",x"2d1f13",x"322416",x"2f2214",x"332517",x"352618",x"342416",x"362617",x"372719",x"342518",x"2f2115",x"342517",x"322316",x"332315",x"302013",x"27190c",x"332315",x"322315",x"312215",x"322316",x"493422",x"5a412b",x"150e07",x"342416",x"352517",x"362719",x"39281a",x"3a2a1b",x"150e07",x"17110a",x"150e07",x"191109",x"191109",x"191109",x"191109",x"1e150b",x"191109",x"1b130b",x"20160d",x"21170f",x"211910",x"231a11",x"261b12",x"261b13",x"221a11",x"20180f",x"211910",x"20170f",x"20160f",x"20180f",x"22180f",x"231a10",x"241911",x"21170f",x"241911",x"21180f",x"21170f",x"241a11",x"241b11",x"241a11",x"231910",x"21180f",x"231910",x"241911",x"261b11",x"231a10",x"21180f",x"241a11",x"241a11",x"241a11",x"241910",x"241911",x"241a11",x"251a12",x"251b11",x"21170f",x"231810",x"1f170e",x"1f170e",x"1d150d",x"21180f",x"20170e",x"22190f",x"231910",x"251b12",x"251b12",x"271c14",x"241a12",x"261c13",x"281f16",x"281e15",x"281e15",x"271d14",x"241c14",x"251c14",x"261c14",x"241b13",x"251b12",x"221a11",x"241b11",x"211810",x"22190f",x"1b130b",x"1f160d",x"20160d",x"20160d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1c0f",x"2f1c0f",x"3a2111",x"27150b",x"3d2311",x"3b2311",x"3b2311",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"1c1108",x"150e07",x"24150a",x"1e1208",x"211409",x"25160a",x"26160a",x"2a180b",x"29180b",x"2b190b",x"29180b",x"25160a",x"25160a",x"24150a",x"2a180b",x"29180b",x"24150a",x"27160a",x"29170a",x"251509",x"221409",x"251409",x"1d1108",x"211309",x"241409",x"201308",x"231409",x"1c1108",x"241509",x"201208",x"241509",x"231409",x"231509",x"27160a",x"25160a",x"26160a",x"2a180b",x"221409",x"231409",x"27160a",x"241509",x"28170a",x"28170a",x"201309",x"27170a",x"25150a",x"27160a",x"27160a",x"211309",x"26160a",x"26160a",x"1b1108",x"26160a",x"221409",x"25150a",x"27160a",x"26180c",x"20140b",x"25160d",x"1d140c",x"1d140c",x"1d140c",x"391f0b",x"341c0b",x"3f240f",x"351e0e",x"301b0c",x"351d0d",x"371f0e",x"38200e",x"351d0d",x"38200f",x"221509",x"28180b",x"2b190b",x"201912",x"1d1610",x"19120c",x"150e07",x"1c1108",x"1c1108",x"24160a",x"1e1209",x"25150a",x"25160a",x"24150a",x"180f07",x"1e1209",x"24150a",x"27170a",x"26160a",x"2b190c",x"221409",x"2a180b",x"211309",x"211409",x"2a190b",x"28170b",x"231509",x"26160a",x"28170a",x"231409",x"28180b",x"25160a",x"27170a",x"29180b",x"27170a",x"27170b",x"27170a",x"24150a",x"27170a",x"27170b",x"26160a",x"2a190b",x"24150a",x"24150a",x"27170a",x"27170a",x"27160a",x"28170a",x"27160a",x"26160a",x"261509",x"1f1208",x"221309",x"211309",x"1f1208",x"1d1108",x"241509",x"26160a",x"27160a",x"201309",x"211308",x"251509",x"241509",x"241509",x"28190c",x"2b1b0f",x"2d1c10",x"2d1d12",x"261a11",x"201710",x"4e2e16",x"3d2411",x"371f0d",x"381f0e",x"412612",x"3f2411",x"432813",x"412511",x"3b2210",x"351d0d",x"3e2411",x"170f07",x"24150a",x"29180b",x"3e2515",x"292019",x"191008",x"1c1108",x"22150b",x"2d1b0e",x"372f27",x"544b41",x"544b41",x"000000",x"000000",x"000000",x"000000"),
(x"866c55",x"866b54",x"5e5246",x"564a3f",x"514438",x"4a3c2f",x"4c3f33",x"483a2d",x"483a2e",x"463a2e",x"46382c",x"46392d",x"44372b",x"493b2f",x"4b3d32",x"4d4034",x"4e4033",x"524234",x"4d3f31",x"514133",x"514235",x"544436",x"554435",x"524233",x"4c3d2f",x"4b3c2e",x"4d3c2d",x"49392c",x"4d3e2f",x"4e3f32",x"4f3f30",x"4c3c2e",x"503e2f",x"4b3b2d",x"4b3b2d",x"4a3a2c",x"4c3b2d",x"4d3d2f",x"4c3b2c",x"524132",x"514032",x"4e3d2e",x"544232",x"544231",x"524132",x"524131",x"503e2e",x"4d3d2f",x"503e30",x"4e3d2f",x"503f31",x"513f2f",x"514031",x"4d3e30",x"4c3c2e",x"47382b",x"4a3a2b",x"4e3d30",x"503e2e",x"4b3c2f",x"4c3c2f",x"4b3c2e",x"4b3b2e",x"493a2d",x"493a2d",x"45372a",x"46382b",x"47392d",x"4c3c2e",x"4c3c2e",x"483a2c",x"493a2c",x"43362b",x"4a3c30",x"4a3c2f",x"473a2f",x"493b2f",x"4c3d31",x"483b30",x"4e4135",x"53453a",x"57493d",x"615143",x"615143",x"241c15",x"231c14",x"271f17",x"231c15",x"201911",x"221a13",x"201811",x"201811",x"211910",x"1f160d",x"1d140b",x"1c130a",x"25190f",x"24190e",x"1f150b",x"21170d",x"20160c",x"291d11",x"2a1d12",x"2a1d11",x"271a0f",x"291c10",x"2a1d11",x"2a1d11",x"2b1e11",x"2f2013",x"2b1d11",x"302114",x"302114",x"312215",x"322316",x"382717",x"3a2818",x"3a2a1a",x"382718",x"382718",x"362618",x"372718",x"3e2c1c",x"3b2a1a",x"382819",x"372618",x"3e2c1c",x"382819",x"3a291a",x"3c2a1a",x"3a2819",x"3e2c1c",x"3a2a1b",x"453222",x"443323",x"453425",x"423223",x"433323",x"443324",x"413123",x"57402e",x"211a14",x"231a11",x"1f150c",x"1d130a",x"1d140b",x"1d140b",x"20160b",x"20160c",x"261a0f",x"23180d",x"23170d",x"22170d",x"24190e",x"23180d",x"24180e",x"24180e",x"281b10",x"23180d",x"281b10",x"281c10",x"291c11",x"23180d",x"291c11",x"2a1d11",x"2e2013",x"2e2114",x"2c1f13",x"291d10",x"2e1f13",x"312214",x"2c1e12",x"322315",x"2c1f12",x"2d1f13",x"322215",x"2a1d11",x"302114",x"312215",x"362516",x"312214",x"2f2114",x"312215",x"322315",x"2d1f13",x"312215",x"342416",x"322315",x"342417",x"352517",x"382718",x"392819",x"43301f",x"523a26",x"150e07",x"312215",x"332416",x"342517",x"39291a",x"3c2a1b",x"150e07",x"150e07",x"150e07",x"181008",x"191109",x"181008",x"181008",x"1d130a",x"181008",x"1d140b",x"1b130b",x"1f160d",x"21180f",x"221810",x"20180f",x"20180f",x"211810",x"23180f",x"20180f",x"231810",x"221810",x"231810",x"20180f",x"20170d",x"21180e",x"1f150c",x"20170d",x"21170e",x"21180e",x"23190f",x"22180f",x"22180f",x"20160d",x"21180e",x"21180e",x"20170d",x"21170e",x"20170d",x"20170d",x"21170d",x"21170d",x"21170e",x"21180f",x"21180d",x"21180e",x"21180f",x"21170e",x"21170e",x"1f160d",x"21170e",x"21180e",x"21170e",x"20170e",x"21170e",x"231910",x"22180f",x"251a11",x"22190f",x"241b12",x"261c12",x"241b11",x"271d14",x"271d14",x"261c13",x"241b13",x"241b12",x"231a11",x"221911",x"221a11",x"20170e",x"20170f",x"1f150c",x"1f150c",x"20150c",x"1e140b",x"1d140a",x"1d140b",x"1d140b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1b0e",x"2d1b0e",x"382111",x"27150b",x"3b2312",x"402511",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"1f1309",x"211409",x"1e1209",x"150e07",x"150e07",x"150e07",x"180f08",x"180f07",x"191008",x"150e07",x"180f08",x"26170b",x"191008",x"160e07",x"160f07",x"160e07",x"1e1209",x"180f08",x"191008",x"150e07",x"150e07",x"150e07",x"1c1108",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"150e07",x"170f07",x"150e07",x"170f07",x"170f07",x"1a1008",x"1d1208",x"1b1108",x"150e07",x"170f07",x"1c1108",x"1e1208",x"150e07",x"1c1108",x"150e07",x"150e07",x"1d1108",x"1b1008",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"1d1108",x"2a180b",x"28180c",x"29190c",x"23150b",x"1b120a",x"1b120a",x"391e0a",x"41230e",x"3e240f",x"351f0f",x"28170a",x"361e0d",x"381f0e",x"3d220f",x"301b0c",x"361f0e",x"23150a",x"28180b",x"321d0d",x"201913",x"1e1811",x"1c150f",x"17110a",x"1e1108",x"1d1108",x"180f08",x"180f08",x"1c1108",x"221409",x"24150a",x"150e07",x"150e07",x"201309",x"1e1209",x"241509",x"1e1208",x"25160a",x"150e07",x"1e1309",x"24160a",x"1e1209",x"1e1208",x"211409",x"241509",x"28180b",x"29180b",x"24150a",x"231509",x"211409",x"211409",x"1f1309",x"201309",x"25160a",x"25160a",x"1e1209",x"23150a",x"26170a",x"221409",x"211409",x"22140a",x"211409",x"211409",x"221409",x"25150a",x"221409",x"1d1108",x"241509",x"221409",x"1f1208",x"201308",x"1d1108",x"1e1108",x"1f1209",x"241509",x"241509",x"251509",x"26160a",x"25160a",x"211409",x"211409",x"26170b",x"301d0f",x"2d1d11",x"2f1e11",x"2a1c11",x"23170f",x"4a2a14",x"3f2511",x"38200e",x"381f0e",x"3e2511",x"361f0e",x"422713",x"3b2210",x"412612",x"351e0d",x"38210f",x"170f07",x"23150a",x"28180b",x"3f2615",x"2e241c",x"191008",x"1c1108",x"22150b",x"2f1c0f",x"3c332a",x"564c42",x"564c42",x"000000",x"000000",x"000000",x"000000"),
(x"8a6f56",x"876e54",x"5d5043",x"54473b",x"524539",x"483b2f",x"4d3e31",x"4a3d31",x"4c3d2e",x"4b3d30",x"4b3d30",x"4a3c2f",x"483a2d",x"4a3b2e",x"493b2e",x"4e3f32",x"4f3f32",x"4f4134",x"504032",x"514132",x"544435",x"594737",x"524133",x"524132",x"4d3d2f",x"4d3c2d",x"503e2f",x"4d3d2f",x"503e2f",x"514030",x"514131",x"4f3e2f",x"503f30",x"524130",x"514131",x"514333",x"564534",x"564332",x"524030",x"513f30",x"574434",x"564433",x"5d4938",x"564334",x"554333",x"4f3e2f",x"524131",x"554231",x"544335",x"4f3f30",x"514031",x"4e3d2e",x"534131",x"564333",x"544131",x"544231",x"544332",x"503f31",x"4e3d2f",x"4f3e30",x"4d3c2d",x"4f3e2d",x"503f2f",x"4d3d2f",x"4f3e2f",x"4e3e30",x"514131",x"4c3e2f",x"504031",x"4a3b2c",x"4b3c2e",x"4d3d2f",x"504032",x"503f32",x"4f4032",x"4f4032",x"504234",x"504134",x"4c3f32",x"504135",x"584a3d",x"5c4e41",x"645446",x"655446",x"271e16",x"281f17",x"231b14",x"271e15",x"211a12",x"221a13",x"251c14",x"201911",x"221910",x"1b130b",x"1e150b",x"21160c",x"23180e",x"23190e",x"241a0f",x"271d11",x"2d2014",x"2c1f13",x"2d1f13",x"2a1e12",x"302215",x"2f2114",x"342518",x"312216",x"332417",x"342516",x"322315",x"342416",x"362618",x"352517",x"342416",x"342315",x"3a2818",x"3a2a1b",x"382718",x"382819",x"3c2a1b",x"392819",x"3c2a1b",x"422f1e",x"3c2a1b",x"42301f",x"44311f",x"412e1d",x"402d1c",x"402f1e",x"413120",x"423322",x"433122",x"483626",x"473525",x"483727",x"493828",x"463526",x"4a3829",x"4a3829",x"644b35",x"231c16",x"211910",x"1d140b",x"1e150b",x"1e150c",x"20160c",x"1e140b",x"23170d",x"21170d",x"23180e",x"261a0f",x"261a0f",x"23180e",x"251a0f",x"2a1d11",x"251a0f",x"24190e",x"261a0f",x"2b1e12",x"2b1e12",x"2a1d11",x"2d2114",x"2f2316",x"312417",x"302215",x"2e2114",x"2d2013",x"322316",x"2f2114",x"312316",x"352618",x"352618",x"382819",x"2c1e12",x"362618",x"332416",x"39281a",x"2e2013",x"2d1f12",x"2e1f12",x"362819",x"362617",x"362618",x"3a291a",x"332416",x"392819",x"352517",x"392819",x"392819",x"3b2a1b",x"392819",x"473322",x"5b432c",x"150e07",x"372a1b",x"37281a",x"39291a",x"3b2a1b",x"3d2c1d",x"150e07",x"150e07",x"150e07",x"1e150c",x"191109",x"191109",x"1d140b",x"191109",x"21170d",x"191109",x"1d140b",x"1e150d",x"1e160c",x"20170e",x"23180e",x"22190f",x"23180f",x"20160d",x"21180e",x"20170e",x"20160d",x"23190f",x"23180f",x"23180e",x"20160d",x"23190f",x"20180e",x"231a10",x"241b11",x"261b11",x"23190f",x"23180f",x"231a10",x"23180f",x"23190f",x"20170e",x"23190f",x"22180f",x"21180e",x"21180e",x"23190f",x"22180f",x"21170e",x"20170d",x"22170d",x"23190f",x"20160d",x"20170d",x"20160d",x"21180e",x"21180e",x"23190f",x"23180f",x"23190f",x"23180f",x"23180e",x"23180f",x"22180f",x"251b12",x"241b11",x"251b11",x"251b11",x"241a11",x"251a10",x"221910",x"241910",x"241a12",x"211910",x"21180f",x"20160d",x"21180e",x"1d140b",x"1e150b",x"1e150b",x"1e140b",x"1f150b",x"1c130a",x"1c130a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e1c10",x"2e1c10",x"351f11",x"27150c",x"3a2312",x"422713",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"25150a",x"1a1008",x"27170a",x"311b0c",x"321c0d",x"331d0d",x"371f0e",x"311c0d",x"301c0d",x"331c0d",x"311c0d",x"321d0d",x"311c0c",x"331d0d",x"361f0f",x"301b0c",x"2e1b0c",x"331d0d",x"301b0b",x"2f1a0a",x"2f1a0b",x"331c0c",x"311c0b",x"331c0c",x"301b0b",x"321c0c",x"2c190b",x"341c0d",x"2f1a0b",x"2c190b",x"2f1a0b",x"2e1a0b",x"271509",x"28170a",x"2f1b0c",x"2c190b",x"341d0d",x"301b0b",x"301b0c",x"2f1a0c",x"301b0c",x"301b0c",x"311c0c",x"2f1a0c",x"311c0c",x"29170a",x"2e1a0b",x"2e190b",x"2f1a0b",x"2e1a0b",x"2c190b",x"311c0c",x"321c0d",x"331c0d",x"331d0d",x"2f1b0c",x"321c0d",x"150e07",x"261509",x"2a180a",x"27160a",x"23150b",x"22150b",x"22150b",x"4c2c14",x"4c2c14",x"38200f",x"2d1a0c",x"25150a",x"371f0e",x"371f0e",x"3a200e",x"341d0d",x"39210f",x"231509",x"25160a",x"321d0d",x"211b14",x"1f1912",x"1b150e",x"1c120b",x"1e1208",x"1d1208",x"201309",x"1e1208",x"211309",x"241509",x"25160a",x"221409",x"211309",x"221309",x"221509",x"241509",x"221409",x"23150a",x"221409",x"211409",x"211409",x"221409",x"25170a",x"24160a",x"27170b",x"29190b",x"24160a",x"23170b",x"25170a",x"211409",x"211409",x"24160a",x"24160a",x"1e1209",x"231409",x"1d1208",x"1d1209",x"201309",x"231509",x"1f1309",x"201409",x"231509",x"1b1108",x"201309",x"1c1108",x"201309",x"1f1309",x"1e1208",x"1b1108",x"160e07",x"170f07",x"170f08",x"1f1309",x"1f1309",x"1d1208",x"1c1108",x"1f1209",x"191008",x"1a1008",x"1b1108",x"1e1209",x"1c1109",x"29190d",x"352011",x"332012",x"2d1d11",x"281a0f",x"492a13",x"3e2411",x"3f2410",x"3f2311",x"442814",x"3d2410",x"402612",x"3c220f",x"3b220f",x"331c0c",x"3f2411",x"180f07",x"24150a",x"27170b",x"3f2616",x"342a21",x"191008",x"1c1108",x"21150b",x"2e1c10",x"372f27",x"564c42",x"564c42",x"000000",x"000000",x"000000",x"000000"),
(x"8c7058",x"8d7058",x"5c4f42",x"504336",x"493b2e",x"45382b",x"463a2d",x"493b2e",x"463a2e",x"473a2d",x"4a3c2f",x"44382d",x"493b2f",x"4a3c2f",x"4c3d2f",x"504031",x"524133",x"554434",x"554435",x"584737",x"534335",x"504134",x"504032",x"524132",x"4e3e2f",x"523f2e",x"524131",x"544131",x"544233",x"503e30",x"4f3d2e",x"523f2e",x"52402f",x"503e2f",x"52402f",x"503d2e",x"554232",x"524030",x"554333",x"584535",x"514131",x"514132",x"574535",x"564333",x"554231",x"524030",x"584534",x"544333",x"564334",x"574535",x"544233",x"5e4a38",x"574535",x"4f3f32",x"544131",x"4f3e31",x"524133",x"534231",x"4d3d2f",x"524030",x"503f30",x"4b3c2e",x"4e3e2f",x"4d3c2e",x"504031",x"4d3d2e",x"514031",x"4d3d2f",x"554435",x"4c392a",x"4e3f32",x"4d3d2f",x"4e4033",x"504133",x"504234",x"4d3f32",x"4c3d2f",x"4a3b2d",x"4c3e31",x"4f4135",x"514134",x"5b4d40",x"655648",x"665648",x"241c15",x"221b14",x"231c14",x"231c15",x"251d15",x"211912",x"241c14",x"241b13",x"231a11",x"1b130b",x"21160d",x"1e140b",x"21170d",x"24180e",x"24190f",x"261a0f",x"271b10",x"2c1e12",x"2c1f13",x"2f2114",x"2a1f13",x"302215",x"2f2214",x"2f2114",x"312215",x"352617",x"332416",x"362719",x"372718",x"3a2a1a",x"382719",x"392819",x"39281a",x"362517",x"382718",x"382718",x"3a2819",x"3a2819",x"362618",x"3b291a",x"3f2d1d",x"3c2a1a",x"3f2d1c",x"402d1d",x"412e1d",x"44301f",x"453220",x"433120",x"463424",x"413021",x"443425",x"483626",x"433425",x"463627",x"493827",x"443425",x"604732",x"201a13",x"241a10",x"21170d",x"20160c",x"1e150b",x"21160d",x"1e150b",x"21160d",x"1f150c",x"25190f",x"25190e",x"291c10",x"25190f",x"24190e",x"2a1d11",x"261b10",x"25190e",x"2d2013",x"2b1e12",x"2c1f12",x"2c1f12",x"2c1f13",x"2f2114",x"342517",x"2a1d11",x"302215",x"332517",x"2e2214",x"2f2215",x"2d2013",x"342416",x"362719",x"332416",x"362718",x"302216",x"332416",x"362618",x"342416",x"352517",x"382719",x"2f2014",x"2e2013",x"312214",x"332316",x"382718",x"362617",x"382718",x"362718",x"362617",x"382819",x"39281a",x"4d3825",x"59412b",x"150e07",x"382719",x"382819",x"332416",x"39291a",x"3b2a1b",x"150e07",x"150e07",x"150e07",x"191109",x"191109",x"1e150b",x"191109",x"21170d",x"191109",x"1e150b",x"1e140b",x"1e150b",x"1e140b",x"1d130b",x"20160c",x"1d140b",x"20160c",x"1d140b",x"1d140b",x"20160c",x"21170d",x"1d140b",x"1e140b",x"21160d",x"21170d",x"21170d",x"21170d",x"23180e",x"251a0f",x"20160c",x"24190f",x"21170d",x"20160d",x"24190f",x"21170d",x"21160d",x"24190e",x"21170d",x"21170d",x"21170d",x"20160c",x"21170d",x"21160c",x"21170d",x"21160d",x"1f150c",x"1d140b",x"20160c",x"1d140b",x"1d140b",x"20150c",x"20160c",x"24190e",x"20160c",x"21160d",x"21160c",x"21170d",x"24190e",x"24190e",x"21160d",x"22170d",x"20160c",x"21170d",x"22170d",x"1d140b",x"21170d",x"1e150b",x"21160d",x"1e150b",x"1e150b",x"1e150b",x"1e150c",x"1e140b",x"1e150b",x"1e140b",x"1e150b",x"1e140b",x"1e140b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1b0f",x"2d1b0f",x"362012",x"26160c",x"382212",x"402512",x"150e07",x"150e07",x"150e07",x"180f07",x"1d1108",x"1b1008",x"1c1108",x"2e1a0b",x"321c0d",x"321c0c",x"311b0c",x"351d0d",x"2e1a0b",x"311b0c",x"321c0c",x"351e0d",x"311b0c",x"351e0d",x"341d0d",x"3a200f",x"3b200e",x"3b210f",x"381f0e",x"3b210e",x"371f0d",x"361e0d",x"381f0e",x"321b0c",x"341d0d",x"341d0c",x"2c170a",x"2f1a0b",x"331c0c",x"351e0d",x"351d0d",x"321c0c",x"331c0c",x"331c0c",x"311c0c",x"331c0d",x"321c0c",x"2f1a0b",x"2f190b",x"2d190b",x"311b0c",x"361e0d",x"311b0b",x"311b0b",x"311b0b",x"341d0d",x"361e0d",x"311b0b",x"30190b",x"311b0b",x"321b0b",x"311b0b",x"321b0c",x"331c0c",x"321c0c",x"301a0b",x"2d190b",x"311b0b",x"150e07",x"211309",x"27160a",x"2d190b",x"24160b",x"22150b",x"22150b",x"4d2d15",x"4d2d15",x"3b2210",x"331d0d",x"2c190b",x"371f0e",x"3d220f",x"331e0d",x"371f0e",x"3b220f",x"231509",x"25160a",x"351f0e",x"211b14",x"1f1912",x"1d1610",x"1e130a",x"231409",x"241509",x"311c0c",x"321c0d",x"311b0d",x"361f0e",x"3a210f",x"351d0d",x"351e0d",x"2e1a0b",x"2f1a0b",x"351e0d",x"321c0c",x"2f1b0c",x"311b0c",x"2d190b",x"2b170a",x"2e190b",x"2e1a0b",x"2f1a0b",x"311b0c",x"301a0b",x"331c0c",x"381f0e",x"351e0d",x"351e0d",x"381f0e",x"341d0d",x"39200e",x"361e0d",x"341d0d",x"331d0d",x"311c0c",x"321c0c",x"341d0d",x"371e0d",x"38200e",x"361e0d",x"361e0d",x"361e0d",x"361e0d",x"351d0d",x"361e0d",x"351e0d",x"2d190b",x"371e0d",x"321b0b",x"2e190a",x"311b0b",x"331c0c",x"341d0d",x"381f0e",x"2f1a0c",x"351e0d",x"311b0b",x"341d0d",x"341d0d",x"160e07",x"24160b",x"28180d",x"2e1c10",x"2c1b10",x"261a10",x"512f16",x"3e2411",x"3d2310",x"3f2512",x"3f2512",x"412612",x"442813",x"3c2411",x"3e2310",x"371f0e",x"39200f",x"180f07",x"23150a",x"26160a",x"3d2515",x"31261d",x"191008",x"1d1208",x"23150b",x"2f1d10",x"3c342d",x"52493e",x"52493e",x"000000",x"000000",x"000000",x"000000"),
(x"8d7158",x"8c7159",x"5d5045",x"524539",x"473a2d",x"423529",x"45382c",x"4b3d30",x"47382b",x"473a2d",x"493a2d",x"48382b",x"46382c",x"4a392b",x"4c3c2e",x"49392a",x"514133",x"554434",x"544334",x"544537",x"564637",x"584636",x"4f3f30",x"544231",x"513f31",x"564333",x"534232",x"584636",x"584535",x"574434",x"524030",x"52402f",x"503f30",x"554232",x"564334",x"544130",x"554230",x"574333",x"544233",x"574534",x"574333",x"594634",x"594736",x"584535",x"534132",x"594635",x"544233",x"594736",x"5a4736",x"5a4737",x"5d4a3a",x"5c4938",x"564334",x"594737",x"574637",x"524131",x"544334",x"554435",x"524132",x"534233",x"5a4635",x"544335",x"504032",x"514031",x"514132",x"504032",x"514132",x"4c3d30",x"4c3c2d",x"4f3f31",x"4d3d30",x"514134",x"4d3d30",x"504134",x"4e4032",x"4e3f31",x"504032",x"4b3d2f",x"4d3d2f",x"4f3f31",x"544538",x"5b4c3f",x"665646",x"645444",x"271e16",x"271e16",x"261e16",x"221b14",x"241b13",x"211912",x"261d15",x"231b12",x"231a11",x"20170e",x"20160c",x"24180e",x"21170d",x"24190f",x"251a0f",x"291c11",x"251a0f",x"302114",x"2c1f12",x"2a1e12",x"2e2013",x"332416",x"312316",x"302215",x"352618",x"362718",x"382718",x"382718",x"3a281a",x"3d2b1c",x"39281a",x"392819",x"3b291a",x"3a2a1a",x"3d2b1b",x"3b2a1a",x"392819",x"3f2d1c",x"3d2b1c",x"3e2d1d",x"3c2a1b",x"443120",x"402d1c",x"402e1d",x"443120",x"412f1f",x"443120",x"453120",x"453222",x"463323",x"433122",x"4b3828",x"463424",x"453425",x"4d3a29",x"4b3827",x"644b34",x"1f1811",x"21180f",x"1e140b",x"1e140b",x"1e140b",x"21170d",x"21170d",x"23180e",x"24190e",x"23180d",x"251a0f",x"25190e",x"261a0f",x"261a0f",x"271b10",x"2c1f12",x"2c1f13",x"291c10",x"2c1e12",x"2c1f13",x"302215",x"2d2014",x"332416",x"2f2114",x"302114",x"2e2013",x"312216",x"302215",x"332416",x"312316",x"332416",x"352618",x"362718",x"352517",x"382718",x"342416",x"3b2a1b",x"352518",x"362618",x"2f2114",x"352517",x"342516",x"312215",x"3a2819",x"382819",x"342517",x"3d2b1c",x"3f2d1d",x"3b2a1b",x"372718",x"372718",x"4d3926",x"5d442e",x"150e07",x"352517",x"372718",x"3b2a1b",x"372718",x"3d2c1c",x"150e07",x"150e07",x"150e07",x"191109",x"191109",x"191109",x"191109",x"21160c",x"1e140b",x"21160d",x"1e150c",x"261a0f",x"21160c",x"261b10",x"20160c",x"20160c",x"20160c",x"1e140b",x"24190e",x"1e150c",x"21160d",x"1f150c",x"20160c",x"21160d",x"21170d",x"24190f",x"25190f",x"20160c",x"20160c",x"23180e",x"20160c",x"24190f",x"21170d",x"21170d",x"22170d",x"24190e",x"24190f",x"24190e",x"23180e",x"21160c",x"24180e",x"24180e",x"21170d",x"21170d",x"21160c",x"24190e",x"23180d",x"20160c",x"23180d",x"24180e",x"21160d",x"24190f",x"261a0f",x"2b1f13",x"23180d",x"24180e",x"24190f",x"271b10",x"25190f",x"23180e",x"20160c",x"23180e",x"20160c",x"24190f",x"271b10",x"21170d",x"22170d",x"24190e",x"21170d",x"1e150b",x"21160c",x"21160c",x"21160d",x"1e140b",x"21170d",x"1e150b",x"1e140b",x"1e140b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1c10",x"2d1c10",x"372112",x"2e1a0e",x"382111",x"3d2311",x"160e07",x"160e07",x"150e07",x"1b1108",x"1f1309",x"24150a",x"241509",x"2e1a0b",x"331d0d",x"321d0d",x"361f0e",x"361f0e",x"3d2310",x"38200e",x"3c230f",x"38200e",x"3d2310",x"39200f",x"37200e",x"3b210f",x"3a200e",x"3a1f0e",x"3a210f",x"3d230f",x"3e2310",x"3c2310",x"38200e",x"371f0e",x"371f0e",x"39200f",x"371f0e",x"38200e",x"39200e",x"38200e",x"351d0d",x"351d0d",x"341d0d",x"301b0b",x"361e0d",x"341d0c",x"351d0d",x"331c0c",x"341d0c",x"321c0c",x"351e0d",x"3a200f",x"38200e",x"361e0d",x"381f0e",x"381f0e",x"39200e",x"371f0e",x"331c0c",x"321b0b",x"341d0c",x"351d0c",x"321c0c",x"311b0c",x"331c0c",x"341c0c",x"301a0b",x"2a170a",x"150e07",x"201309",x"26160a",x"221409",x"23150b",x"1f130a",x"1f130a",x"4b2b15",x"4b2b15",x"39210f",x"331d0d",x"2f1a0c",x"361f0e",x"371f0e",x"341c0d",x"3a200f",x"3a210e",x"231509",x"27170b",x"331d0e",x"221b14",x"201912",x"1d1710",x"24170d",x"25150a",x"26160a",x"311b0c",x"321c0c",x"301b0c",x"331d0d",x"39200f",x"331d0d",x"3a210f",x"39200f",x"361e0e",x"3c220f",x"38200e",x"3a210f",x"311c0c",x"351e0d",x"321d0d",x"2f1b0c",x"351e0d",x"351e0e",x"341e0d",x"3a210f",x"3a200f",x"371f0e",x"381f0e",x"3b220f",x"371f0e",x"38200f",x"371f0e",x"38200f",x"3a210f",x"3e2310",x"361e0e",x"39200f",x"3a210f",x"38200e",x"351e0d",x"341d0c",x"351d0d",x"3a210f",x"3a210f",x"3c2210",x"371f0e",x"38200e",x"361f0e",x"3b220f",x"351d0d",x"38200e",x"371f0e",x"361e0d",x"371f0d",x"371f0d",x"371f0d",x"351d0c",x"321c0c",x"311b0c",x"321c0c",x"160e07",x"25160b",x"2d1b0f",x"2d1c11",x"2d1c10",x"23180f",x"4d2c15",x"3e2411",x"39200e",x"432713",x"3b210f",x"412712",x"432813",x"3b2210",x"3b2210",x"3a210f",x"39210f",x"170f07",x"23150a",x"24150a",x"3d2515",x"30271f",x"191008",x"1d1108",x"23150b",x"2d1c0f",x"352d25",x"554c41",x"554c41",x"000000",x"000000",x"000000",x"000000"),
(x"8b6f57",x"8e7159",x"5e5145",x"514438",x"4c3f34",x"46392d",x"48392d",x"42362a",x"46382b",x"4a3b2e",x"483a2d",x"48392c",x"45372b",x"473a2d",x"4f3f30",x"513f31",x"514133",x"4f3f31",x"554233",x"534132",x"564435",x"554333",x"503f31",x"4d3d2e",x"513f2f",x"4d3d2e",x"513f2f",x"524132",x"524131",x"544132",x"523f2f",x"4f3d2d",x"534030",x"584331",x"584331",x"564232",x"574331",x"574533",x"5d4837",x"5a4533",x"5b4836",x"574534",x"554232",x"564333",x"564333",x"564433",x"544233",x"5a4735",x"5b4737",x"5b4736",x"5c4939",x"5a4737",x"5c4a3a",x"5c4938",x"564637",x"564435",x"544336",x"564535",x"554334",x"534233",x"524132",x"544335",x"524232",x"534335",x"594737",x"564536",x"554435",x"514031",x"514031",x"504133",x"544334",x"534133",x"544336",x"524233",x"504032",x"524234",x"4d3e31",x"4b3c2e",x"4a3b2e",x"4c3d30",x"56473a",x"574739",x"635141",x"625142",x"241c14",x"251d15",x"241c14",x"241c14",x"241b13",x"241c13",x"231a12",x"221911",x"20180f",x"1e140b",x"23180e",x"23180e",x"21170d",x"24190e",x"2a1d12",x"2a1d11",x"2a1d11",x"2d1f13",x"302215",x"2d2013",x"2f2115",x"372719",x"322316",x"352517",x"332416",x"362618",x"3a291a",x"392819",x"382819",x"362617",x"392819",x"382718",x"3c2a1a",x"3a2919",x"372618",x"352416",x"372618",x"392819",x"3a2919",x"3d2b1c",x"3b2a1a",x"3f2d1c",x"412f1e",x"432f1e",x"422f1e",x"43301f",x"453220",x"433120",x"463222",x"4b3726",x"4a3827",x"473524",x"473526",x"473626",x"483625",x"4a3827",x"634a33",x"1d1710",x"20160d",x"1e140b",x"1e150b",x"1d140b",x"20160c",x"1d140b",x"20160c",x"25190e",x"23180d",x"22170d",x"23180d",x"271b10",x"281c10",x"291c11",x"2d1f12",x"291c11",x"291d11",x"291c11",x"2c1f12",x"302215",x"2e2114",x"2c1f13",x"322316",x"2f2115",x"352518",x"2f2114",x"312316",x"312316",x"2d2013",x"362718",x"392819",x"372819",x"362617",x"332416",x"3a291a",x"342416",x"342416",x"332315",x"352517",x"322315",x"332415",x"312214",x"2e2013",x"322316",x"3b291a",x"3b2a1b",x"3a2919",x"3a291a",x"3a291a",x"3a291a",x"4e3825",x"59412c",x"150e07",x"352517",x"382819",x"3c2b1c",x"372719",x"39281a",x"150e07",x"150e07",x"150e07",x"1e150b",x"21170d",x"1f150c",x"23180e",x"20160c",x"1e140b",x"1d140b",x"23170d",x"22170d",x"24190e",x"281b10",x"21170c",x"20150c",x"21160c",x"24190e",x"23180d",x"291c11",x"251a0f",x"251a0f",x"21160d",x"291c11",x"261a0f",x"24190f",x"24190f",x"24190e",x"261a0f",x"25190f",x"2b1e13",x"261a0f",x"2b1e12",x"2b1e13",x"291d11",x"2a1d11",x"271b10",x"22170d",x"23180e",x"23180d",x"261a0f",x"23180d",x"281b10",x"281b10",x"22170d",x"22170d",x"23180d",x"22170d",x"23180d",x"271b10",x"23180d",x"291c11",x"20160c",x"2b1e12",x"23180e",x"261a0f",x"2c1f12",x"24190f",x"2a1d12",x"261b10",x"21160d",x"25190f",x"251a0f",x"21160d",x"24190f",x"251a0f",x"23180e",x"24190e",x"24190f",x"22170d",x"21160c",x"251a0f",x"21160d",x"20160c",x"25190e",x"20150c",x"20160c",x"20160c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1c10",x"2d1c10",x"362012",x"2e1a0e",x"362011",x"3d2310",x"150e07",x"150e07",x"150e07",x"1f1208",x"1d1208",x"211309",x"221409",x"2f1b0c",x"351f0e",x"341d0d",x"361f0e",x"361f0e",x"39200f",x"381f0e",x"351d0d",x"371f0e",x"3b200e",x"371f0e",x"3d2310",x"3a210f",x"3c210f",x"371e0d",x"371e0d",x"39200e",x"3b200e",x"3b220f",x"39200f",x"351e0d",x"341d0c",x"331c0c",x"361e0d",x"381f0e",x"341c0d",x"351d0d",x"361e0d",x"321b0c",x"311b0b",x"311a0b",x"311a0b",x"2f190a",x"2f190b",x"2f1a0b",x"311b0c",x"341d0c",x"301b0b",x"301a0b",x"30190b",x"321b0b",x"341c0c",x"361d0c",x"351d0d",x"331c0c",x"331c0c",x"331c0b",x"2e180a",x"311a0b",x"301a0b",x"2d180a",x"321b0b",x"311a0b",x"311a0b",x"28160a",x"150e07",x"201208",x"28160a",x"2a180b",x"27160a",x"231409",x"231409",x"472812",x"472812",x"3c2310",x"331d0d",x"2e1b0c",x"3a210f",x"311c0d",x"3a210f",x"39200e",x"361e0d",x"24150a",x"28180b",x"341e0e",x"221c15",x"211a14",x"1f1710",x"25160b",x"26160a",x"25150a",x"311b0c",x"301b0c",x"2e1a0c",x"341d0d",x"331d0d",x"341d0d",x"351e0d",x"38200e",x"371f0e",x"351d0d",x"341d0c",x"371e0d",x"311b0c",x"311b0b",x"321c0c",x"311b0c",x"2c180a",x"2f1a0b",x"371e0e",x"39200f",x"3a210f",x"39210f",x"39200f",x"361e0d",x"3a210f",x"381f0e",x"371f0e",x"331c0c",x"371f0e",x"371f0e",x"2f1b0c",x"351e0d",x"3c220f",x"3a210f",x"381f0d",x"361d0d",x"331c0d",x"361e0d",x"39200e",x"3a210f",x"39210f",x"38200e",x"361e0d",x"381f0e",x"39200e",x"39200e",x"361e0d",x"351e0d",x"351e0d",x"351d0d",x"311b0b",x"2e190b",x"2f1a0b",x"311b0b",x"2e190a",x"150e07",x"25170b",x"29190e",x"2f1d11",x"2a1c11",x"25180f",x"4f2e16",x"412511",x"3b210f",x"402511",x"341d0d",x"412613",x"392110",x"39200f",x"3a210f",x"39200f",x"3a2210",x"170f07",x"22150a",x"25160a",x"3f2717",x"352a22",x"191008",x"1c1108",x"23150b",x"2f1d11",x"382f27",x"564c42",x"564c42",x"000000",x"000000",x"000000",x"000000"),
(x"856b53",x"856b54",x"5a4e41",x"54483c",x"463a30",x"44392f",x"43362a",x"433529",x"47392c",x"43362a",x"47382c",x"46392e",x"433629",x"483a2c",x"4b3b2e",x"504133",x"514234",x"4c3c2e",x"4c3b2c",x"4b3c2d",x"4f3f31",x"514131",x"554233",x"554333",x"554332",x"524132",x"574333",x"554232",x"554232",x"554230",x"534030",x"503d2d",x"53402f",x"54402e",x"523f2d",x"564230",x"503c2b",x"513c2c",x"574330",x"5c4633",x"554232",x"5a4635",x"544132",x"564333",x"544131",x"544232",x"524131",x"574332",x"584433",x"594535",x"584535",x"594737",x"5b4939",x"5c4a3a",x"5e4a38",x"624d3b",x"594736",x"544233",x"5b4737",x"5a4737",x"594635",x"564433",x"564536",x"554536",x"544334",x"524132",x"554434",x"4e4032",x"47392c",x"4c3c2f",x"514032",x"4f3f32",x"4b3b2e",x"4d3e30",x"514235",x"504134",x"483b2e",x"483a2c",x"493b2d",x"4d3e31",x"514336",x"57473b",x"615143",x"635244",x"251c14",x"251d15",x"261d15",x"261c14",x"251c14",x"231b13",x"231b13",x"231b12",x"20160d",x"191109",x"1d140b",x"20160c",x"20160c",x"291d11",x"281b10",x"271b0f",x"23180d",x"281b10",x"2d1f13",x"281c10",x"2d1f13",x"322316",x"322416",x"312215",x"332416",x"332416",x"382819",x"3b291a",x"39281a",x"3a291a",x"382718",x"3b291a",x"3c2a1a",x"3a2919",x"402e1d",x"3d2c1d",x"3b291a",x"3d2b1b",x"3f2c1c",x"3e2c1d",x"3f2c1c",x"422f1f",x"3e2b1b",x"412e1d",x"44311f",x"473221",x"412d1d",x"3c2b1b",x"3b291a",x"412f1f",x"423020",x"433121",x"453222",x"463424",x"473524",x"473423",x"58402c",x"1d160f",x"1f160d",x"21160d",x"21160d",x"1e140b",x"1d140b",x"22170d",x"251a0f",x"23180d",x"23180e",x"2d2014",x"25190f",x"281b10",x"291c11",x"2a1d12",x"261a0f",x"2b1e12",x"2c1e12",x"281c10",x"251a0f",x"2f2114",x"2c1e12",x"2c1f12",x"271a0f",x"2f2114",x"2d1f13",x"342416",x"312215",x"2f2114",x"312215",x"322315",x"322315",x"352517",x"352517",x"322316",x"39281a",x"352517",x"372718",x"352517",x"392819",x"392819",x"392819",x"3a2a1b",x"372618",x"332416",x"3c2a1b",x"3b2a1b",x"3a281a",x"39281a",x"372718",x"3b2a1a",x"4a3623",x"59402a",x"150e07",x"302214",x"2d1f12",x"312214",x"382719",x"382718",x"150e07",x"150e07",x"150e07",x"20160c",x"20160c",x"22170d",x"22170d",x"291c11",x"261a0f",x"23180e",x"22170d",x"20150c",x"23180e",x"281c10",x"251a0f",x"2b1e13",x"23180d",x"281b10",x"291c11",x"24190f",x"23180e",x"23180e",x"22170d",x"251a0f",x"25190f",x"2b1e12",x"281c10",x"21170d",x"1f150b",x"261a0f",x"24190e",x"2c1f12",x"291c11",x"2d2013",x"2c1f12",x"20160c",x"2a1d11",x"22170d",x"281b10",x"261a0f",x"2b1e12",x"291c11",x"281b10",x"24190e",x"2b1e12",x"23180d",x"23180e",x"271c11",x"23180d",x"22170d",x"2b1d12",x"24190f",x"291d11",x"291c11",x"25190e",x"2a1d11",x"25190f",x"291d11",x"23180d",x"21170d",x"24180e",x"23180e",x"20160c",x"25190f",x"23180e",x"23180e",x"23180d",x"23180d",x"22170d",x"24190e",x"24190e",x"21160d",x"23180e",x"23180e",x"20160c",x"22170d",x"23180d",x"23180d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e1c10",x"2e1c10",x"372112",x"2f1b0f",x"362011",x"3a2210",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"27160a",x"24150a",x"311c0d",x"341d0d",x"361f0e",x"371f0e",x"311b0c",x"311b0b",x"2e180a",x"2d170a",x"2d190a",x"351d0c",x"331c0c",x"371f0d",x"3a210f",x"3b210f",x"39200e",x"3c220f",x"2c190b",x"341c0c",x"371f0e",x"3b210f",x"39200f",x"361e0d",x"351d0d",x"381f0e",x"38200e",x"311a0b",x"351e0d",x"39200f",x"3b210f",x"361e0d",x"361e0d",x"3a200e",x"341c0c",x"321c0c",x"351d0d",x"331c0c",x"2c170a",x"341d0c",x"351d0d",x"341c0c",x"361d0d",x"321b0b",x"341c0c",x"361e0d",x"361e0d",x"371f0d",x"321b0c",x"301a0b",x"311a0b",x"2f1a0b",x"301a0b",x"311b0b",x"311a0b",x"2c180a",x"2d190b",x"150e07",x"1f1208",x"251509",x"231409",x"221409",x"1f1208",x"1f1208",x"492a13",x"492a13",x"3e2411",x"321c0d",x"2e1b0c",x"3c230f",x"3f2311",x"3c2210",x"3b220f",x"39210f",x"25150a",x"26160a",x"331d0d",x"231c15",x"201912",x"1d1710",x"26180c",x"28170a",x"25160a",x"351e0e",x"331c0c",x"2f1b0c",x"321c0c",x"2e1a0b",x"351d0d",x"351e0e",x"351d0d",x"371f0d",x"351d0d",x"351d0d",x"39200e",x"38200e",x"331d0d",x"371f0e",x"381f0e",x"341d0d",x"341d0d",x"371f0e",x"38200f",x"371f0e",x"361f0e",x"381f0e",x"38200e",x"341d0d",x"341d0d",x"351d0d",x"2b180a",x"2d170a",x"2b170a",x"301a0b",x"321c0c",x"351d0d",x"3a210f",x"39200e",x"371f0e",x"351e0e",x"381f0e",x"351d0d",x"351d0d",x"381f0e",x"38200e",x"3a210f",x"371f0e",x"39200e",x"3a210f",x"351d0d",x"321c0c",x"3a210f",x"39200f",x"381f0e",x"311b0c",x"341d0d",x"341d0d",x"351d0d",x"18110a",x"28180c",x"29190f",x"2d1c11",x"291b11",x"241910",x"4b2a13",x"3b2310",x"402612",x"3d2410",x"3e2310",x"432813",x"3a210f",x"3b2310",x"37200f",x"3b2210",x"351e0e",x"170f07",x"23150a",x"27170b",x"402817",x"3b3027",x"191008",x"1d1108",x"22150b",x"432e21",x"2e251e",x"51483e",x"51483e",x"000000",x"000000",x"000000",x"000000"),
(x"886d54",x"886c55",x"574b3f",x"504338",x"493d33",x"4b3d30",x"43372c",x"41352a",x"45372b",x"42352a",x"46382c",x"44372b",x"493b2e",x"493b2e",x"4f3f31",x"4e3e2f",x"513f2f",x"4d3c2e",x"4f3d2d",x"513f2f",x"4e3c2d",x"554131",x"574333",x"574435",x"584434",x"554333",x"584535",x"524130",x"564433",x"554130",x"513e2e",x"513d2b",x"56412f",x"54402f",x"543f2d",x"503d2c",x"54412f",x"55412f",x"564230",x"594532",x"4e3e2e",x"544130",x"564232",x"564332",x"584534",x"594633",x"5b4735",x"5a4533",x"5b4534",x"594433",x"5b4735",x"5a4635",x"5b4837",x"5c4837",x"5d4a39",x"5c4837",x"604b38",x"5a4736",x"5e4a37",x"594635",x"5a4736",x"584635",x"574637",x"584738",x"544537",x"584737",x"523f31",x"4e3e30",x"4e3e30",x"4c3c2f",x"504132",x"4f3f31",x"4f3f33",x"504133",x"514032",x"4f3f31",x"4e3e30",x"4c3c2e",x"4e3e31",x"4b3c2f",x"524133",x"57483b",x"625142",x"615142",x"261d15",x"271e16",x"271d15",x"241b12",x"241a12",x"231a11",x"231911",x"20180f",x"1e150b",x"1e140b",x"1d140b",x"1d140b",x"23180e",x"251a0f",x"25190e",x"281b0f",x"2a1d11",x"281b10",x"2a1d11",x"2c1e12",x"2d1f13",x"312215",x"342416",x"332416",x"3a2a1a",x"3b2a1b",x"3b2a1b",x"3c2a1b",x"3a291a",x"3e2c1c",x"3d2b1c",x"3f2d1d",x"3f2d1d",x"412f1f",x"412f1f",x"43301f",x"3f2d1c",x"3d2b1c",x"412e1e",x"402e1d",x"44311f",x"43301f",x"432f1e",x"432f1f",x"43301f",x"43301f",x"3a2819",x"3b2818",x"402e1d",x"43301f",x"42301f",x"463321",x"463321",x"453322",x"463324",x"463423",x"634b34",x"1d160f",x"211910",x"1e140b",x"1e140b",x"1e140b",x"1e140b",x"21170d",x"271b10",x"271b10",x"2b1e12",x"261a0f",x"291c11",x"2a1d11",x"291c11",x"291c11",x"2a1d11",x"2f2114",x"2c1e12",x"2b1e12",x"2d1f13",x"312215",x"2b1d11",x"2e1f12",x"2c1f12",x"322315",x"2e2013",x"2d1f13",x"2d1f13",x"322416",x"362617",x"372719",x"352618",x"3a291a",x"39291a",x"3a291a",x"3a291a",x"3c2b1b",x"3a291a",x"3a291a",x"372819",x"3c2b1b",x"3c2b1c",x"3d2b1b",x"3a291a",x"3b2a1b",x"39281a",x"3a291a",x"3a291a",x"3f2d1d",x"3c2a1b",x"39281a",x"4b3724",x"58402b",x"181008",x"312214",x"322315",x"362517",x"342416",x"392819",x"150e07",x"150e07",x"150e07",x"1e140b",x"24190f",x"22170d",x"271b10",x"23180e",x"251a0f",x"261a0f",x"24180e",x"261a10",x"271b10",x"22170d",x"2b1e12",x"261a0f",x"23180e",x"261a10",x"261a0f",x"2b1e12",x"261a0f",x"251a0f",x"2a1d11",x"281b10",x"291c11",x"251a0f",x"23170d",x"25190e",x"291c11",x"281b10",x"281c10",x"271b10",x"2b1e12",x"281c10",x"2c1e12",x"291d11",x"2a1e12",x"2d2013",x"2c1f13",x"291c11",x"2b1e12",x"2d2013",x"2a1d11",x"302215",x"271b10",x"2d2013",x"24190f",x"291d11",x"2d1f13",x"2a1d11",x"261a0f",x"261a0f",x"2a1d11",x"251a0f",x"23170d",x"281b10",x"291d11",x"2c1f13",x"22160c",x"22170d",x"271b10",x"25190e",x"23180e",x"271b10",x"24190e",x"20160c",x"22170d",x"21160d",x"24190f",x"22170d",x"271b10",x"251a0f",x"20160c",x"261a0f",x"24180e",x"24190e",x"24190f",x"24190f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e1d11",x"2e1d11",x"331f11",x"311d0f",x"382111",x"3c2311",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"23150a",x"27170b",x"361f0e",x"321c0d",x"2e1a0b",x"3b220f",x"351e0d",x"351e0d",x"371e0e",x"3a200e",x"351d0d",x"351d0d",x"331d0c",x"3a200e",x"3a200e",x"3d220f",x"3a200e",x"381f0e",x"381f0e",x"3b210f",x"39200e",x"3a210f",x"39200f",x"3a210f",x"361f0e",x"341d0c",x"321c0c",x"351d0d",x"371f0d",x"3a200f",x"3a200e",x"351d0d",x"39200e",x"39200f",x"3a200e",x"391f0e",x"351e0d",x"321c0c",x"331c0c",x"301a0b",x"341d0c",x"351d0c",x"3c210e",x"391f0e",x"391f0e",x"331b0b",x"321b0c",x"381f0e",x"361e0d",x"361e0d",x"321b0b",x"331b0b",x"2e190a",x"311b0b",x"321b0b",x"311a0b",x"2a170a",x"150e07",x"1d1108",x"251509",x"211309",x"201208",x"1c1108",x"1c1108",x"492b14",x"492b14",x"3e2512",x"2d1a0b",x"25150a",x"3c220f",x"3a210f",x"38200f",x"3b220f",x"371f0e",x"25150a",x"29180b",x"301c0c",x"231c15",x"1f1912",x"1f150f",x"2a190d",x"211409",x"211409",x"2c190b",x"321c0c",x"331c0c",x"321c0c",x"301a0b",x"341d0d",x"321c0c",x"381f0e",x"39200e",x"371f0e",x"38200f",x"3a210f",x"361f0f",x"3b2210",x"3a2210",x"3c2310",x"402512",x"3c2311",x"3c2311",x"3f2411",x"3f2411",x"3b2210",x"39210f",x"3b210f",x"38200e",x"3a210f",x"39200f",x"381f0e",x"311c0c",x"351d0d",x"311c0c",x"381f0d",x"351d0d",x"371f0d",x"371f0e",x"371f0e",x"361e0d",x"361e0d",x"381f0e",x"39200e",x"3d2310",x"3b220f",x"3c220f",x"3a210f",x"361e0d",x"331c0c",x"351d0c",x"361e0d",x"361e0d",x"361e0d",x"341d0c",x"351d0d",x"361f0e",x"371f0e",x"371e0d",x"18110a",x"24160b",x"29190f",x"2e1d11",x"2c1c11",x"271a11",x"4a2a13",x"3d2411",x"3f2512",x"3d2311",x"402511",x"452914",x"3d2310",x"38200f",x"3a2210",x"3d2411",x"361f0e",x"180f08",x"23150a",x"28180b",x"3f2817",x"3c332c",x"190f08",x"1d1208",x"26170c",x"462f22",x"27211a",x"4e453b",x"4e453b",x"000000",x"000000",x"000000",x"000000"),
(x"8c7058",x"8a6d55",x"5b4e42",x"514438",x"4e4236",x"493d31",x"44362b",x"45372a",x"423529",x"43362a",x"45372a",x"49392c",x"47382b",x"493a2c",x"4e3d2e",x"514030",x"4f3f31",x"503f2f",x"4c3c2d",x"513f30",x"564535",x"594434",x"5a4635",x"564534",x"594636",x"594738",x"584636",x"584534",x"564231",x"4e3c29",x"4e3c2c",x"523d2c",x"584230",x"594330",x"5c4531",x"59432f",x"59432f",x"55412f",x"584331",x"57412e",x"53402f",x"5a4533",x"5a4533",x"5b4633",x"5b4634",x"5f4a36",x"5c4735",x"5f4a38",x"5b4836",x"574332",x"5c4835",x"584533",x"5d4736",x"5d4734",x"5e4734",x"604a35",x"554434",x"574432",x"614b38",x"5d4936",x"594535",x"584533",x"544230",x"554435",x"594737",x"544536",x"574535",x"564434",x"4f3e31",x"534133",x"4d3e31",x"514031",x"4b3c2f",x"504133",x"554433",x"534234",x"514030",x"514031",x"4d3b2d",x"4b3c2e",x"4d3f32",x"5a4a3b",x"615040",x"625142",x"231b13",x"251c13",x"251c14",x"251c13",x"231911",x"231a11",x"221910",x"20160d",x"1e140b",x"1d130a",x"21170c",x"22170d",x"23180e",x"21160d",x"23180e",x"291c10",x"2d2013",x"281c10",x"2c1e12",x"2f2114",x"2d1f12",x"302215",x"362718",x"372719",x"382719",x"39291a",x"3c2b1c",x"3a291a",x"3d2c1d",x"402e1e",x"463323",x"402f1f",x"443221",x"412f1f",x"493523",x"423120",x"433120",x"453221",x"443121",x"412e1e",x"422f1e",x"3f2c1b",x"3e2b1b",x"402d1d",x"43301f",x"493522",x"4a3522",x"43301e",x"43301f",x"473321",x"422f1e",x"402e1d",x"432f1f",x"473423",x"4b3726",x"4b3725",x"5c432e",x"1c160f",x"22180f",x"21170d",x"21170d",x"22180e",x"22180e",x"22180e",x"261b10",x"2b1e12",x"281c11",x"281c11",x"271c11",x"271c11",x"2b1e13",x"2b1e12",x"251a0f",x"24180e",x"281c10",x"2b1e11",x"2f2114",x"342517",x"2f2114",x"312215",x"362618",x"322315",x"312214",x"2c1e12",x"302114",x"362718",x"3a2a1a",x"352517",x"382719",x"352618",x"3a2a1b",x"3b2a1b",x"362719",x"423020",x"3f2e1e",x"402f1f",x"3a2a1b",x"433020",x"423120",x"3d2c1d",x"3f2e1e",x"3f2d1e",x"3c2b1c",x"3c2a1b",x"3d2b1b",x"382718",x"382718",x"392819",x"523c28",x"59412c",x"191109",x"3a291a",x"3a281a",x"392819",x"362617",x"362617",x"150e07",x"150e07",x"150e07",x"23180e",x"23180e",x"21170d",x"2b1e13",x"271b10",x"261b10",x"281c11",x"281c11",x"2c1f13",x"2f2115",x"2d2014",x"2c1f13",x"2b1f13",x"2b1e13",x"2d2014",x"2f2115",x"261a0f",x"2d1f12",x"271b0f",x"271a0f",x"271b10",x"2d2013",x"2a1d11",x"2d2013",x"2f2114",x"2b1e12",x"2e2013",x"312214",x"2a1d11",x"281b10",x"2a1d12",x"2e2014",x"2e2114",x"2d2013",x"2c1f13",x"2b1e13",x"2d1f13",x"2e2114",x"302215",x"2e2114",x"322417",x"312316",x"2f2115",x"2c1f13",x"302216",x"2f2115",x"2f2115",x"2b1e13",x"291c11",x"2d1f12",x"2b1d11",x"271a0f",x"2b1e11",x"2b1e12",x"2e2013",x"2b1e12",x"2d1f13",x"291d11",x"25190e",x"25190e",x"261a0f",x"24190e",x"24190f",x"24190e",x"251a0f",x"261a0f",x"24190f",x"271c11",x"24190f",x"2a1d12",x"251a0f",x"251a0f",x"251a0f",x"281c11",x"281c11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1c11",x"2d1c11",x"311d11",x"362011",x"331e10",x"341d0e",x"150e07",x"150e07",x"150e07",x"1a1008",x"1d1108",x"231409",x"1e1208",x"2a170a",x"2f1a0b",x"341d0d",x"341d0d",x"321c0c",x"301b0b",x"321b0c",x"341d0c",x"351d0d",x"321c0d",x"361e0d",x"341c0c",x"361e0d",x"39200e",x"351d0d",x"3a200e",x"3a200e",x"351e0d",x"341d0d",x"3b210f",x"381f0e",x"371f0e",x"341d0c",x"321c0c",x"351d0d",x"381f0e",x"38200e",x"3c210f",x"3b200e",x"371f0e",x"381f0d",x"371e0d",x"341c0c",x"351d0d",x"351d0d",x"351e0d",x"381f0e",x"371f0e",x"38200e",x"39200f",x"341c0c",x"361e0d",x"381f0e",x"3f2411",x"3d2310",x"3a210f",x"361e0d",x"321b0b",x"321b0b",x"321b0b",x"351d0d",x"391f0d",x"371e0d",x"371f0e",x"331c0d",x"150e07",x"1f1208",x"2e190b",x"2c180b",x"29190c",x"21140a",x"21140a",x"462814",x"462814",x"3c2311",x"2e1a0b",x"2a180b",x"3a210f",x"3c2210",x"321c0d",x"371f0e",x"39200f",x"27160a",x"28170a",x"321d0d",x"221b15",x"201912",x"1d140d",x"26160a",x"2a180b",x"26160a",x"321c0c",x"2f1a0b",x"331c0c",x"2f1a0b",x"321c0c",x"331c0c",x"331d0d",x"351e0d",x"341e0d",x"39200f",x"371f0e",x"381f0e",x"341d0d",x"381f0e",x"361f0e",x"341d0d",x"361f0e",x"331c0d",x"321c0c",x"381f0e",x"361e0d",x"331c0c",x"301b0c",x"341d0d",x"361e0d",x"361e0d",x"351d0d",x"351d0c",x"351d0d",x"361e0d",x"321c0c",x"351e0d",x"341d0c",x"341c0c",x"381f0d",x"361e0d",x"351d0d",x"371f0e",x"3a200e",x"351d0d",x"381f0e",x"381f0e",x"361e0d",x"361e0d",x"341d0d",x"361e0d",x"361e0d",x"38200e",x"39200e",x"38200e",x"361e0d",x"351d0d",x"331c0c",x"331c0c",x"361e0d",x"170f07",x"25170c",x"301e11",x"322013",x"2f1e12",x"281b11",x"492913",x"3d2411",x"3d2310",x"3b2310",x"351e0d",x"3d2310",x"3f2411",x"3d2311",x"38200f",x"3c2311",x"3a210f",x"150e07",x"24150a",x"2a190b",x"3a200f",x"383028",x"190f08",x"1d1208",x"23160b",x"38291f",x"2b241d",x"4b4339",x"4b4339",x"000000",x"000000",x"000000",x"000000"),
(x"856951",x"8e7158",x"5e5144",x"55483b",x"4c3f33",x"483b2f",x"413428",x"413429",x"43362a",x"45372b",x"44372b",x"44362a",x"443529",x"47392b",x"4f3d2d",x"4b3b2d",x"4d3c2f",x"503f2f",x"514030",x"4e3e2e",x"513f2f",x"544030",x"534030",x"534131",x"574433",x"574434",x"594636",x"554333",x"564333",x"564130",x"54402f",x"564231",x"5a4531",x"574330",x"56412f",x"5a4430",x"54402d",x"5a4330",x"5d4530",x"57412d",x"543f2d",x"513e2d",x"54412f",x"554131",x"574331",x"5c4735",x"584433",x"594433",x"5e4835",x"594432",x"554131",x"574331",x"564332",x"57422f",x"5c4531",x"5a4431",x"584331",x"574230",x"584532",x"5a4533",x"574331",x"5b4533",x"544233",x"584331",x"564334",x"5b4938",x"564536",x"544333",x"4e3d2f",x"544133",x"503f31",x"4e4134",x"4c3d30",x"4f3e2f",x"554333",x"534130",x"4c3c2e",x"493a2d",x"48382b",x"4c3c2d",x"514032",x"554436",x"5a493a",x"5d4c3c",x"201810",x"221a11",x"1f1710",x"211910",x"21180f",x"21180f",x"1f160d",x"1d130a",x"1d140b",x"1e140b",x"20160c",x"23180e",x"23180d",x"2e2013",x"25190f",x"281c10",x"281c10",x"291c11",x"2b1e11",x"2b1d11",x"2b1d11",x"312215",x"322316",x"332316",x"3a291a",x"38281a",x"382718",x"382718",x"3d2b1b",x"3f2c1c",x"3b2a1a",x"3d2b1b",x"422f1f",x"3e2c1c",x"3e2b1c",x"402d1d",x"453120",x"422f1e",x"422f1e",x"422e1d",x"3f2c1c",x"3e2c1c",x"45311f",x"43301f",x"432f1e",x"463320",x"432f1e",x"45311f",x"3e2b1b",x"44301f",x"44301f",x"402d1c",x"422e1d",x"433020",x"463323",x"443222",x"5c432e",x"1d1610",x"231910",x"20160c",x"20160c",x"21160d",x"20150c",x"22170d",x"291c11",x"25190f",x"281c10",x"23180e",x"291d11",x"251a0f",x"2c1f12",x"291c10",x"2a1d11",x"291c11",x"2b1e11",x"291c11",x"2e2013",x"342517",x"302114",x"322316",x"312214",x"312215",x"312215",x"2f2013",x"2f2013",x"312215",x"362617",x"362618",x"392819",x"3a291a",x"382718",x"3a2819",x"382818",x"3b2a1a",x"392819",x"382718",x"3f2d1d",x"3b291a",x"382718",x"3e2c1c",x"362618",x"382818",x"3d2b1c",x"372617",x"3f2d1c",x"3e2c1c",x"3c2a1a",x"3d2b1c",x"493522",x"543f29",x"191109",x"382818",x"342416",x"372718",x"372718",x"342416",x"150e07",x"150e07",x"150e07",x"24190e",x"20160c",x"23180e",x"23180d",x"20160c",x"291c10",x"23180e",x"22170d",x"271b10",x"251a0f",x"2a1d11",x"2a1d11",x"2b1e12",x"2b1e12",x"2d1f12",x"2a1d11",x"291c10",x"2a1d11",x"2b1e12",x"2b1e11",x"2b1d12",x"2e2013",x"2d2013",x"2c1e12",x"312215",x"291c11",x"271b10",x"2b1e12",x"2b1e11",x"2b1d11",x"2d1f13",x"271b10",x"2d1f13",x"2c1e12",x"2d1f13",x"2c1e12",x"2c1e12",x"2d1f12",x"2b1e12",x"291d11",x"291d11",x"2d1f13",x"2a1d11",x"2e2013",x"2f2114",x"2f2114",x"2e2013",x"2e2013",x"2b1d11",x"2a1d11",x"2d1f13",x"2d1f13",x"291c11",x"2b1d11",x"2f2114",x"291d11",x"2c1f12",x"281b10",x"291c11",x"24190e",x"23180d",x"261a0f",x"271b10",x"20150c",x"22170d",x"25190f",x"251a0f",x"25190e",x"281c10",x"23180e",x"23180e",x"24190e",x"22170d",x"281c10",x"281c10",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c1c10",x"2c1c10",x"2e1c10",x"331f12",x"311d0f",x"3b2310",x"160e07",x"160e07",x"150e07",x"150e07",x"221409",x"201208",x"201308",x"2c190b",x"311c0c",x"341d0d",x"361e0d",x"351d0d",x"351e0d",x"331c0c",x"301b0c",x"331c0c",x"351d0d",x"39200e",x"38200e",x"38200e",x"381f0e",x"371f0e",x"371e0d",x"331c0c",x"331c0c",x"341d0c",x"341d0c",x"371f0d",x"381f0e",x"351e0d",x"331d0d",x"321c0c",x"361d0d",x"3c220f",x"3f2411",x"3f2411",x"3c210f",x"39200e",x"3f2411",x"3c2210",x"381f0e",x"361d0d",x"3c2210",x"3d220f",x"361e0d",x"38200e",x"371e0e",x"3c220f",x"3a210f",x"381f0e",x"351d0d",x"381f0e",x"341d0c",x"39200e",x"3c220f",x"3b210e",x"3c210f",x"311a0b",x"341c0c",x"301a0b",x"2f1a0b",x"2e1a0b",x"150e07",x"1e1208",x"2d1a0d",x"2d1a0d",x"27170c",x"22150b",x"22150b",x"4a2a15",x"4a2a15",x"3b2210",x"2e1a0b",x"29180b",x"39200f",x"38200f",x"39210f",x"38200e",x"38200f",x"28170a",x"2a180b",x"321d0e",x"221b14",x"1f1812",x"1b140c",x"231409",x"26160a",x"241509",x"301b0b",x"2d190b",x"2e190b",x"2e190b",x"2f1a0b",x"311b0c",x"311c0c",x"341d0d",x"361f0d",x"38200f",x"39200f",x"3a210f",x"39200f",x"351e0d",x"331c0d",x"331d0d",x"301a0b",x"311c0c",x"371f0e",x"381f0e",x"351d0d",x"341d0d",x"311c0c",x"331d0d",x"2d190b",x"351e0d",x"371f0d",x"361e0d",x"341c0c",x"371f0d",x"351d0d",x"341d0d",x"381f0e",x"38200f",x"381f0e",x"351e0d",x"371f0d",x"311b0c",x"331c0c",x"311b0b",x"341d0c",x"371f0d",x"3a200e",x"371f0e",x"351e0d",x"39200e",x"331c0c",x"351e0d",x"3a210f",x"3a2210",x"39200e",x"351d0d",x"39200f",x"3c2311",x"3a210f",x"170f07",x"28180c",x"311e10",x"311f13",x"2f1e13",x"281b11",x"4a2a14",x"3d2310",x"3e2411",x"3a200f",x"381f0e",x"3c2311",x"3e2411",x"402612",x"361f0e",x"3d2411",x"39200f",x"180f07",x"24150a",x"211309",x"443024",x"2b241c",x"191008",x"1d1208",x"1f1309",x"2c2017",x"302821",x"4d443b",x"4d443b",x"000000",x"000000",x"000000",x"000000"),
(x"846954",x"816751",x"5e5044",x"54473a",x"504235",x"4d3f33",x"493c30",x"46392d",x"45372b",x"493a2d",x"46382b",x"44362a",x"493829",x"48392b",x"513f2e",x"4f3e2f",x"513f30",x"513f30",x"554232",x"564434",x"564333",x"554333",x"534130",x"544232",x"5a4837",x"5b4838",x"594736",x"5a4736",x"584535",x"574332",x"574331",x"55412f",x"584330",x"594332",x"57422f",x"594330",x"58422e",x"5c4531",x"5d4732",x"5b4431",x"5a432f",x"59432e",x"5b4430",x"584432",x"5f4835",x"5b4533",x"5e4834",x"594433",x"5c4736",x"594534",x"594432",x"594331",x"57412f",x"5a4432",x"59432f",x"5c4632",x"574534",x"5b4633",x"594330",x"5a4531",x"584331",x"574331",x"564331",x"54402f",x"5a4634",x"584636",x"594838",x"574535",x"554335",x"4f4033",x"554536",x"554537",x"4f3f32",x"4f3f32",x"534335",x"4d3d2f",x"4e3e30",x"4c3c2d",x"4b3b2d",x"493b2e",x"4f3f32",x"4d3f31",x"5c4a3c",x"5c4b3c",x"20170f",x"21180f",x"20180f",x"211810",x"20170e",x"20170d",x"20160c",x"1d140b",x"1d140b",x"1d130b",x"1c130a",x"1f150b",x"20150c",x"2a1d12",x"261a10",x"261a0f",x"2a1d11",x"2f2114",x"332416",x"322316",x"322316",x"312215",x"3a291a",x"3a291a",x"3e2c1c",x"3a291a",x"382718",x"3a291a",x"3f2c1c",x"3c2a1b",x"3b291a",x"402d1d",x"3f2c1c",x"3e2c1c",x"422f1f",x"42301f",x"433020",x"443120",x"483322",x"432f1e",x"422f1e",x"43301f",x"402d1c",x"422f1e",x"422f1e",x"43301f",x"4a3623",x"483422",x"4a3623",x"473221",x"473321",x"44311f",x"422e1e",x"4a3625",x"473523",x"463423",x"5f4630",x"1d1710",x"231910",x"20160c",x"1d140b",x"20160c",x"20150c",x"251a0f",x"23180d",x"291c11",x"24190f",x"261b10",x"271b10",x"2c1f13",x"291c11",x"2a1d11",x"291d11",x"2c1f12",x"281b10",x"291d11",x"2a1d11",x"2e2114",x"302215",x"322316",x"302215",x"382719",x"392819",x"382719",x"352517",x"322416",x"382819",x"372718",x"3c2b1b",x"372718",x"3e2b1c",x"3a291a",x"3a291a",x"372718",x"392819",x"3b2a1b",x"3b291a",x"402e1e",x"3d2b1c",x"3a2a1b",x"3e2d1d",x"3d2c1c",x"3e2c1c",x"3d2b1b",x"352517",x"372618",x"382819",x"3a291a",x"4f3a26",x"4d3925",x"191109",x"382719",x"3b2a1b",x"39281a",x"3b2a1b",x"3b2a1a",x"150e07",x"150e07",x"150e07",x"251a0f",x"261a0f",x"23180e",x"281c10",x"20160c",x"291c11",x"22170d",x"24190e",x"23180e",x"2e2013",x"251a0f",x"281c10",x"2e2114",x"2d1f13",x"2e2014",x"2d1f13",x"2c1e12",x"271b10",x"2a1d11",x"291d11",x"2a1d11",x"2e1f13",x"2e2114",x"322416",x"2f2114",x"2f2214",x"322316",x"322416",x"2f2114",x"302114",x"2e2013",x"302215",x"2d1f13",x"2d2013",x"332416",x"2e2013",x"2c1f13",x"2e2014",x"302114",x"2d1f13",x"2f2114",x"2e2013",x"2d1f13",x"2e2013",x"2a1d12",x"312216",x"332416",x"312215",x"2c1e12",x"312215",x"322315",x"2b1e12",x"2c1e12",x"2e1f13",x"2d1f13",x"302215",x"2d2013",x"2b1f12",x"2f2114",x"2b1e12",x"261a0f",x"281b10",x"281c10",x"2a1d11",x"251a0f",x"23180e",x"2b1e12",x"2a1d11",x"2a1d12",x"291c11",x"271b10",x"271b10",x"2b1e12",x"261a0f",x"261a0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b1b10",x"2b1b10",x"2c1c11",x"301d0f",x"311d0f",x"2d190c",x"180f07",x"180f07",x"170f07",x"160e07",x"1e1209",x"24150a",x"221409",x"331d0d",x"371f0e",x"3a200f",x"361e0d",x"381f0e",x"341c0c",x"351d0c",x"341d0c",x"331c0c",x"361e0d",x"381f0d",x"361e0d",x"2b180b",x"371f0e",x"381f0e",x"39200e",x"39200e",x"361e0d",x"341d0d",x"391f0e",x"381f0e",x"3d2310",x"3c2310",x"3a2210",x"3b2210",x"3b2210",x"3a210f",x"3c2210",x"3c2210",x"3c2310",x"3e2410",x"3c2210",x"341d0c",x"351d0d",x"39200e",x"3e2310",x"3a200e",x"3e2310",x"3c220f",x"3a200e",x"3d220f",x"39200e",x"2f1a0b",x"3b210e",x"3a200d",x"3a1f0d",x"391f0d",x"341d0c",x"301b0b",x"361f0d",x"38200e",x"361f0e",x"351e0d",x"331d0d",x"361e0d",x"150e07",x"23160b",x"28180c",x"2d1a0d",x"2a1a0c",x"22150b",x"22150b",x"412512",x"412512",x"3d2411",x"2e1a0c",x"2e1a0c",x"351e0e",x"3c2310",x"3e2411",x"3c2310",x"331d0d",x"27160a",x"2d1a0c",x"301b0c",x"201913",x"1d1710",x"171009",x"201208",x"261509",x"28170b",x"351e0d",x"311c0d",x"311b0c",x"341d0d",x"38200f",x"38200e",x"39200e",x"351d0d",x"361e0d",x"361e0d",x"38200f",x"3d2311",x"3b2310",x"3d2411",x"3b2210",x"3a210f",x"361f0e",x"351e0d",x"3a210f",x"3a210f",x"361f0e",x"3d2310",x"3a220f",x"3b220f",x"361f0e",x"301b0c",x"341d0c",x"331c0c",x"381f0d",x"341d0c",x"331c0c",x"331d0c",x"301b0b",x"351d0d",x"3a200f",x"39200f",x"381f0e",x"39200e",x"371e0e",x"321c0c",x"371f0e",x"301b0c",x"371f0e",x"39210f",x"3d2310",x"38200f",x"3c2210",x"39210f",x"3a210f",x"39210f",x"3a210f",x"3c2310",x"3a220f",x"341d0d",x"331c0c",x"170f07",x"2b1a0d",x"311e10",x"311f12",x"2c1d11",x"271b11",x"472711",x"38200e",x"3f2411",x"381f0e",x"371f0e",x"442914",x"3a2210",x"3e2411",x"361e0d",x"412612",x"39210f",x"181008",x"231509",x"1f1208",x"422e21",x"332c24",x"190f08",x"1d1108",x"1f1209",x"281c14",x"3a332b",x"4a4138",x"4a4138",x"000000",x"000000",x"000000",x"000000"),
(x"8a6f56",x"8b6f57",x"5a4c3f",x"56473b",x"504236",x"4b3e32",x"4c3f32",x"45392e",x"45382d",x"47392c",x"483a2d",x"4b3b2d",x"49382a",x"4f3d2e",x"4e3f30",x"534030",x"584536",x"564434",x"5b4837",x"5a4737",x"5b4837",x"5a4635",x"5b4735",x"5c4937",x"614d3a",x"5f4b39",x"5d4a39",x"5b4737",x"5b4635",x"5b4736",x"594432",x"5a4534",x"5c4835",x"5c4836",x"5f4936",x"5c4633",x"5a4431",x"5f4732",x"5c4431",x"5a4330",x"5c442f",x"5d4530",x"54402f",x"5c4431",x"5a4430",x"594432",x"604934",x"624b37",x"604b38",x"604a37",x"5f4835",x"5d4634",x"5a4532",x"554130",x"5a4534",x"5c4734",x"644c37",x"5c4733",x"5d4834",x"614a37",x"5d4735",x"5e4631",x"584331",x"584330",x"5c4631",x"594736",x"594839",x"5c4a38",x"584636",x"554334",x"574637",x"544436",x"524234",x"514031",x"504032",x"4f3e2f",x"4b3a2b",x"503f30",x"4c3c2d",x"503f30",x"514134",x"564739",x"635041",x"635040",x"1f160e",x"1d150d",x"21170e",x"21170e",x"21180f",x"1f150c",x"1e150c",x"1f150c",x"1e140b",x"1e140b",x"1d140b",x"23180e",x"24190f",x"261a10",x"2d1f13",x"2d2014",x"2f2114",x"2e2014",x"2e2115",x"302114",x"312215",x"342517",x"39281a",x"3b2a1b",x"39281a",x"392819",x"3c2b1b",x"3c2a1b",x"3e2c1d",x"3f2d1d",x"422f1f",x"433120",x"463221",x"443120",x"493523",x"483423",x"4a3725",x"463322",x"483423",x"4c3825",x"463220",x"453120",x"43301f",x"473221",x"453221",x"473321",x"483422",x"4c3825",x"493422",x"4a3524",x"4b3725",x"44301f",x"473321",x"483523",x"493424",x"493624",x"5f4630",x"1a140d",x"23190f",x"21160d",x"21170d",x"21170d",x"24190e",x"21170d",x"24190f",x"24190e",x"2c1f13",x"2b1e13",x"2c2014",x"2d2014",x"271b10",x"2f2115",x"2e2013",x"2b1e12",x"2e2014",x"2f2114",x"2e2114",x"2e2014",x"352618",x"362719",x"342517",x"362719",x"352618",x"382718",x"342417",x"382819",x"382819",x"3a291a",x"3b2a1a",x"352517",x"412f1e",x"3c2b1b",x"3d2b1c",x"3f2d1d",x"412e1e",x"3e2d1d",x"3e2c1d",x"3c2a1b",x"473422",x"422f1f",x"413020",x"3d2b1c",x"42301f",x"3f2d1d",x"3f2d1d",x"3b2a1a",x"422f1e",x"3e2c1c",x"5b432e",x"4d3825",x"191109",x"3a2a1b",x"3a291a",x"3c2b1c",x"3c2b1c",x"3a2919",x"150e07",x"150e07",x"150e07",x"261a0f",x"23180e",x"2c1f13",x"261b10",x"261a0f",x"271b10",x"2a1d11",x"2a1d11",x"271b10",x"2a1d12",x"261b10",x"2e2114",x"2d2014",x"2c1f14",x"302215",x"2c1f13",x"2b1e12",x"2a1d11",x"2b1e12",x"2d1f13",x"2d2013",x"302215",x"302215",x"2e2114",x"312316",x"2f2114",x"332417",x"2e2115",x"312215",x"2e2013",x"2e2014",x"322316",x"342517",x"322316",x"352518",x"2e2014",x"342517",x"332417",x"332416",x"332316",x"332417",x"302215",x"332416",x"352618",x"302215",x"362719",x"302215",x"302215",x"2f2115",x"332416",x"342416",x"2b1d12",x"322316",x"332417",x"2e2014",x"302215",x"2d2014",x"2f2114",x"2c1f13",x"2a1d12",x"281c10",x"25190f",x"2b1d12",x"261a0f",x"291d11",x"291d11",x"2c1f13",x"24190e",x"2c1f12",x"2f2114",x"2a1d11",x"2a1d11",x"2a1d12",x"281c10",x"281c10",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291b10",x"291b10",x"2b1c10",x"2e1c0f",x"2f1d0f",x"2f1b0c",x"1a1008",x"1a1008",x"180f07",x"180f08",x"1c1108",x"150e07",x"241509",x"2c190b",x"2d190b",x"321c0c",x"311b0b",x"301b0b",x"2e190b",x"341c0c",x"301a0b",x"331c0c",x"381f0d",x"351d0d",x"39200d",x"381f0d",x"381f0e",x"3f2410",x"3c220f",x"361f0e",x"361e0d",x"351c0c",x"381f0e",x"3a210f",x"361f0e",x"39210f",x"38200e",x"3a210f",x"351d0d",x"351d0d",x"341d0d",x"331c0c",x"351d0d",x"341c0c",x"351c0c",x"301a0b",x"381f0d",x"39200e",x"3b210f",x"3c210f",x"39200e",x"3b210f",x"3a200e",x"39200e",x"331c0b",x"341c0b",x"381f0d",x"391f0d",x"3b200e",x"311b0b",x"381f0d",x"321b0b",x"371f0e",x"351d0d",x"38200e",x"38200e",x"351e0d",x"331d0d",x"17100a",x"26170c",x"29190e",x"2b1a0e",x"2c1b0f",x"24170d",x"24170d",x"422511",x"422511",x"392110",x"311c0d",x"2b190b",x"38200f",x"3b2210",x"3b2210",x"351e0e",x"361f0e",x"28170a",x"2c190b",x"301b0c",x"1f1811",x"1d1710",x"17110a",x"27170a",x"28180b",x"29180b",x"321c0c",x"311b0c",x"2f1a0b",x"2f1a0b",x"341e0e",x"36200f",x"38200f",x"39200e",x"381f0e",x"38200e",x"38200e",x"341d0d",x"361e0d",x"321c0c",x"39200e",x"351e0d",x"351e0d",x"311c0c",x"371f0e",x"331c0d",x"341c0d",x"351d0c",x"341c0c",x"331c0c",x"311b0b",x"301a0b",x"2e190b",x"331c0b",x"331c0c",x"331c0c",x"351d0c",x"361e0d",x"341d0d",x"2f1a0b",x"321c0c",x"311c0c",x"341e0d",x"3a210f",x"321c0c",x"2e180a",x"371e0d",x"39200f",x"3b220f",x"3a210f",x"39200f",x"38200f",x"361e0d",x"371e0d",x"2b180b",x"321c0c",x"331c0c",x"311b0b",x"2f190b",x"2f190b",x"311b0c",x"170f07",x"2a1a0c",x"311e11",x"332013",x"2e1d12",x"291d13",x"482812",x"39200e",x"3e2310",x"381f0e",x"3a200f",x"422713",x"3c2311",x"3d2411",x"331c0c",x"37200f",x"3d2310",x"191008",x"24150a",x"201208",x"422f23",x"3b332b",x"190f08",x"1d1108",x"1e1208",x"2a2018",x"413930",x"4a4037",x"4a4037",x"000000",x"000000",x"000000",x"000000"),
(x"7f6551",x"836752",x"584c40",x"57493c",x"534537",x"4a3d30",x"4a3c31",x"45382c",x"493a2d",x"4b3c2f",x"47392c",x"47382b",x"4c3c2d",x"4b3b2c",x"523f2f",x"503e2e",x"544332",x"5a4636",x"584635",x"584637",x"594735",x"594634",x"5c4938",x"5d4938",x"5c4838",x"594635",x"574535",x"574333",x"594735",x"564131",x"5a4634",x"5c4938",x"5e4a39",x"5a4736",x"5a4635",x"644d38",x"584330",x"5b442f",x"5b4430",x"5e4935",x"5e4632",x"5e4733",x"5e4733",x"5d4530",x"634c36",x"664b34",x"5d4836",x"614b36",x"5e4835",x"5f4a38",x"5f4936",x"5f4936",x"5c4633",x"5e4734",x"624b38",x"594532",x"594332",x"584331",x"55422f",x"564130",x"594431",x"57412f",x"55402e",x"513d2d",x"513f2e",x"56402f",x"534333",x"5b4737",x"5b4838",x"564434",x"554536",x"58483a",x"564537",x"564434",x"524231",x"4e3f31",x"4a3b2d",x"4b3a2c",x"4d3b2c",x"473829",x"4f3e2e",x"574739",x"5f4e3e",x"5e4e3e",x"22180f",x"21170e",x"1b130b",x"20170e",x"1d140b",x"1d140b",x"1d130b",x"1c130a",x"1c130a",x"1c130a",x"1e140b",x"20160c",x"261a0f",x"271a0f",x"2a1d11",x"302214",x"302215",x"2e2013",x"332417",x"3a291a",x"362618",x"3a291a",x"3a291a",x"402e1e",x"3d2c1c",x"3e2c1c",x"3f2c1c",x"3b2a1a",x"3e2b1b",x"422f1f",x"412f1f",x"422f1f",x"453221",x"453221",x"493523",x"473322",x"402d1d",x"412e1d",x"412e1d",x"3e2b1b",x"402d1c",x"3e2a1a",x"3f2b1b",x"3d2a19",x"422f1d",x"442e1d",x"3f2d1c",x"4a3623",x"4a3624",x"432f1e",x"473322",x"493523",x"473322",x"483424",x"473524",x"4a3726",x"634b33",x"1b150e",x"21180e",x"20150c",x"20160c",x"21160d",x"21170d",x"251a0f",x"251a0f",x"2b1e12",x"251a0f",x"271b10",x"2b1e11",x"271b10",x"271b10",x"281b10",x"291d11",x"271a0f",x"25190e",x"2a1d11",x"2a1d11",x"2d1e12",x"332416",x"342517",x"302215",x"382718",x"352518",x"3a291a",x"3b2a1b",x"3e2d1d",x"3a291a",x"362719",x"3b2b1b",x"3c2a1b",x"3a2919",x"382718",x"3e2b1b",x"3e2c1c",x"39291a",x"402e1e",x"352618",x"3d2c1c",x"443221",x"402e1e",x"3d2b1b",x"392819",x"3c2a1a",x"3b2919",x"3c2b1b",x"3a2818",x"3c2919",x"3b2919",x"533c27",x"442f1e",x"181008",x"3b2a1b",x"3c2b1c",x"3a2819",x"3a2a1b",x"3c2b1c",x"281c11",x"150e07",x"150e07",x"271b10",x"271b10",x"291c11",x"281b10",x"271b10",x"281c10",x"261a0f",x"2a1d12",x"2b1f13",x"2b1f13",x"2d1f13",x"312316",x"2c1f13",x"291c11",x"271b10",x"291c11",x"2b1e11",x"291d11",x"271a0f",x"2d1e12",x"2a1d11",x"2a1d11",x"2f1f13",x"281c10",x"302214",x"332417",x"312215",x"352618",x"332417",x"362719",x"312216",x"2f2115",x"352618",x"332517",x"332416",x"322315",x"302114",x"322315",x"352617",x"39291a",x"372719",x"322416",x"312216",x"312316",x"352618",x"2d1f12",x"2b1e12",x"312215",x"302214",x"2b1e11",x"2e1f12",x"2d1e12",x"2d1e12",x"281c10",x"2b1d11",x"2a1d11",x"342517",x"332417",x"2c1f12",x"2a1d12",x"2c1f13",x"2a1d12",x"2d1f13",x"271b10",x"2a1d12",x"2f2115",x"291c11",x"2c1e12",x"271b10",x"2a1d11",x"2d2013",x"2c1f13",x"2b1f13",x"291d11",x"291d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281a0f",x"281a0f",x"29190e",x"2f1c0f",x"2d1a0f",x"331d0d",x"1b1108",x"1b1108",x"190f08",x"160f07",x"1e1208",x"251509",x"1e1208",x"2b170a",x"2d180a",x"2f1a0b",x"341d0c",x"38200e",x"39200e",x"361e0d",x"341d0d",x"3a200e",x"3c220f",x"3c220f",x"3b210f",x"3a200e",x"321b0b",x"331c0c",x"351d0c",x"361e0d",x"3a200e",x"3c230f",x"38200f",x"3c220f",x"38200e",x"3b210f",x"361e0d",x"3a210f",x"3a210f",x"3a210f",x"39200e",x"39200f",x"3a210f",x"3b210f",x"39200e",x"381f0e",x"38200e",x"381f0e",x"371e0d",x"341d0c",x"351d0d",x"361d0d",x"39200e",x"381f0d",x"381f0d",x"391f0d",x"351d0c",x"331c0b",x"301a0a",x"321c0b",x"2e1a0a",x"311b0b",x"321b0c",x"331c0d",x"341d0d",x"341e0d",x"371f0e",x"381f0e",x"17110a",x"27190e",x"2e1c0f",x"2e1c0f",x"2a1a0f",x"24180f",x"24180f",x"462711",x"462711",x"3d2411",x"321d0d",x"28170b",x"38200f",x"3e2411",x"3b2210",x"311c0c",x"331c0c",x"2b190b",x"2b180b",x"2f1a0c",x"1d160f",x"1b150e",x"171009",x"1f1309",x"28170a",x"28170a",x"361e0d",x"351d0d",x"311c0c",x"2d190b",x"2c180a",x"311b0c",x"2d190b",x"2f1a0b",x"351d0d",x"3a210f",x"351e0d",x"361f0e",x"2a180b",x"301b0b",x"351d0d",x"361e0d",x"341c0c",x"301a0b",x"351d0c",x"361e0d",x"371e0d",x"341c0c",x"311b0b",x"311a0b",x"331c0c",x"331d0d",x"2f1b0c",x"381f0e",x"361e0d",x"371e0d",x"341d0d",x"381f0e",x"38200e",x"331c0c",x"321c0c",x"2e190b",x"321b0c",x"331c0c",x"371e0d",x"39200e",x"3c2310",x"381f0e",x"39200e",x"371f0e",x"331c0d",x"3b220f",x"3a210f",x"3a210f",x"361f0e",x"311c0d",x"3b2210",x"3a210f",x"371f0e",x"3a210f",x"371f0e",x"18110a",x"2c1a0d",x"2c1c11",x"2e1d11",x"312014",x"2b1c13",x"472812",x"381f0e",x"402512",x"3e220f",x"402512",x"3d2411",x"3d2311",x"3f2512",x"371f0d",x"3b2210",x"3a210f",x"181008",x"25160a",x"211309",x"534538",x"50473d",x"190f08",x"1d1108",x"1e1208",x"332b24",x"4d433a",x"4b4239",x"4b4239",x"000000",x"000000",x"000000",x"000000"),
(x"806751",x"806752",x"5a4d41",x"594b3e",x"504336",x"4e4034",x"493b2f",x"4a3b2e",x"493a2d",x"49392c",x"4e3e2d",x"4e3e2f",x"503f2e",x"4c3c2c",x"514032",x"53402f",x"564433",x"594534",x"5b4736",x"5d4735",x"574534",x"5e4935",x"5d4937",x"5e4b37",x"5c4836",x"594636",x"564332",x"594434",x"554231",x"544232",x"5e4836",x"614c39",x"624d3a",x"624d3b",x"614e3d",x"624b38",x"614936",x"5d4631",x"604733",x"5d4734",x"5e452f",x"5e4530",x"604832",x"5d4732",x"644c36",x"624a34",x"634b37",x"674e38",x"664e3a",x"664f3a",x"644d39",x"5f4937",x"664d38",x"5c4531",x"604936",x"5a4634",x"614933",x"5e4731",x"5d4733",x"5a4330",x"5c4531",x"55412f",x"554230",x"584331",x"56412f",x"5c4633",x"554231",x"594535",x"594635",x"564434",x"554535",x"584737",x"5a4737",x"5c4735",x"594735",x"534232",x"4d3d2d",x"4b3b2d",x"503f30",x"534132",x"574536",x"574739",x"614e3d",x"614f3f",x"1e150b",x"1f150c",x"1f150c",x"1f150c",x"1e140b",x"1d140b",x"1d140b",x"1e140b",x"1c130a",x"1c130a",x"20160c",x"261a0f",x"281c10",x"261a0f",x"2c1f12",x"2c1f13",x"2f2115",x"322316",x"302114",x"372719",x"3a291a",x"3c2b1c",x"3d2c1c",x"402f1f",x"433120",x"3f2d1d",x"3f2d1d",x"422f1f",x"3d2c1c",x"402e1e",x"443220",x"453221",x"473422",x"4a3624",x"4a3524",x"4b3724",x"4a3522",x"45311f",x"473220",x"3d2a19",x"412d1c",x"422f1c",x"473220",x"493422",x"432f1e",x"473320",x"473220",x"503b27",x"4d3825",x"463220",x"473321",x"4b3624",x"453221",x"473423",x"4c3827",x"4e3b29",x"694f37",x"1b150e",x"23190f",x"22180d",x"22170d",x"22180e",x"251a0f",x"24190f",x"251a0f",x"251a0f",x"2b1e12",x"281c11",x"291d11",x"25190f",x"2a1d11",x"271a0f",x"281b0f",x"23180d",x"2e2013",x"352517",x"322315",x"332416",x"342416",x"39291a",x"362719",x"3a281a",x"3d2b1c",x"3f2d1d",x"3a291a",x"3e2c1d",x"3f2d1e",x"402f1f",x"443221",x"402f1e",x"3c2a1b",x"453120",x"412f1e",x"402e1e",x"3d2c1c",x"3d2c1c",x"463322",x"423120",x"412f1f",x"443220",x"43301e",x"402d1c",x"3e2c1c",x"3c2919",x"3c2919",x"3e2b1a",x"3e2c1b",x"3d2b1c",x"573d29",x"503a26",x"191109",x"39291a",x"3a2a1b",x"362618",x"3b2a1a",x"3d2c1c",x"322416",x"150e07",x"150e07",x"291d12",x"281c11",x"251a0f",x"2d1f13",x"2d2014",x"271b10",x"2c1e13",x"2e2014",x"2a1e12",x"2c1f13",x"281c11",x"2f2115",x"322416",x"2b1e12",x"2e2013",x"2c1f12",x"291c10",x"281b0f",x"2d1f12",x"2a1d11",x"332416",x"2e1f13",x"2e2013",x"312215",x"312215",x"312316",x"342417",x"342416",x"312316",x"352618",x"362719",x"37281a",x"38291b",x"37281a",x"322416",x"342517",x"362719",x"342517",x"372719",x"372719",x"352618",x"37281a",x"352618",x"362619",x"352618",x"332416",x"332416",x"312215",x"302013",x"2d1f12",x"2b1d11",x"342416",x"332416",x"302114",x"2e2014",x"312215",x"312215",x"342517",x"2b1e12",x"2d2013",x"2b1e12",x"2b1e12",x"302215",x"2c1f13",x"312316",x"302316",x"302216",x"271b10",x"2f2115",x"2d2013",x"322416",x"2e2014",x"2d1f13",x"2d2014",x"2d2014",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281a0f",x"281a0f",x"29190e",x"2b1a0f",x"2b1a0e",x"2c190b",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"1b1108",x"211309",x"1b1008",x"29170a",x"2d190a",x"2e190b",x"301b0b",x"371f0e",x"361e0d",x"341d0d",x"38200e",x"402410",x"3a200f",x"39200e",x"351d0d",x"361e0d",x"38200e",x"3d2310",x"38200f",x"3d2410",x"3d2310",x"3a210f",x"381f0e",x"351d0d",x"361e0d",x"38200f",x"3c2310",x"3b210f",x"361f0e",x"331d0d",x"371e0d",x"351d0c",x"371e0d",x"3a210f",x"39200e",x"341d0c",x"361d0d",x"351d0c",x"3a200e",x"371f0e",x"341d0c",x"331c0c",x"371e0d",x"371f0d",x"341d0d",x"351d0c",x"391f0d",x"381f0d",x"391f0d",x"351d0c",x"2f1a0a",x"381f0d",x"301a0b",x"351e0d",x"351d0d",x"341c0c",x"331c0c",x"2c180a",x"19130c",x"23160d",x"2b1a0f",x"291a0f",x"281a10",x"24170f",x"24170f",x"462712",x"462712",x"3b2310",x"321d0d",x"201309",x"38200f",x"351e0d",x"311c0c",x"28160a",x"321c0c",x"2b190b",x"2b180b",x"311c0d",x"1b140d",x"19130c",x"171009",x"1e1108",x"221309",x"241409",x"2c180a",x"2c180a",x"2a1709",x"291509",x"211107",x"221107",x"211107",x"241208",x"2d180a",x"2d190a",x"2c180a",x"301b0b",x"321c0b",x"311b0c",x"301a0b",x"331c0c",x"361e0d",x"371f0d",x"361e0d",x"321b0c",x"331c0c",x"341c0c",x"321b0b",x"311b0b",x"2f1a0b",x"381f0e",x"311c0c",x"371f0e",x"371f0e",x"311b0c",x"3a210f",x"38200e",x"341d0d",x"2f1a0b",x"351e0d",x"39200e",x"3d2311",x"38210f",x"3d2310",x"3c2310",x"38200e",x"361e0d",x"351d0d",x"361f0e",x"3c2311",x"39200f",x"39200e",x"361e0d",x"351d0d",x"331c0c",x"341c0c",x"351e0d",x"341d0d",x"2f1a0b",x"331c0c",x"181009",x"28190d",x"301f13",x"301e12",x"2e1f15",x"271a11",x"462711",x"3a200f",x"361e0d",x"3b220f",x"422712",x"402512",x"3c2310",x"3f2411",x"351d0d",x"3c220f",x"3c220f",x"150e07",x"24150a",x"221409",x"544a3f",x"544b41",x"190f07",x"1d1208",x"1e1209",x"52493f",x"4f463d",x"4f463d",x"4f463d",x"000000",x"000000",x"000000",x"000000"),
(x"7b634f",x"7b6450",x"5d5145",x"56493b",x"4d3f32",x"514235",x"514234",x"4e3f32",x"4b3c2f",x"4b3d2f",x"49392b",x"4f3c2b",x"4c3a2c",x"503f30",x"514031",x"554231",x"5a4736",x"574535",x"564333",x"564332",x"584534",x"604a37",x"5b4736",x"5b4736",x"5a4636",x"574534",x"574434",x"574534",x"594635",x"5d4735",x"584534",x"5b4938",x"5c4a39",x"614d3c",x"614d3d",x"624e3c",x"5d4837",x"5f4935",x"614a35",x"5d4732",x"5f4732",x"5e4730",x"5c452f",x"5f4833",x"58402c",x"614a34",x"604833",x"624a34",x"674e37",x"664e38",x"604833",x"614a36",x"644e38",x"614935",x"584432",x"544130",x"584330",x"604832",x"5c4633",x"5b4632",x"5c4632",x"58432e",x"584330",x"564330",x"544130",x"584432",x"584230",x"5f4835",x"57422f",x"574332",x"564434",x"584636",x"584535",x"584534",x"534133",x"4d3c2e",x"47382a",x"4b3b2d",x"4d3c2d",x"534132",x"574738",x"594a3c",x"5c4c3e",x"5c4c3d",x"1f150b",x"1f150c",x"1e140b",x"1d140b",x"1d130a",x"1f150b",x"20150c",x"20150c",x"1f150b",x"1c130a",x"1d130a",x"21170d",x"271b10",x"291c11",x"2a1d11",x"302214",x"2c1e12",x"302215",x"3a291b",x"382819",x"3b2a1b",x"3d2c1c",x"382819",x"3e2c1d",x"3a2919",x"412f1f",x"42301f",x"402e1d",x"443220",x"402d1d",x"3f2d1b",x"3f2d1d",x"473321",x"453221",x"463220",x"45311f",x"422e1d",x"432f1d",x"432f1e",x"412e1d",x"3f2c1b",x"3e2a1a",x"412e1c",x"3e2c1b",x"422f1e",x"463220",x"45301f",x"493522",x"493422",x"4e3824",x"4c3825",x"4a3624",x"483422",x"483522",x"483623",x"463323",x"5d432e",x"1c160f",x"23190f",x"21170d",x"22180e",x"20160c",x"20150b",x"21160d",x"271b10",x"2f2115",x"291c11",x"2a1d11",x"24180e",x"24180d",x"291c11",x"271b10",x"291d11",x"271a0f",x"2c1f12",x"2c1f12",x"302114",x"332416",x"322315",x"382819",x"362618",x"352517",x"3d2c1d",x"412f1f",x"3d2b1c",x"3c2a1b",x"3f2d1d",x"3e2c1d",x"362617",x"3f2e1e",x"3f2d1d",x"422f1d",x"42301e",x"3f2c1c",x"3c2a1a",x"422f1e",x"43311f",x"42301f",x"3f2d1c",x"382718",x"3b291a",x"3e2c1b",x"3d2a1a",x"3d2b1b",x"3b2919",x"392717",x"3e2c1b",x"3d2c1b",x"5d432d",x"4d3825",x"191109",x"342517",x"3a2a1a",x"3b2a1a",x"3c2b1c",x"3d2c1d",x"291c11",x"150e07",x"150e07",x"24190f",x"281c10",x"24190f",x"2a1d11",x"24190e",x"2e2114",x"291c11",x"24190e",x"2c1e12",x"2d1f13",x"2d2013",x"2b1e12",x"2c1e12",x"291c10",x"2c1e12",x"271b10",x"2b1e11",x"281b10",x"291c10",x"2c1f12",x"291c11",x"2d1f13",x"2b1e12",x"2c1e12",x"302114",x"352618",x"352617",x"312316",x"362619",x"3b2a1b",x"332416",x"352517",x"352518",x"342416",x"302215",x"352517",x"352517",x"372819",x"372718",x"352517",x"342517",x"3a291a",x"372719",x"332416",x"332416",x"322215",x"302114",x"332315",x"322315",x"2f2113",x"332315",x"2a1d11",x"2f2014",x"312215",x"322316",x"312214",x"2e2013",x"342517",x"332416",x"342517",x"312316",x"2f2114",x"302214",x"2e2013",x"2e2014",x"2c1e12",x"2e2114",x"2e2014",x"302215",x"2c1f13",x"2b1d12",x"2b1e11",x"2c1e12",x"2d1f13",x"2d1f13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291a10",x"291a10",x"28180d",x"2d1c0f",x"2a190c",x"331d0d",x"1c1108",x"1c1108",x"1b1108",x"180f07",x"1d1108",x"1b1108",x"211309",x"2c180b",x"2f1a0b",x"2f190b",x"321c0c",x"331d0d",x"3a210f",x"3a2210",x"3a2210",x"3b2210",x"3c2310",x"391f0e",x"381f0d",x"38200e",x"381f0e",x"3a210f",x"371e0d",x"371e0d",x"381f0e",x"3c220f",x"351e0d",x"321b0b",x"2f190b",x"351e0d",x"351e0d",x"361e0d",x"351d0d",x"351e0d",x"3a200f",x"39200e",x"39200e",x"371f0d",x"391f0e",x"371f0e",x"381f0e",x"371e0d",x"361e0d",x"361e0d",x"341c0c",x"301a0b",x"341c0c",x"331c0d",x"341d0d",x"371f0e",x"38200e",x"341d0c",x"391f0d",x"3c210e",x"331c0b",x"361e0d",x"331c0d",x"381f0e",x"301a0b",x"2d190b",x"331d0d",x"371f0e",x"19130c",x"281a10",x"2a1b0f",x"2e1c10",x"291c12",x"221910",x"221910",x"4b2b14",x"4b2b14",x"3c2311",x"2c190b",x"2a180b",x"371f0e",x"351e0e",x"311c0c",x"361e0d",x"301a0b",x"29180a",x"2c180b",x"2f1b0c",x"1a130c",x"19130c",x"171009",x"1e1208",x"28170a",x"26160a",x"331c0d",x"341d0d",x"321c0c",x"29170a",x"281609",x"2e190b",x"341d0d",x"361e0e",x"351e0d",x"351d0d",x"351e0d",x"371f0e",x"341d0d",x"361e0d",x"381f0d",x"311b0c",x"361d0d",x"381f0d",x"3a210e",x"3a210f",x"3a200f",x"361e0d",x"371e0d",x"341c0c",x"361e0d",x"371f0d",x"311c0d",x"351e0e",x"3c2310",x"3b2310",x"38200f",x"39200f",x"351d0d",x"371f0e",x"361e0e",x"37200e",x"371f0e",x"301a0b",x"3a200e",x"38200e",x"331d0d",x"2f1a0b",x"301a0b",x"341d0c",x"331c0c",x"361e0d",x"381f0e",x"371f0e",x"371f0e",x"38200e",x"371f0e",x"341d0d",x"351d0d",x"331d0c",x"351d0d",x"17110a",x"25180e",x"2b1b10",x"312016",x"2c1e13",x"2b1d13",x"452711",x"3d220f",x"3e2410",x"3c230f",x"412712",x"3e2411",x"3b220f",x"3b210f",x"351d0d",x"3b220f",x"3d2410",x"412411",x"24150a",x"221409",x"544a3f",x"544b41",x"150e07",x"150e07",x"150e07",x"544b41",x"50463d",x"4e453c",x"4e453c",x"000000",x"000000",x"000000",x"000000"),
(x"6f5b4a",x"6d5947",x"584c3f",x"524438",x"504235",x"514336",x"4f4033",x"4a3b2e",x"4f4133",x"4f3f32",x"503f30",x"4e3d2d",x"513e2e",x"503e2e",x"564332",x"554535",x"5a4737",x"5b4736",x"594734",x"624b37",x"5b4635",x"5d4734",x"5b4633",x"604b38",x"5f4937",x"5a4532",x"5f4834",x"604936",x"5f4a37",x"614c3a",x"644f3d",x"5b4736",x"5d4835",x"624c38",x"604c3a",x"604b37",x"624b39",x"5c4734",x"5e4734",x"5f4631",x"654c34",x"604832",x"634b34",x"5d4733",x"634a33",x"634b33",x"664c35",x"664c34",x"684e36",x"684d36",x"674f3a",x"664e3a",x"674f3a",x"5b4635",x"624c36",x"5e4836",x"634b37",x"604834",x"624933",x"664e39",x"654b35",x"604a36",x"624a36",x"5a432f",x"57422e",x"5a4532",x"584432",x"5c452f",x"5a442f",x"5a4533",x"5c4836",x"594635",x"5c4938",x"564537",x"554331",x"4d3c2d",x"47372a",x"4a392b",x"4e3c2d",x"514031",x"544436",x"5d4c3d",x"614e3e",x"5f4d3d",x"20160c",x"1e150b",x"1e150b",x"1e140b",x"1e140b",x"20160c",x"20150c",x"1e150c",x"21160d",x"21170d",x"24190f",x"23180d",x"261a0e",x"291c10",x"2e2013",x"2e2014",x"312315",x"2f2114",x"362618",x"382819",x"3d2b1c",x"3b2a1b",x"402f1f",x"3d2c1c",x"402d1c",x"3f2d1d",x"43301f",x"422f1e",x"453221",x"433120",x"473322",x"493523",x"473321",x"4a3523",x"4c3623",x"473221",x"463220",x"44301e",x"422f1e",x"483423",x"4b3523",x"4a3523",x"4b3724",x"432f1c",x"412d1b",x"493320",x"4f3925",x"483422",x"483321",x"473221",x"4a3523",x"4c3623",x"4e3a27",x"4d3827",x"4f3b29",x"443323",x"58402b",x"1d1711",x"21180f",x"21170d",x"22180e",x"21170d",x"24190f",x"251a0f",x"261a0f",x"261b10",x"2a1d11",x"2b1e12",x"2a1d11",x"281c10",x"281b10",x"302215",x"2d1f13",x"2e2014",x"312216",x"2f2113",x"2f2113",x"342415",x"352517",x"352517",x"392819",x"3b2a1a",x"3b2a1b",x"3a291a",x"412f1f",x"402e1e",x"3f2e1e",x"3f2d1d",x"402d1c",x"3c2a1b",x"3e2c1c",x"3f2d1d",x"463321",x"412e1e",x"412e1e",x"3e2c1d",x"422f1e",x"42301f",x"3f2d1c",x"402e1d",x"45311f",x"432f1d",x"402d1c",x"453220",x"453120",x"443120",x"473322",x"3d2b1a",x"584028",x"4c3622",x"191109",x"392819",x"352517",x"382719",x"3a291a",x"3d2b1c",x"24190f",x"150e07",x"150e07",x"24190f",x"21160c",x"24190e",x"24190e",x"261a0f",x"302215",x"2f2115",x"2d1f13",x"2d2014",x"2c1e12",x"2a1d11",x"302214",x"322316",x"291d11",x"2c1f12",x"2d1f13",x"302215",x"2d1f13",x"2e2014",x"312216",x"2d1f11",x"2e2012",x"312114",x"332416",x"352517",x"312215",x"342416",x"352517",x"302215",x"362719",x"332517",x"37281a",x"362618",x"382718",x"382819",x"392819",x"392819",x"372719",x"372819",x"372819",x"3c2b1c",x"362617",x"392819",x"382819",x"3a291a",x"362617",x"342416",x"332416",x"352517",x"332416",x"352518",x"352618",x"322314",x"2e2012",x"312113",x"302214",x"352517",x"2f2014",x"322316",x"302214",x"302215",x"312316",x"312216",x"2e2114",x"2d1f13",x"322315",x"302214",x"332416",x"2e2013",x"302215",x"2f2115",x"2d2013",x"312316",x"2d2013",x"2d2013",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281a0f",x"281a0f",x"28190e",x"2c1b0f",x"29190c",x"2e1a0b",x"1e1208",x"1e1208",x"1c1108",x"180f07",x"1d1108",x"241509",x"241509",x"311b0c",x"311b0b",x"301b0b",x"2f1a0b",x"311b0c",x"301a0b",x"361e0d",x"341d0d",x"301b0b",x"341c0c",x"351d0c",x"321b0b",x"361e0d",x"38200e",x"3a210f",x"3c2210",x"3c220f",x"3a220f",x"3f2511",x"3f2511",x"38200e",x"3b220f",x"3a220f",x"3a210f",x"321c0c",x"301a0b",x"2d170a",x"321b0b",x"331c0c",x"361e0d",x"391f0e",x"3a200e",x"341d0c",x"351d0d",x"351d0c",x"351d0c",x"381f0e",x"3d2310",x"39210f",x"371f0d",x"361f0e",x"371f0d",x"351d0d",x"371f0e",x"371f0d",x"351d0d",x"351d0d",x"341d0c",x"391f0e",x"361e0d",x"361e0d",x"341d0d",x"2b180b",x"2e1a0b",x"341c0c",x"19130c",x"27190f",x"2d1c10",x"301e13",x"2d1d12",x"241910",x"241910",x"4a2a14",x"4a2a14",x"3a2210",x"311c0d",x"27160a",x"341d0d",x"3a200f",x"371f0e",x"361f0e",x"321b0c",x"2a180b",x"2d190b",x"311c0c",x"19120b",x"17100a",x"171009",x"1e1208",x"241509",x"221309",x"351e0d",x"311d0d",x"2a180b",x"301c0c",x"321d0d",x"301c0d",x"341e0e",x"331d0d",x"311c0c",x"301b0c",x"2f1a0c",x"2f1b0c",x"301c0c",x"321c0d",x"2e1a0c",x"311c0d",x"2f1a0b",x"321c0c",x"2f1a0c",x"331d0c",x"331d0d",x"2e1a0b",x"2f1b0c",x"321c0c",x"2c190b",x"2c180b",x"301b0c",x"2b180b",x"2d1a0b",x"2d190b",x"2c190b",x"28170a",x"2c190b",x"2b190b",x"2e1a0c",x"2b190b",x"311c0c",x"2f1b0c",x"2e1a0b",x"2f1a0c",x"2b180b",x"2e190b",x"301b0c",x"321c0c",x"2d190b",x"331d0d",x"301c0d",x"28170a",x"2e1a0b",x"301b0c",x"28160a",x"311c0c",x"2d190b",x"2d1a0b",x"301b0b",x"18110a",x"2a1a10",x"2e1f14",x"2f2015",x"2c2016",x"2a1d14",x"452611",x"3a200e",x"3b220f",x"361e0d",x"3c2310",x"3c210f",x"39210f",x"3e2310",x"351e0d",x"3d2310",x"3f2512",x"391f0d",x"391f0d",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"544b41",x"50463d",x"4e453c",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"695849",x"685647",x"5d5144",x"53473b",x"504337",x"4d3f33",x"4f4033",x"4a3d31",x"4b3c2f",x"4a3b2e",x"513f2f",x"4b3a2c",x"503f30",x"554233",x"534132",x"534030",x"584333",x"584332",x"574332",x"5a4633",x"5b4734",x"5f4935",x"5c4837",x"5a4533",x"594432",x"5c4734",x"5b4635",x"5e4837",x"604b38",x"624c38",x"5a4533",x"604935",x"5a4534",x"5f4936",x"5f4935",x"5b4634",x"5a4533",x"5e4733",x"5e4833",x"5b4532",x"5c4530",x"614832",x"5e4531",x"5f4732",x"5d4633",x"5e4530",x"5e4732",x"634932",x"654c34",x"604733",x"644b36",x"674f3a",x"644c38",x"604a37",x"634c38",x"5f4a36",x"624a35",x"684e38",x"634b35",x"644b37",x"614934",x"614a35",x"5c4735",x"614b38",x"574331",x"584331",x"5a4431",x"56412f",x"55412e",x"513d2d",x"574332",x"534131",x"594838",x"5c4a39",x"504030",x"4b3a2b",x"4e3d2d",x"4f3d2e",x"4d3c2d",x"4c3b2e",x"544435",x"5b493a",x"5e4d3f",x"5d4d3f",x"1d140b",x"1d140b",x"1d140b",x"20160c",x"20160c",x"1e140b",x"20160c",x"20160c",x"1e140b",x"21160d",x"1f150b",x"25190e",x"22170c",x"291c10",x"2e1f13",x"25190e",x"291c10",x"2f2013",x"302114",x"392819",x"3e2c1d",x"3d2b1b",x"402d1d",x"3d2a1b",x"422f1e",x"412e1e",x"44301f",x"43301e",x"422f1e",x"412e1d",x"43301f",x"45311f",x"463220",x"473220",x"4a3421",x"45301f",x"432f1e",x"483321",x"473221",x"463120",x"4a3623",x"483322",x"432f1d",x"432f1d",x"3d2a1a",x"412d1b",x"483321",x"432e1d",x"3f2c1b",x"422f1d",x"483321",x"493422",x"4e3926",x"4a3624",x"4a3625",x"473423",x"5c442d",x"1c160f",x"21180f",x"21180e",x"23180e",x"23180d",x"23180e",x"23180e",x"291d11",x"25190e",x"25190e",x"25190e",x"2a1d11",x"2b1e12",x"2c1e12",x"2c1e12",x"2b1e12",x"2f2114",x"2d1f11",x"2e2012",x"2d1f12",x"2e2012",x"332316",x"332315",x"302113",x"342416",x"3e2c1c",x"3c2a1b",x"3c2b1c",x"402d1d",x"402d1d",x"3a2819",x"3f2d1d",x"402d1d",x"3b2a1b",x"3b2a1a",x"422f1d",x"3f2c1c",x"3b2a1b",x"3d2b1b",x"43301f",x"3f2d1c",x"412e1d",x"412e1d",x"45301f",x"43301f",x"412e1d",x"3e2b1b",x"402e1e",x"43301f",x"412d1b",x"402d1c",x"543b26",x"45321e",x"191109",x"312214",x"2e2013",x"302114",x"382718",x"39281a",x"281c11",x"150e07",x"150e07",x"25190f",x"261a0f",x"261a0f",x"24180e",x"291c10",x"291c11",x"281c10",x"291c11",x"2b1e12",x"2d2013",x"312214",x"2e2013",x"2c1e12",x"2a1d11",x"2d1f13",x"2a1d11",x"2c1e12",x"2f2114",x"2d1f13",x"2c1e11",x"312114",x"281b0f",x"2d1f12",x"2f2114",x"2f2013",x"302113",x"2f2113",x"2d1f13",x"332416",x"332416",x"352617",x"342416",x"322316",x"362618",x"342416",x"362618",x"372718",x"372718",x"322316",x"332416",x"342516",x"342416",x"342416",x"362618",x"342416",x"322315",x"312316",x"2e2013",x"312214",x"332416",x"332416",x"342415",x"342315",x"302113",x"2d1e11",x"2f2114",x"2e1f13",x"322214",x"2b1e12",x"322215",x"2f2114",x"2e2014",x"2f2114",x"2f2114",x"312215",x"2a1d11",x"322315",x"302114",x"2b1d11",x"2b1d11",x"312215",x"2d1f13",x"2d2013",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"27190f",x"27190f",x"27190f",x"2a1a0e",x"2a1a0e",x"24150a",x"24150a",x"1d1208",x"1c1108",x"170f07",x"1b1008",x"1f1208",x"1e1208",x"170f07",x"180f08",x"150e07",x"180f08",x"170f07",x"170f07",x"1a1008",x"1a1008",x"1b1108",x"170f07",x"1b1008",x"1c1108",x"1f1309",x"1b1108",x"1e1208",x"1f1208",x"201309",x"1b1008",x"1f1309",x"1f1309",x"1f1309",x"221509",x"1e1208",x"1c1208",x"1d1209",x"180f08",x"1b1108",x"1b1108",x"1b1008",x"1f1209",x"1e1208",x"1e1208",x"1d1108",x"1d1209",x"1f1209",x"1b1008",x"170f07",x"1c1108",x"191008",x"150e07",x"150e07",x"160f07",x"160e07",x"1b1008",x"1c1108",x"191008",x"1c1108",x"1b1008",x"1f1209",x"1d1209",x"1c1108",x"190f08",x"191008",x"170f07",x"150e07",x"19120c",x"23170e",x"2e1c11",x"301d11",x"2c1d12",x"251911",x"251911",x"3e230f",x"402410",x"2d1a0c",x"2f1b0c",x"1e1108",x"371f0e",x"381f0e",x"38200e",x"371f0e",x"321c0c",x"29180b",x"2b180b",x"2f1c0d",x"171009",x"171009",x"150e07",x"1f1208",x"231409",x"211309",x"1d1108",x"170f07",x"1c1108",x"180f07",x"1b1108",x"180f08",x"150e07",x"180f07",x"1d1108",x"1d1108",x"170f07",x"1b1008",x"1d1108",x"1c1108",x"211309",x"1f1209",x"251509",x"1e1208",x"1d1108",x"1d1108",x"170f07",x"201208",x"231409",x"221409",x"221409",x"1d1208",x"1d1108",x"1f1208",x"170f07",x"150e07",x"1f1209",x"1d1208",x"211409",x"231409",x"150e07",x"170f07",x"191008",x"1b1008",x"150e07",x"1d1108",x"201309",x"26160a",x"1f1209",x"25160a",x"241509",x"24150a",x"201309",x"170f07",x"1c1108",x"180f08",x"201309",x"1f1208",x"1c1108",x"1a1008",x"1c1108",x"28170c",x"2b1b11",x"2f2016",x"312115",x"2f2117",x"241a12",x"462813",x"321c0d",x"351e0e",x"38200f",x"371f0e",x"3d2310",x"3d2311",x"3c2210",x"341c0c",x"3c220f",x"3e2310",x"391f0d",x"391f0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"645546",x"655649",x"5b4d41",x"584b3e",x"4f4235",x"4c3e32",x"4b3c2f",x"4d3e30",x"4c3d30",x"4c3d2f",x"4a3a2c",x"4c3b2c",x"4f3e31",x"4f3d2e",x"503e2e",x"513e2d",x"513f2e",x"56422f",x"594331",x"584331",x"5b4736",x"5b4633",x"5d4633",x"5e4834",x"5d4734",x"574332",x"594533",x"5c4735",x"624b37",x"614b39",x"604b37",x"5e4835",x"604a36",x"604a35",x"624b38",x"5e4834",x"5c4734",x"604a35",x"614934",x"5e4632",x"614a34",x"624932",x"5f4631",x"604832",x"5c442f",x"604630",x"5f4631",x"5e452f",x"634a33",x"644b36",x"634c37",x"644b34",x"634d3a",x"624b38",x"624b38",x"614b36",x"634c37",x"5d4935",x"614934",x"604731",x"624931",x"5f4936",x"604a35",x"5c4938",x"594532",x"584432",x"5c4733",x"574130",x"55412e",x"58432f",x"5a4534",x"5a4431",x"5e4a36",x"564536",x"503e2d",x"4b3b2c",x"4a3a2c",x"4c3a2b",x"4c392b",x"4c3c2d",x"514031",x"58483a",x"57493c",x"58493c",x"1f150b",x"1d140b",x"1c130a",x"1f150b",x"1d140b",x"1d140b",x"1f150b",x"1f150b",x"20160c",x"1f150c",x"1e140b",x"22170d",x"22170d",x"25190e",x"2a1d11",x"2a1d11",x"2a1d11",x"342416",x"362517",x"3a2819",x"3f2d1c",x"3e2b1c",x"3c2a1a",x"402e1d",x"3d2b1b",x"402d1c",x"412e1d",x"3e2b1b",x"432f1e",x"432f1e",x"432f1e",x"432f1f",x"473321",x"432f1e",x"412c1c",x"45311f",x"45301f",x"412e1d",x"402d1c",x"412e1c",x"422e1d",x"45301f",x"392818",x"3b2918",x"3f2c1b",x"412d1b",x"463220",x"432f1d",x"44301e",x"473220",x"483320",x"493421",x"4b3724",x"483423",x"443222",x"493624",x"5c432e",x"1d1710",x"231910",x"21170d",x"22170d",x"22170d",x"22170d",x"25190f",x"281c11",x"271b10",x"26190e",x"271a0f",x"2a1d11",x"271b10",x"281b10",x"281c10",x"2e1f13",x"2d1f13",x"2a1c10",x"2e1f12",x"2a1c10",x"322214",x"352517",x"342416",x"372617",x"3d2a1b",x"392819",x"3a2819",x"412e1e",x"3f2c1c",x"3c2a1a",x"402e1d",x"3b291a",x"402d1c",x"3c2a1a",x"3b291a",x"3c2a1b",x"3e2c1c",x"3e2c1c",x"3f2d1c",x"422f1e",x"3f2c1c",x"3d2a1a",x"3e2c1b",x"473220",x"402d1d",x"3a2819",x"3e2c1b",x"412d1d",x"3f2c1c",x"372717",x"3d2b1a",x"46321f",x"47331f",x"191009",x"332315",x"2f2013",x"362617",x"392819",x"3a2919",x"25190f",x"150e07",x"150e07",x"291c11",x"22170d",x"24180e",x"271b10",x"2c1e12",x"291c11",x"2a1d11",x"2c1e12",x"2a1d11",x"2e2014",x"2b1d11",x"2b1d11",x"2a1d11",x"2c1e12",x"2f2014",x"2a1d11",x"2e2013",x"2e1f13",x"342416",x"281b0f",x"2d1e11",x"2c1e11",x"2b1e11",x"2f2013",x"2e2013",x"322315",x"322315",x"322315",x"312215",x"3b2a1a",x"362517",x"302114",x"342517",x"342417",x"342416",x"362517",x"312215",x"352517",x"372618",x"352517",x"342417",x"372718",x"362517",x"322214",x"342416",x"322315",x"342417",x"2e2013",x"302114",x"342416",x"362517",x"2e1f12",x"2e2012",x"2f2013",x"2f2113",x"2c1e12",x"2f2113",x"2f2013",x"2c1e12",x"2e1f13",x"332416",x"322316",x"2a1d11",x"281b10",x"2e2014",x"2d1f12",x"291c10",x"2b1d11",x"312215",x"291c11",x"2c1e12",x"2b1e12",x"2a1d12",x"291d11",x"291d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24180f",x"24180f",x"241910",x"2a1a0e",x"2a1a0f",x"341e0f",x"2c190b",x"1e1208",x"1c1108",x"180f08",x"150e07",x"211409",x"27170b",x"2a190b",x"211409",x"25160a",x"25160a",x"26160a",x"221409",x"25160a",x"211409",x"25160a",x"27170a",x"27170a",x"25150a",x"27170a",x"201309",x"221409",x"26160a",x"2a190b",x"29170b",x"2d1a0c",x"2d1a0c",x"2c1a0b",x"2a180b",x"28170b",x"2d1a0c",x"27170a",x"28170a",x"28170a",x"27160a",x"241509",x"241509",x"28160a",x"251509",x"241409",x"241409",x"221309",x"231409",x"211309",x"1e1208",x"231509",x"180f07",x"1f1309",x"26160a",x"231409",x"26160a",x"28170a",x"231409",x"241409",x"241509",x"241509",x"26160a",x"27170a",x"1f1209",x"1f1209",x"1a1008",x"211309",x"26170b",x"26180d",x"2e1d11",x"301f13",x"2a1c11",x"1f1710",x"1f1710",x"523521",x"412511",x"2c190b",x"2e1b0c",x"241409",x"361f0e",x"361e0d",x"3a210f",x"39200e",x"321c0c",x"26160a",x"2a180b",x"351f0e",x"160f09",x"150e07",x"150e07",x"180f07",x"1d1108",x"1f1208",x"27160a",x"241509",x"211308",x"211308",x"211308",x"231409",x"251509",x"231409",x"241409",x"221309",x"241409",x"211309",x"251509",x"241509",x"28160a",x"29170a",x"27170a",x"27160a",x"28170b",x"2d1a0c",x"2c1a0b",x"2e1b0c",x"2b190b",x"2b190b",x"24150a",x"2a180b",x"27160a",x"27170a",x"1d1208",x"27170a",x"2a190b",x"27160a",x"231509",x"26160a",x"27160a",x"221409",x"1e1208",x"1f1309",x"28170a",x"2a180b",x"2e1a0c",x"2c1a0b",x"28170a",x"29180b",x"25160a",x"2d1a0c",x"2b190b",x"2a180b",x"29170a",x"241509",x"251509",x"27160a",x"241509",x"261509",x"211309",x"28180b",x"2c1d12",x"2c1e14",x"2c1f15",x"261d17",x"3d200d",x"3f2411",x"3a210f",x"3a210f",x"3c2310",x"361e0d",x"381f0e",x"402512",x"3e2411",x"331c0c",x"3b2210",x"381f0e",x"39200e",x"39200e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"665647",x"675748",x"5c4e42",x"57483c",x"514336",x"4d3e31",x"4c3d2f",x"4c3d2f",x"504132",x"514031",x"4e3e30",x"52402f",x"4f3c2c",x"513e2e",x"513d2d",x"513f2f",x"544232",x"53402d",x"584432",x"594433",x"614a37",x"5e4835",x"5e4936",x"5e4733",x"5b4532",x"5e4835",x"634a36",x"5c4733",x"614934",x"614b36",x"67503c",x"614a36",x"5e4937",x"644d39",x"644d3a",x"654d39",x"634b38",x"634c38",x"654d36",x"624a34",x"5d4730",x"5f4631",x"58422e",x"5f4630",x"5d4630",x"5b442e",x"58412d",x"584230",x"5c4731",x"604832",x"604933",x"614834",x"664f3a",x"634c3a",x"634d3a",x"674f3a",x"654d39",x"634b35",x"684f38",x"614a36",x"604935",x"624934",x"614a35",x"614b37",x"5f4b39",x"634c3a",x"5f4835",x"574231",x"5d4733",x"5f4935",x"604a36",x"584534",x"5b4937",x"5e4c3c",x"4f3e30",x"4c3b2c",x"4a3a2c",x"463729",x"473628",x"4c3b2d",x"504132",x"57483a",x"594a3c",x"594a3c",x"1e150b",x"1d140b",x"20160c",x"1d140b",x"1d140b",x"20160c",x"21160d",x"20150c",x"20150b",x"1f150b",x"251a0f",x"22170d",x"22170d",x"2b1e12",x"2c1e12",x"2f2014",x"2b1e11",x"342516",x"362618",x"3c2a1a",x"3b2a1a",x"3d2b1b",x"3c2a1a",x"3b2919",x"3e2c1b",x"3c2a1a",x"3d2a1a",x"3f2c1b",x"3d2b1b",x"3f2d1c",x"3f2d1c",x"44301f",x"44311f",x"453120",x"483321",x"45311f",x"473220",x"4a3522",x"4a3522",x"48331f",x"46311f",x"422e1c",x"4d3825",x"432f1e",x"463120",x"473221",x"493321",x"4a3422",x"473220",x"4f3925",x"4a3623",x"463220",x"453120",x"4d3725",x"453222",x"453221",x"5c432d",x"1d1710",x"21180f",x"23180e",x"1f150b",x"21170d",x"21170d",x"22170d",x"291d11",x"251a0f",x"281c10",x"2b1d11",x"2a1d11",x"2a1d11",x"2d2013",x"2b1e11",x"2d1f12",x"2a1d11",x"362619",x"322315",x"322315",x"342416",x"322315",x"3a291a",x"382718",x"3d2b1b",x"382819",x"3d2b1b",x"3b291a",x"3f2c1c",x"3a291a",x"3e2b1b",x"3e2d1b",x"3b2a1a",x"382617",x"332315",x"3a2919",x"3b291a",x"3c2a1a",x"3c2a1b",x"412e1e",x"3d2b1c",x"412e1d",x"402d1c",x"412d1d",x"412e1d",x"402d1d",x"3f2c1b",x"422e1d",x"3f2d1b",x"443120",x"402e1d",x"563c29",x"563e2a",x"191109",x"372718",x"352517",x"3a291a",x"3a291a",x"352517",x"271b0f",x"150e07",x"150e07",x"281b10",x"261a0f",x"23180d",x"271b10",x"2b1d11",x"281c10",x"291c10",x"2a1d11",x"2c1e12",x"2b1e12",x"2e2014",x"2e2013",x"312215",x"2a1d11",x"312215",x"322315",x"2f2013",x"322315",x"322214",x"372819",x"312215",x"2e2013",x"382719",x"382718",x"322315",x"352517",x"322316",x"362618",x"352517",x"342416",x"342416",x"362617",x"362617",x"352517",x"332315",x"322215",x"302114",x"352516",x"322315",x"342416",x"382718",x"352617",x"372718",x"342416",x"342516",x"2e1f13",x"362618",x"342416",x"342416",x"2f2013",x"2f2013",x"3a291a",x"312215",x"342416",x"362617",x"342416",x"342416",x"322215",x"342516",x"362618",x"312215",x"342416",x"322315",x"2d1f12",x"2d1f13",x"2e2013",x"2b1e11",x"2d1f13",x"2d1f13",x"2e2013",x"2c1f12",x"2f2013",x"2a1d11",x"2e2113",x"2e2113",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"20170e",x"20170e",x"21160e",x"25170d",x"27180d",x"301c0e",x"2c190b",x"1c1108",x"1b1008",x"180f07",x"150e07",x"1d1108",x"201208",x"1d1108",x"221409",x"201308",x"27160a",x"26160a",x"28170a",x"26160a",x"26160a",x"231409",x"231409",x"28160a",x"231409",x"261509",x"241509",x"251509",x"251509",x"2c190b",x"27160a",x"2a180a",x"2a170a",x"28160a",x"2b180a",x"271609",x"251509",x"241409",x"221208",x"201108",x"201108",x"271509",x"221309",x"251509",x"241409",x"251509",x"241409",x"29160a",x"281609",x"27160a",x"281609",x"201208",x"201208",x"1d1108",x"251509",x"231409",x"251509",x"251409",x"241409",x"27160a",x"28160a",x"241409",x"231409",x"2c190b",x"26160a",x"28170a",x"25160a",x"2b180b",x"2a190c",x"2f1c0f",x"2a1b10",x"2a1c11",x"261a11",x"1d160f",x"1d160f",x"4c2e1b",x"3d2310",x"2c190b",x"27160a",x"231409",x"361e0d",x"331c0d",x"38200e",x"361f0e",x"361f0e",x"221409",x"27170a",x"2f1c0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"1a1008",x"1e1108",x"1d1108",x"221409",x"231409",x"211308",x"1d1108",x"180f07",x"1c1108",x"1f1208",x"1c1108",x"241509",x"211308",x"1f1208",x"241409",x"231409",x"221409",x"231409",x"221409",x"251509",x"231409",x"231409",x"1d1108",x"221309",x"211309",x"261609",x"27160a",x"251509",x"231409",x"231409",x"231409",x"1d1108",x"1c1108",x"211309",x"221409",x"241409",x"201208",x"1b1108",x"251509",x"221409",x"26160a",x"201208",x"221309",x"201208",x"201208",x"1f1208",x"1e1108",x"1f1108",x"1c1007",x"201208",x"241409",x"231409",x"201208",x"231409",x"1f1208",x"21140a",x"231810",x"251b14",x"271e16",x"231d16",x"4a2a14",x"39200e",x"39200f",x"381f0e",x"351d0d",x"321b0c",x"3a210f",x"3e2310",x"3c210f",x"361e0d",x"3d2411",x"351d0d",x"3d220f",x"3d220f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"625244",x"625345",x"5b4f42",x"534438",x"4d3f31",x"4b3d30",x"4d3d30",x"4b3c2f",x"524132",x"514234",x"534131",x"514030",x"584331",x"523f2e",x"54402f",x"54402e",x"5a4533",x"5a4533",x"5a4532",x"5c4633",x"604a37",x"614b38",x"5e4936",x"604a36",x"604a36",x"5d4835",x"5b4531",x"654d39",x"654e38",x"68503a",x"604a36",x"664e38",x"664d37",x"5f4936",x"604935",x"624c38",x"634c37",x"5f4a36",x"644c36",x"644d39",x"6a5038",x"654e38",x"5c4632",x"614b35",x"644c36",x"674e36",x"5e4633",x"634b36",x"664e37",x"614934",x"5b4532",x"634934",x"644b35",x"664d36",x"68503b",x"674e39",x"6a513b",x"684f3a",x"664e3b",x"654d38",x"634d39",x"634d37",x"614a37",x"5f4836",x"5c4735",x"5b4633",x"5c4532",x"5c4632",x"5b4531",x"5b4633",x"5e4836",x"5e4b39",x"624f3d",x"5e4c3a",x"534333",x"513f30",x"4f3e2e",x"503e2e",x"4d3b2c",x"503e2e",x"564434",x"564638",x"5b4b3d",x"5b4c3e",x"1e150b",x"1d140b",x"1e140b",x"1e140b",x"1d140b",x"20160c",x"21160c",x"21160d",x"21170d",x"21170d",x"22180d",x"281b10",x"24180d",x"271b0f",x"271a0f",x"2d1f12",x"2b1e11",x"302114",x"382718",x"3e2c1c",x"402e1e",x"423120",x"43301f",x"402f1f",x"42301f",x"473322",x"422f1e",x"493422",x"473321",x"483421",x"412e1d",x"45311f",x"422f1e",x"473220",x"4a3522",x"4a3421",x"473320",x"4a3522",x"4b3622",x"493422",x"483421",x"4c3724",x"493421",x"4b3522",x"483320",x"45301e",x"3f2b1a",x"463220",x"44301e",x"432f1e",x"483321",x"4b3623",x"503b27",x"4c3a27",x"4d3927",x"4a3726",x"684e36",x"1d1610",x"231910",x"251a10",x"21160d",x"23180e",x"22170d",x"24190e",x"291c11",x"281c10",x"291d11",x"251a0f",x"291c10",x"291c10",x"2b1e12",x"322316",x"332416",x"332416",x"2c1e12",x"302114",x"342415",x"322214",x"332315",x"362617",x"392819",x"352516",x"3d2b1b",x"3e2c1c",x"473322",x"40301f",x"433120",x"402f1e",x"443120",x"43301f",x"3b2a1a",x"422f1e",x"3d2b1c",x"44311f",x"3a2819",x"3e2c1c",x"3f2d1c",x"44301f",x"43301f",x"43301e",x"43301e",x"3d2b1b",x"3e2c1c",x"402e1d",x"412f1e",x"412f1e",x"3c2a1b",x"3e2c1c",x"4e3824",x"4b3522",x"181008",x"352517",x"342416",x"342416",x"342416",x"382719",x"261a10",x"150e07",x"150e07",x"291d11",x"2c1f13",x"2c1f13",x"2c1f12",x"2c1e12",x"2b1e12",x"2f2114",x"281b10",x"302114",x"2d1f12",x"2e2013",x"322316",x"332416",x"342517",x"312215",x"322315",x"302114",x"362718",x"362618",x"2e1f13",x"302114",x"302114",x"2f2013",x"302013",x"322315",x"332315",x"302114",x"362618",x"39281a",x"3a291a",x"342618",x"362719",x"362718",x"3a2a1b",x"362719",x"342416",x"382819",x"3d2b1b",x"372718",x"352517",x"362617",x"312215",x"342416",x"382719",x"372718",x"312215",x"372718",x"382718",x"382819",x"352517",x"3a291a",x"362517",x"332316",x"322214",x"2f2013",x"302013",x"312215",x"312214",x"2d1f13",x"342416",x"342517",x"362619",x"342618",x"352618",x"302215",x"352518",x"352618",x"312215",x"302114",x"2f2114",x"2f2114",x"312215",x"2b1e11",x"2d1f12",x"2d1f12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d150d",x"1d150d",x"1f160f",x"20160e",x"27180e",x"2c1a0c",x"2d1a0c",x"1d1108",x"1b1008",x"180f07",x"150e07",x"150e07",x"150e07",x"191008",x"1d1208",x"1e1208",x"201309",x"1f1208",x"201309",x"221309",x"180f07",x"201309",x"221409",x"241509",x"201309",x"27160a",x"25150a",x"27160a",x"29170a",x"26160a",x"241509",x"241509",x"221409",x"27160a",x"221409",x"261609",x"231409",x"241509",x"251509",x"251509",x"211309",x"27160a",x"241509",x"241509",x"26160a",x"25150a",x"241509",x"28170a",x"241509",x"241509",x"231409",x"25150a",x"211409",x"29170b",x"29180b",x"26160a",x"1f1208",x"28170a",x"27170a",x"27160a",x"24150a",x"25160a",x"29180b",x"2b190b",x"2a180b",x"231409",x"231509",x"211309",x"1f130a",x"1f150d",x"1b150e",x"1d150d",x"1d1710",x"1d160f",x"1d160f",x"51301a",x"452812",x"311b0b",x"2c1a0b",x"231409",x"321c0c",x"361e0d",x"331c0c",x"3b210f",x"341e0e",x"1e1208",x"231409",x"29180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"170f07",x"1b1008",x"150e07",x"171009",x"1d160f",x"201a13",x"231c15",x"231d16",x"4d2c14",x"381f0e",x"381f0e",x"3a200f",x"351e0d",x"321b0b",x"3b2311",x"361e0e",x"361f0e",x"38200e",x"3b2311",x"341d0d",x"361d0c",x"361d0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"635344",x"685748",x"5d4e40",x"524336",x"4f4032",x"4a3d30",x"4e4032",x"514032",x"4f3f2f",x"5a4636",x"574434",x"514132",x"5b4533",x"54412f",x"554230",x"534030",x"5a4534",x"5a4535",x"5b4735",x"5e4836",x"634a37",x"5f4b38",x"664c38",x"624b38",x"604b37",x"644e3a",x"634c38",x"604936",x"684e35",x"684e36",x"664d36",x"684f39",x"69513a",x"674f3b",x"664f3b",x"674f3b",x"6a513d",x"6a513a",x"6e543d",x"67503a",x"664f39",x"67503b",x"664e3a",x"654d38",x"684f3a",x"634a35",x"654c37",x"614935",x"624a35",x"614934",x"614934",x"644a36",x"644b35",x"654b35",x"694e38",x"674e38",x"644b36",x"6a513c",x"634c38",x"664d38",x"684f3a",x"604936",x"604935",x"5f4733",x"604935",x"614a36",x"614a35",x"5d4734",x"674e38",x"654f3c",x"66513f",x"65513f",x"604c3b",x"5c4a39",x"5c4634",x"54402f",x"523f2f",x"503e2d",x"4f3d2d",x"513e2e",x"554436",x"59483a",x"5d4e40",x"5c4d3f",x"20150c",x"20150c",x"20160c",x"1e140b",x"1d140b",x"20160c",x"1d140b",x"20150c",x"21170d",x"21160c",x"22170d",x"281c10",x"291d11",x"291c11",x"2a1d11",x"312214",x"362617",x"342416",x"3f2d1d",x"3c2b1c",x"453221",x"412f1e",x"453221",x"473321",x"453120",x"432f1e",x"412f1e",x"432f1e",x"45311f",x"44311f",x"453120",x"432f1e",x"473320",x"44301f",x"483321",x"4a3422",x"483321",x"453120",x"4a3422",x"45311f",x"473320",x"473220",x"493320",x"493321",x"4e3824",x"4d3623",x"4a3421",x"493321",x"4f3824",x"4c3623",x"4e3825",x"4f3a27",x"4d3926",x"4f3a27",x"533c2a",x"4d3927",x"684d35",x"1d1710",x"241910",x"23180d",x"23180d",x"20160c",x"20160c",x"22170d",x"24190e",x"24190e",x"2a1d11",x"23180e",x"2d1f12",x"2b1e12",x"2b1e12",x"2d1f12",x"302214",x"322315",x"332315",x"2e2013",x"362617",x"352516",x"3b2919",x"362617",x"3a2819",x"3b291a",x"3f2d1d",x"412f1f",x"453221",x"433120",x"433120",x"3f2e1d",x"402e1d",x"3e2c1c",x"402d1d",x"3f2c1c",x"402d1c",x"3b2a1a",x"3c2a1b",x"432f1e",x"402d1c",x"3d2a1a",x"422e1d",x"453120",x"422f1d",x"44311f",x"432f1e",x"382618",x"42301e",x"3f2c1c",x"3d2b1a",x"3f2c1c",x"563f29",x"533c27",x"191109",x"372617",x"392819",x"382718",x"372719",x"3c2b1c",x"23180e",x"150e07",x"150e07",x"2a1d11",x"2b1e12",x"2a1d11",x"2f2114",x"281c10",x"251a0f",x"2d1f12",x"2d1f13",x"2b1e11",x"2d1f13",x"2d1f13",x"322315",x"2f2013",x"342516",x"342416",x"2f2114",x"2f2114",x"332416",x"362617",x"2e1f12",x"312214",x"2f2114",x"372718",x"342416",x"332315",x"3b2a1a",x"362617",x"3a291a",x"3a2a1b",x"362719",x"3a291a",x"372719",x"362718",x"372718",x"342416",x"39281a",x"342416",x"382818",x"342516",x"372718",x"362617",x"372618",x"332316",x"382718",x"372718",x"342516",x"342416",x"362617",x"332315",x"392819",x"342416",x"322215",x"362617",x"342416",x"392818",x"342416",x"372617",x"342416",x"2f2114",x"312216",x"372819",x"352618",x"372819",x"3a291a",x"302215",x"2e2013",x"2e2013",x"322316",x"2e2013",x"312215",x"2b1d11",x"2b1d12",x"302114",x"2e2013",x"2e2013",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"1c140d",x"20160e",x"28190e",x"2f1d0f",x"351f0f",x"1d1108",x"1a1008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a130c",x"1c150f",x"1b140e",x"1b140e",x"1c150e",x"1c150e",x"50321d",x"4a2c12",x"2e1b0b",x"301c0c",x"2b190b",x"331c0d",x"341d0d",x"2a160a",x"331d0c",x"3c2310",x"1a1008",x"1e1208",x"27170b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"1d1710",x"211b14",x"221b15",x"231c15",x"4d2c15",x"3a2110",x"3a210e",x"39210f",x"38200e",x"341d0c",x"3d2410",x"38200f",x"3d2411",x"331d0d",x"3e2512",x"371f0e",x"3a1f0d",x"3a1f0d",x"38200f",x"331d0d",x"361e0d",x"38200e",x"341c0c",x"39200e",x"371e0d",x"361f0d",x"3d230e",x"361e0d",x"3f230f",x"3e230f",x"000000",x"000000"),
(x"6b5949",x"6b5848",x"5d4e40",x"504236",x"4b3d31",x"47382b",x"4a3c2e",x"4d3d2f",x"534133",x"584536",x"554232",x"503f2f",x"5a4533",x"574331",x"564232",x"5b4734",x"5b4736",x"5c4835",x"5b4635",x"614b38",x"634d3a",x"654f3c",x"644e3a",x"644c38",x"695340",x"66503c",x"644d39",x"674e39",x"604835",x"624b36",x"644d38",x"664d38",x"68503a",x"654e3a",x"6b533e",x"69503b",x"674e39",x"664f3b",x"624d3c",x"6a513d",x"6b523b",x"6b533d",x"6c523c",x"624d39",x"6c523d",x"664e39",x"67503a",x"685039",x"6a503a",x"674e37",x"624933",x"664d37",x"694e36",x"694f37",x"6a5038",x"624b37",x"614936",x"604a36",x"634b36",x"654d37",x"604a36",x"624b36",x"634c38",x"5f4935",x"604934",x"614a35",x"5d4632",x"5b4532",x"5b4533",x"5d4836",x"5f4b39",x"644d3b",x"634e3b",x"5c4936",x"584534",x"4f3d2c",x"524030",x"4f3e2e",x"54402f",x"554232",x"574636",x"5b4b3b",x"615042",x"605041",x"1d140b",x"1e140b",x"20160c",x"1d140b",x"20150c",x"1d140b",x"20150c",x"20160c",x"20160c",x"20160c",x"23180d",x"281b10",x"291c11",x"2d1f12",x"291c11",x"302114",x"2c1d11",x"322214",x"352516",x"3e2c1c",x"402e1d",x"493523",x"453220",x"3f2d1c",x"483422",x"463220",x"45311f",x"4b3623",x"4a3624",x"493421",x"45301e",x"473221",x"483321",x"483422",x"4d3623",x"432f1e",x"45301f",x"45311f",x"463220",x"483421",x"4d3723",x"4a3522",x"4c3522",x"483320",x"4b3623",x"493421",x"4b3522",x"46321f",x"3e2a19",x"422d1c",x"45311f",x"4f3825",x"4e3825",x"503c29",x"4c3927",x"483423",x"6c5037",x"1c150e",x"271b11",x"24190e",x"22180e",x"23180d",x"20160c",x"23180e",x"291c11",x"261a0f",x"2a1d11",x"291c11",x"2d1f12",x"2b1e11",x"2e1f13",x"332416",x"312214",x"362618",x"342416",x"342416",x"352517",x"322315",x"322315",x"362617",x"322214",x"382617",x"372718",x"3f2d1c",x"422f1e",x"443120",x"402e1e",x"3a2819",x"43311f",x"3d2b1c",x"402e1d",x"3e2d1c",x"412f1f",x"3c2a1a",x"3d2b1b",x"3d2b1b",x"3f2c1c",x"402d1d",x"473220",x"402d1d",x"3c2a1a",x"412d1d",x"412d1c",x"3f2c1c",x"382718",x"432f1e",x"3d2b1c",x"3d2b1b",x"553e29",x"563e29",x"150e07",x"342416",x"2d1d11",x"302113",x"312214",x"392819",x"281c10",x"150e07",x"150e07",x"271a0f",x"271b10",x"2a1d11",x"302114",x"2f2114",x"312316",x"2d1f12",x"2e1f13",x"322316",x"2f2014",x"2d2013",x"342416",x"312215",x"2f2114",x"2d1f12",x"322315",x"332416",x"342416",x"362618",x"342416",x"362517",x"332416",x"342416",x"352517",x"312215",x"2e1d11",x"302113",x"352517",x"3a291a",x"362618",x"3a2a1b",x"3a2a1b",x"362617",x"3b2a1b",x"3a291a",x"342517",x"3d2c1c",x"3c2b1c",x"3a2919",x"362517",x"3f2c1c",x"372718",x"39281a",x"342416",x"362517",x"2d1f12",x"332315",x"332416",x"342516",x"342416",x"342416",x"362517",x"342416",x"372718",x"322315",x"322315",x"342415",x"28190e",x"322214",x"2f2013",x"322315",x"362618",x"362719",x"352517",x"302114",x"332517",x"332416",x"2e2013",x"332417",x"342517",x"2b1d11",x"2c1e12",x"2d2013",x"302214",x"302214",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b140d",x"1e150e",x"24170d",x"301e0f",x"341e0e",x"1c1008",x"1a1008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"19120b",x"1a140d",x"1b150e",x"1b140e",x"1c140e",x"2e1a0b",x"2b190a",x"492b13",x"3a230e",x"36200e",x"311d0c",x"311b0c",x"3a210f",x"2e190a",x"331c0c",x"3a220f",x"170f07",x"190f08",x"1a1108",x"180f07",x"211308",x"201309",x"221409",x"1f1208",x"1b1008",x"1a1007",x"1c1108",x"1d1108",x"1f1208",x"201308",x"201308",x"201309",x"1e1209",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"201309",x"1f1208",x"241409",x"1f1309",x"201209",x"221409",x"241509",x"221409",x"211309",x"201309",x"221409",x"201309",x"1f1309",x"201208",x"1d1108",x"231409",x"221409",x"231409",x"221409",x"1f1309",x"201309",x"211309",x"231409",x"26160a",x"23150a",x"201309",x"25160a",x"24150a",x"25150a",x"28170a",x"26160a",x"28180b",x"29180b",x"28180b",x"27170a",x"211409",x"26160a",x"25160a",x"22150a",x"23150a",x"25160a",x"23150a",x"23150a",x"2c1a0c",x"311d0d",x"37200f",x"37200f",x"331e0d",x"4b2b15",x"3a210f",x"38200e",x"3a210f",x"2e1a0b",x"351e0e",x"3d2410",x"3d2410",x"3e2512",x"361f0e",x"392210",x"3a210f",x"422511",x"2d1a0b",x"38200f",x"331d0d",x"361e0d",x"38200e",x"341c0c",x"39200e",x"371e0d",x"361f0d",x"3d230e",x"361e0d",x"3f230f",x"3e230f",x"3e230f",x"000000"),
(x"7f6651",x"826852",x"605143",x"56473a",x"514133",x"4d3d30",x"544333",x"4d3d30",x"554334",x"584635",x"5a4634",x"544130",x"503c2b",x"54402e",x"54412f",x"574330",x"5f4936",x"5d4836",x"5d4836",x"614b37",x"654e3a",x"654e3a",x"614b38",x"6b5542",x"69523f",x"664f3b",x"624c38",x"624b38",x"674e39",x"664e3a",x"68503c",x"715740",x"6c533d",x"6f553f",x"6f5640",x"6d543d",x"68513f",x"69513c",x"6e563f",x"6a533f",x"6d5640",x"6a513d",x"6d5440",x"69523e",x"69503c",x"644f3c",x"69523f",x"695039",x"6e543d",x"664d38",x"695039",x"654c36",x"6a4f36",x"6a4f36",x"684f38",x"674e38",x"654c36",x"604832",x"634c37",x"654d3a",x"664d37",x"654f3a",x"664f3b",x"695139",x"634c38",x"644b35",x"614a36",x"6a5139",x"604934",x"614b37",x"67513e",x"67503d",x"664f3b",x"5e4a38",x"5f4936",x"574330",x"4f3c2c",x"4e3b2c",x"4e3c2d",x"513f2f",x"554334",x"5d4c3c",x"645243",x"645242",x"20160c",x"20160c",x"1d140b",x"1e140b",x"1f150b",x"1f150b",x"20160c",x"20160c",x"21160d",x"21170d",x"24190f",x"2d1f13",x"2a1d12",x"332416",x"2f2115",x"312316",x"392819",x"3a2819",x"422f1f",x"422f1f",x"453220",x"43301f",x"473321",x"432f1d",x"3e2a1a",x"402d1c",x"46311f",x"45311f",x"4b3623",x"453220",x"4b3522",x"473220",x"473320",x"483321",x"483320",x"46311f",x"47321f",x"432f1d",x"493422",x"4e3724",x"4e3824",x"513b28",x"4f3a26",x"523b28",x"503b26",x"503b26",x"4f3926",x"533d28",x"4f3925",x"4e3824",x"4f3925",x"523b28",x"4d3825",x"503b27",x"503a28",x"493422",x"5a402b",x"1b150e",x"21170e",x"22170d",x"23180e",x"23180e",x"23180e",x"23180d",x"291c10",x"261a0f",x"281c10",x"2b1d11",x"2b1d11",x"2c1e12",x"2d1f13",x"2d1f13",x"322316",x"332417",x"362719",x"3c2b1c",x"392919",x"362718",x"3e2d1d",x"402e1d",x"412e1d",x"3c2a1a",x"453220",x"43301f",x"402e1e",x"412f1e",x"43301f",x"3f2d1c",x"3b2919",x"3c2a1a",x"3c2a1a",x"3b291a",x"3f2c1c",x"3f2d1c",x"402d1d",x"3d2b1b",x"3f2c1c",x"45311f",x"44301e",x"43301e",x"402d1c",x"3c2a1a",x"402d1d",x"43301f",x"43301f",x"443120",x"433120",x"463322",x"5a422b",x"5b432d",x"150e07",x"3d2b1c",x"3a291a",x"392818",x"3c2a1b",x"3c2b1c",x"24190f",x"150e07",x"150e07",x"2a1d11",x"23180d",x"281c10",x"281b10",x"291c11",x"2d2013",x"2d1f13",x"2f2014",x"2d1f12",x"332416",x"342516",x"342416",x"342516",x"2d1f12",x"342415",x"352617",x"312315",x"3a281a",x"362719",x"372719",x"352517",x"392819",x"3a2a1a",x"38281a",x"3d2b1c",x"3a291a",x"382718",x"3c2a1b",x"3c2b1c",x"3a291a",x"392819",x"3b2a1a",x"382718",x"332315",x"312214",x"382718",x"392819",x"3d2b1b",x"372718",x"372718",x"392818",x"3a2919",x"382819",x"362617",x"332316",x"342417",x"322214",x"322316",x"372718",x"382719",x"362719",x"3b2a1b",x"3b2a1a",x"3d2c1c",x"362718",x"38281a",x"3d2c1c",x"382819",x"342416",x"362618",x"362718",x"342517",x"302214",x"362617",x"312214",x"2f2013",x"2e2013",x"2d1f13",x"2b1e12",x"2f2114",x"2e2114",x"2b1d11",x"2d1f12",x"2e2013",x"2e2013",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24180e",x"24180e",x"1c150d",x"271a0f",x"291a0f",x"321e10",x"3b2211",x"3d210f",x"3e220e",x"412410",x"422410",x"442611",x"432510",x"3c200e",x"3a1f0d",x"40230e",x"442611",x"452712",x"482912",x"422510",x"412410",x"432510",x"432510",x"3c200d",x"3e210e",x"40230f",x"422510",x"452611",x"442511",x"452611",x"492913",x"482913",x"4c2b14",x"482913",x"472813",x"482913",x"4d2d15",x"4c2c14",x"482812",x"462711",x"4b2b14",x"432611",x"462914",x"442712",x"442712",x"3f2310",x"432611",x"402410",x"402410",x"452711",x"462712",x"452611",x"422410",x"422410",x"482912",x"472913",x"422411",x"482913",x"492a14",x"492a13",x"492a14",x"4a2b14",x"4a2b14",x"482913",x"4d2c15",x"4a2c15",x"4b2c15",x"4c2c15",x"492a14",x"4b2b15",x"4d2d16",x"492b14",x"402410",x"412511",x"472913",x"3f230f",x"3e240f",x"38210d",x"371f0d",x"331d0c",x"381f0e",x"361e0d",x"38200e",x"371f0e",x"381f0e",x"211309",x"1f1309",x"1d1108",x"2e1a0b",x"341d0d",x"351d0d",x"371e0d",x"381e0d",x"3c210e",x"3e230f",x"3f2310",x"3e220f",x"391f0d",x"381e0c",x"381e0d",x"381f0d",x"3a200e",x"381f0d",x"381f0d",x"3a200e",x"3a200e",x"3c210f",x"3d220f",x"3d220e",x"3b200d",x"3b200d",x"3a200e",x"381f0d",x"3f220f",x"3f230f",x"3d210e",x"3a200d",x"3b200d",x"442610",x"452711",x"452711",x"452611",x"432510",x"3d220f",x"3f230f",x"3b200d",x"391f0d",x"3b200e",x"442611",x"422511",x"3d210f",x"3b200e",x"412410",x"412511",x"442712",x"452712",x"442712",x"4a2a14",x"4a2a14",x"4a2a14",x"472812",x"452712",x"412411",x"4a2a14",x"462813",x"482a14",x"4a2812",x"432611",x"442712",x"492a13",x"492812",x"442611",x"462711",x"442611",x"3f230f",x"381f0e",x"3b200e",x"402510",x"39200e",x"371f0e",x"3f2411",x"3e220f",x"3e240f",x"3e2510",x"402510",x"442712",x"4c2c15",x"4e2d15",x"512f17",x"4d2d15",x"4b2c15",x"4d2d15",x"4c2d15",x"492b14",x"482a14",x"482a12",x"4b2d13",x"4e2e13",x"543213",x"4f2e13",x"4f2e13",x"000000"),
(x"826851",x"82674f",x"5f5043",x"534336",x"504133",x"493b2f",x"4c3c2e",x"534133",x"4b3b2e",x"4d3d2e",x"513f2e",x"523e2d",x"564231",x"523f2d",x"564230",x"5c4633",x"554332",x"594634",x"594433",x"5b4736",x"634c39",x"624e3b",x"69523f",x"6c5744",x"69513c",x"654e38",x"654e3b",x"644d39",x"654d38",x"634c38",x"674f3b",x"6b513c",x"71563e",x"66503c",x"69513c",x"684f3a",x"684f3a",x"69503a",x"6a513c",x"6a513c",x"6b523e",x"69513d",x"68503b",x"66503e",x"685241",x"675240",x"68503d",x"68513d",x"664e38",x"644d37",x"654c37",x"634b37",x"664d37",x"634b36",x"614a34",x"654d37",x"654c37",x"644c37",x"674d36",x"674e38",x"664e39",x"695039",x"6a503a",x"685039",x"664e38",x"5f4834",x"644c36",x"5d4633",x"5d4634",x"5d4734",x"604b38",x"644d3a",x"614a37",x"5a4735",x"5c4632",x"4e3c2d",x"513e2e",x"4f3c2d",x"4e3c2c",x"4f3d2d",x"513f31",x"574738",x"5d4c3e",x"604f40",x"1c130a",x"1c130a",x"1c130a",x"1d130a",x"1d140b",x"20150c",x"20160c",x"20160c",x"20160c",x"21170d",x"23180e",x"291d11",x"2c1f12",x"2c1f12",x"2e2013",x"302114",x"352517",x"342416",x"3c2a1a",x"3d2b1b",x"422e1d",x"402d1d",x"3f2d1c",x"3f2c1b",x"45311f",x"412e1d",x"422f1d",x"412e1d",x"432f1e",x"45311f",x"432e1d",x"432f1e",x"44301e",x"432f1e",x"432f1d",x"45311f",x"46311f",x"483320",x"4c3523",x"4c3623",x"4e3824",x"533c27",x"533b27",x"4a3522",x"473321",x"483321",x"4d3623",x"473220",x"4a3422",x"44311e",x"473321",x"4c3623",x"493421",x"483523",x"483422",x"433121",x"61472f",x"1c150e",x"20170d",x"22170d",x"1f150b",x"1f150b",x"20160c",x"23180d",x"21160c",x"281b10",x"261a0f",x"271b10",x"2b1e11",x"2d1f12",x"2e2013",x"2e2013",x"312215",x"322416",x"342416",x"322316",x"382819",x"382718",x"3d2a1b",x"372718",x"3c2a1a",x"382718",x"402d1c",x"3f2c1c",x"422e1d",x"3f2d1c",x"3e2c1b",x"3c2b1a",x"3a2819",x"3c2a1a",x"3c2a1a",x"392819",x"392819",x"3e2c1b",x"392718",x"392819",x"402d1c",x"3e2b1b",x"3d2b1a",x"3f2d1c",x"3d2b1a",x"3d2a1a",x"3a2819",x"3f2c1c",x"43301e",x"422f1e",x"473221",x"412e1e",x"553e29",x"563f29",x"150e07",x"332416",x"362618",x"342416",x"352517",x"372718",x"1e140b",x"150e07",x"150e07",x"291d11",x"22170d",x"281b10",x"2b1d11",x"291c11",x"281c10",x"2c1e12",x"2a1d11",x"2a1d11",x"2f2113",x"2a1d11",x"312214",x"332315",x"312215",x"312215",x"362618",x"312215",x"372718",x"342517",x"342416",x"362617",x"3a291a",x"382718",x"322316",x"372718",x"312215",x"332315",x"362618",x"392819",x"392819",x"362618",x"3a2819",x"392819",x"372618",x"302114",x"342417",x"332316",x"352516",x"352517",x"342416",x"332415",x"342516",x"2f2114",x"342416",x"362617",x"352517",x"352517",x"342416",x"382718",x"372718",x"3a291a",x"3d2b1b",x"3a281a",x"3a291a",x"3a2819",x"3a2819",x"322315",x"352517",x"332315",x"352517",x"322315",x"302114",x"322316",x"312215",x"312214",x"352517",x"2d1f13",x"2b1e12",x"302114",x"2c1e12",x"2e2013",x"291c10",x"2a1d11",x"2f2013",x"2f2013",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24170f",x"24170f",x"1f160f",x"291a0f",x"2d1c11",x"2c1a0e",x"311d0f",x"351d0e",x"341c0c",x"371f0d",x"351d0c",x"331c0c",x"391f0d",x"321a0b",x"321b0b",x"331b0b",x"341c0b",x"341d0c",x"3c220f",x"3c210f",x"3c220f",x"3b210e",x"39200e",x"3b210e",x"381e0d",x"3a200e",x"391f0e",x"3a200e",x"402410",x"412410",x"402510",x"422611",x"412612",x"402511",x"3d220f",x"2f180a",x"3c220f",x"3f2411",x"3c2310",x"3f2310",x"3d2310",x"39200e",x"3a200e",x"3d2411",x"402512",x"3f2511",x"3d2411",x"3e2411",x"412612",x"422613",x"402512",x"412512",x"472914",x"3b2210",x"39210f",x"3d2310",x"3f2410",x"3d2310",x"402511",x"3f2511",x"3e2410",x"412511",x"3e2310",x"3f2511",x"3d2310",x"3a210f",x"3a200e",x"361e0d",x"331c0c",x"39200e",x"38200f",x"37200f",x"3b220f",x"37200e",x"39210f",x"351e0e",x"321c0c",x"38200e",x"38200f",x"361f0e",x"39200f",x"371f0e",x"38200e",x"351e0d",x"361e0d",x"211309",x"1f1209",x"221409",x"27170a",x"29170a",x"2b180b",x"2f1b0c",x"301b0c",x"351d0d",x"341d0d",x"311b0c",x"341d0d",x"331d0c",x"311c0c",x"331d0d",x"331c0c",x"2e1a0b",x"301b0b",x"311b0b",x"2d190b",x"2d190b",x"341c0c",x"311b0b",x"301b0b",x"311b0b",x"2f1a0b",x"321b0c",x"2d190b",x"2d190b",x"331c0c",x"2f190a",x"361d0b",x"2c170a",x"321a0b",x"361e0d",x"371e0d",x"39200e",x"3c220f",x"3b210f",x"321c0c",x"341d0d",x"361d0d",x"351d0d",x"3a200f",x"331c0c",x"321c0d",x"3d220f",x"3c220f",x"3b210f",x"38200f",x"3c220f",x"3b210f",x"2f190b",x"311b0b",x"331d0e",x"39210f",x"3c2310",x"3e2410",x"3d2310",x"391f0e",x"3a210f",x"452914",x"3a2210",x"3a2210",x"3e2511",x"422612",x"402612",x"402511",x"3f2512",x"3b2210",x"3c2310",x"3d2310",x"412611",x"3f2410",x"412511",x"442712",x"442813",x"3f2410",x"3f2511",x"3a210e",x"3c230f",x"412510",x"422610",x"402510",x"39200d",x"3b210d",x"38200d",x"3b210e",x"3e2410",x"3a210e",x"3e240f",x"462a11",x"482b12",x"4a2c11",x"44290f",x"44290f",x"000000"),
(x"856b55",x"866b54",x"5b4c3f",x"564739",x"4f3f31",x"4f3f32",x"4b3d2f",x"4c3d2f",x"4b3a2c",x"524031",x"4f3d2f",x"564231",x"523f2e",x"584331",x"5f4733",x"584230",x"5a4431",x"5c4532",x"5d4836",x"5e4937",x"644d3a",x"664f3c",x"6a5341",x"6a5340",x"6a513d",x"664e3a",x"654d39",x"634d39",x"67503d",x"644c38",x"69503c",x"6c533b",x"6d523a",x"6a523d",x"684f3b",x"6d543e",x"68503b",x"6d533e",x"684f38",x"644c37",x"654e3a",x"654d38",x"644c38",x"5c4837",x"69523e",x"6a5340",x"6a513d",x"674f3b",x"684e39",x"674d36",x"684f38",x"664e38",x"654e3a",x"674e39",x"674e39",x"644c36",x"644b36",x"634c37",x"654c36",x"664e38",x"674e38",x"6a513b",x"6a5039",x"6d523a",x"684e37",x"634b35",x"674f39",x"614935",x"644c37",x"614a36",x"5c4734",x"5c4735",x"604a36",x"5c4837",x"574433",x"594331",x"523f2e",x"533f2f",x"564230",x"4f3d2e",x"503e30",x"554335",x"625143",x"625041",x"1c130a",x"181008",x"1d130a",x"1c130a",x"1c130a",x"1d130a",x"23180d",x"20160c",x"23180e",x"23180e",x"261a0f",x"291d11",x"2b1d11",x"2f2114",x"2e2013",x"332416",x"352517",x"3a2919",x"3c2a1a",x"3a291a",x"3f2c1b",x"412d1c",x"402d1c",x"422e1e",x"432f1e",x"493421",x"4a3522",x"442f1e",x"463120",x"46311f",x"45311e",x"45311f",x"422f1d",x"402c1b",x"44301e",x"412e1c",x"432f1d",x"483320",x"4d3723",x"4d3623",x"4d3724",x"4e3824",x"4c3623",x"4e3824",x"503925",x"493422",x"4a3522",x"4b3623",x"4b3523",x"473220",x"483320",x"4a3422",x"412e1d",x"473421",x"473321",x"493523",x"5d432d",x"1b150e",x"241a0f",x"21160c",x"22170d",x"21170c",x"21160c",x"24180e",x"21160c",x"281b0f",x"271b10",x"291c10",x"281b0f",x"281c10",x"2e2013",x"302114",x"312215",x"362617",x"352517",x"3a281a",x"3a2819",x"352517",x"3b291a",x"3e2b1a",x"3c2a1a",x"3f2c1c",x"3a2919",x"392819",x"3a2819",x"3e2c1b",x"3e2b1b",x"382718",x"402d1c",x"3d2b1b",x"3f2d1c",x"3d2a1a",x"3c2a1a",x"3b2919",x"3c291a",x"3f2d1c",x"3c2b1a",x"3f2b1a",x"45311f",x"3b2919",x"3b2819",x"3e2c1b",x"3e2b1b",x"432f1e",x"3f2c1c",x"43301f",x"483421",x"463220",x"543d27",x"523c28",x"150e07",x"352517",x"372718",x"382718",x"352516",x"372618",x"20160c",x"150e07",x"150e07",x"271b10",x"2a1d11",x"2c1e12",x"2c1f12",x"2b1e11",x"2f2114",x"302114",x"2e2013",x"2f2013",x"2f2113",x"291c10",x"2f2014",x"302113",x"302113",x"342416",x"362517",x"322215",x"352517",x"382719",x"362618",x"3b2a1a",x"3a2819",x"372718",x"342416",x"3b291a",x"3e2b1c",x"322315",x"362617",x"362517",x"362617",x"372617",x"372618",x"392819",x"3b291a",x"372718",x"3a2819",x"332315",x"352517",x"352516",x"362617",x"3a2919",x"332315",x"332214",x"362517",x"332314",x"332214",x"352517",x"382718",x"352517",x"392819",x"352617",x"362618",x"362617",x"362617",x"372718",x"382718",x"3b291a",x"372718",x"332416",x"312214",x"332315",x"2f2013",x"302115",x"2f2114",x"322316",x"342416",x"2e1f13",x"312215",x"2b1e12",x"312215",x"2e2013",x"2c1e12",x"2c1f12",x"2c1e12",x"2c1e12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24180f",x"24180f",x"24180f",x"281a0f",x"362212",x"2e1b0e",x"331e0f",x"351e0e",x"351d0d",x"371f0d",x"381f0e",x"331c0c",x"2f190a",x"31190a",x"351d0c",x"361d0c",x"371e0c",x"3a200e",x"371e0d",x"371e0d",x"3b210f",x"3d220f",x"3d220f",x"3a200e",x"3d230f",x"3b210f",x"3c220f",x"3e2310",x"402511",x"3e2410",x"3f2410",x"412511",x"3f2411",x"3a210e",x"402511",x"402511",x"3e2310",x"3d230f",x"402410",x"3e2310",x"3a200e",x"39200e",x"39200e",x"341d0d",x"3d2411",x"38200e",x"321b0c",x"3a200f",x"3c220f",x"3e2410",x"3c220f",x"3c2210",x"3a210f",x"391f0d",x"361d0c",x"311a0b",x"371e0d",x"361e0d",x"371e0d",x"391f0e",x"39200e",x"39200e",x"331d0c",x"381f0d",x"381f0d",x"351e0d",x"361e0d",x"311c0c",x"381f0d",x"361e0d",x"371e0d",x"341c0c",x"341c0d",x"321c0c",x"331c0d",x"311c0c",x"311c0c",x"311c0c",x"311c0c",x"2d190b",x"331c0c",x"311c0c",x"331c0c",x"341c0c",x"351d0d",x"1f1208",x"201308",x"1b1108",x"221409",x"2a180b",x"2f1b0c",x"311c0c",x"361e0d",x"37200d",x"361f0d",x"341d0c",x"311c0b",x"2d1a0b",x"381f0e",x"301b0c",x"331c0c",x"331d0c",x"301b0c",x"311b0c",x"321c0c",x"311c0c",x"371f0e",x"321c0c",x"351d0c",x"311b0b",x"301a0b",x"321c0c",x"331c0d",x"351d0c",x"2e190a",x"2e170a",x"321a0b",x"351d0c",x"361d0c",x"321b0c",x"321c0c",x"39200e",x"39200e",x"3b210e",x"381f0e",x"3c220f",x"331c0c",x"351e0d",x"3c220f",x"371f0e",x"3d2310",x"3e2310",x"402511",x"3d2310",x"3d2310",x"39200f",x"39200e",x"3b210f",x"3a220f",x"371f0e",x"371f0e",x"3c2210",x"3d210f",x"361e0d",x"3d2310",x"3a200f",x"3e2411",x"3f2411",x"331c0c",x"3a200e",x"422611",x"3e2411",x"3c220f",x"3c210f",x"3a210f",x"371f0e",x"351c0c",x"341c0b",x"3a200e",x"3a200e",x"39200e",x"3a200e",x"3e230f",x"3a200e",x"38200d",x"39200d",x"371f0d",x"371f0c",x"3b210e",x"3b210e",x"38200d",x"361f0c",x"39200e",x"371f0c",x"37200d",x"3d230e",x"3f250e",x"442810",x"492b11",x"43280f",x"43280f",x"000000"),
(x"866b54",x"8b6f57",x"5d4f42",x"534335",x"4d3e32",x"504032",x"514031",x"503e30",x"513f30",x"574433",x"594432",x"564332",x"5b4533",x"5e4735",x"5e4732",x"634c37",x"614b37",x"624b37",x"654e3b",x"5c4837",x"654e3a",x"69523e",x"6c543f",x"6a523d",x"674f3a",x"6c523a",x"634b36",x"624c3a",x"5d4736",x"69513d",x"6b533f",x"6e553f",x"68503b",x"6f553d",x"6c533c",x"6c533c",x"67503c",x"684e3a",x"684e39",x"614a36",x"5e4734",x"684f38",x"684f3a",x"654d39",x"654f3c",x"6a533f",x"6e543f",x"6b533d",x"70553d",x"695039",x"6f543c",x"664d35",x"664e3a",x"694f3a",x"6c513b",x"6c533d",x"69503b",x"684f39",x"674e39",x"644b37",x"634a34",x"6b5038",x"6c523a",x"6f553c",x"6a5038",x"674e39",x"674d38",x"624b36",x"594432",x"5f4732",x"604834",x"5e4936",x"5d4836",x"634d3a",x"5a4736",x"5b4531",x"5a4432",x"564231",x"554130",x"584533",x"584534",x"5a4839",x"665443",x"645242",x"1d140b",x"1d140b",x"1d140b",x"1d140b",x"1d140b",x"1f150c",x"1f150b",x"1e140b",x"1e140b",x"23180d",x"21160c",x"2c1f13",x"2c1f12",x"2d1f13",x"312316",x"342516",x"362517",x"3a291a",x"3c2a1a",x"3c2a1a",x"3d2a1a",x"402d1c",x"43301f",x"45301f",x"432f1e",x"4b3623",x"483321",x"4e3825",x"4c3723",x"4e3723",x"4c3723",x"422f1c",x"473220",x"493321",x"473220",x"4b3522",x"483421",x"493422",x"483320",x"442f1d",x"3c2919",x"4c3623",x"4c3623",x"553e2a",x"4d3723",x"4d3724",x"4b3623",x"4c3623",x"473220",x"463220",x"46321f",x"483320",x"422e1d",x"493623",x"4a3625",x"493524",x"664a33",x"1b140d",x"23180e",x"24190f",x"21160d",x"23180d",x"23180e",x"23180d",x"271b10",x"281c10",x"281b10",x"2c1e12",x"2b1e11",x"2b1e11",x"2a1d11",x"2e1f12",x"2a1c11",x"342517",x"3b291a",x"3d2c1c",x"342416",x"3a291a",x"39281a",x"3f2c1b",x"3a2819",x"3a291a",x"3e2c1b",x"3c2a19",x"3b2919",x"443120",x"443120",x"3d2a1a",x"43301f",x"44311f",x"44301f",x"402e1e",x"43301f",x"3d2b1b",x"412f1e",x"3e2b1a",x"3a2919",x"412e1d",x"3f2c1c",x"422f1e",x"3f2d1c",x"3c2a1a",x"3a2919",x"3c2919",x"372617",x"443120",x"463221",x"4a3625",x"503926",x"4c3725",x"23180e",x"322316",x"302215",x"342517",x"302214",x"312214",x"1f150b",x"150e07",x"150e07",x"2b1e11",x"312215",x"2f2114",x"2d1f13",x"312215",x"322316",x"322316",x"2f2114",x"2b1e11",x"2f2013",x"322316",x"332416",x"322215",x"312215",x"312215",x"362617",x"332315",x"2e1f13",x"342517",x"382718",x"3a291a",x"382718",x"372718",x"3b2a1b",x"382819",x"352517",x"362617",x"3a2919",x"362516",x"3a2819",x"3b2a1b",x"3b2a1b",x"392819",x"382819",x"3b291a",x"3b2a1a",x"402e1e",x"3c2b1b",x"3b2a1a",x"3b2a1a",x"382817",x"3a2819",x"382818",x"352517",x"392819",x"362617",x"362517",x"362517",x"332315",x"2f2013",x"362718",x"322316",x"352618",x"322316",x"372718",x"372718",x"382819",x"322215",x"342417",x"342416",x"342416",x"2e2013",x"382819",x"382818",x"312215",x"372718",x"352517",x"322316",x"2e2114",x"322315",x"2e2013",x"2f2114",x"291d10",x"2f2014",x"2f2014",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25190f",x"25190f",x"251910",x"2e1d11",x"301d11",x"362011",x"382111",x"351e0f",x"381f0e",x"39200f",x"351d0c",x"341d0c",x"351d0d",x"361d0c",x"341c0c",x"361d0c",x"371e0d",x"371e0d",x"351c0c",x"361e0c",x"371e0d",x"3a200e",x"391f0d",x"3b210f",x"3a200e",x"3b210e",x"361e0d",x"371e0d",x"361d0d",x"361d0d",x"3b210f",x"3b210f",x"3d230f",x"3b210f",x"371f0e",x"3c230f",x"371f0e",x"3b210f",x"3e2310",x"3d2210",x"3b210f",x"3a210f",x"3a210f",x"39200e",x"311a0b",x"3c220f",x"3c2310",x"3e2411",x"3f2411",x"3c220f",x"351e0e",x"3b210f",x"3b210f",x"3f2410",x"39200e",x"3b220f",x"39200e",x"3b220f",x"3b220f",x"3a200e",x"381f0e",x"3a200e",x"321b0c",x"371e0d",x"381f0e",x"371f0d",x"3a210e",x"3c220f",x"39200f",x"3b220f",x"39210f",x"3d2310",x"3e2310",x"331d0d",x"331d0d",x"311c0c",x"2c190b",x"2e1a0b",x"2e190b",x"28160a",x"301a0b",x"341d0c",x"321c0c",x"311b0c",x"311b0b",x"211409",x"1b1107",x"211308",x"241609",x"311c0c",x"331e0c",x"37200c",x"341f0c",x"36200c",x"3a220d",x"38200d",x"38200d",x"311d0c",x"351f0c",x"371f0d",x"361f0d",x"321c0c",x"331d0d",x"301b0c",x"331d0d",x"311b0c",x"2f1a0b",x"341d0c",x"351e0d",x"321c0c",x"331d0d",x"2f1b0b",x"2f1a0b",x"321c0c",x"311b0c",x"321b0c",x"311b0b",x"341c0c",x"321c0c",x"2f1a0b",x"301a0b",x"331c0c",x"331c0c",x"331c0c",x"301b0c",x"321c0c",x"321c0c",x"39200e",x"381f0e",x"371e0d",x"361d0d",x"361e0d",x"371f0d",x"39200e",x"3b210f",x"3b210f",x"361f0e",x"361f0e",x"341c0c",x"39200e",x"371f0e",x"3b210f",x"361d0d",x"39200f",x"381f0d",x"3b220f",x"361d0c",x"381f0e",x"3e2310",x"3f2411",x"3d2411",x"3a210f",x"3c2210",x"3d2310",x"3a210f",x"3c210f",x"3f2410",x"3e2310",x"3e230f",x"3b210f",x"3f2410",x"3c220f",x"381f0e",x"391f0e",x"371e0d",x"3a200e",x"3c210e",x"3c220e",x"3b210e",x"3d240f",x"3e240f",x"3f240f",x"3d230f",x"432711",x"402611",x"412610",x"422610",x"442810",x"45290f",x"43280f",x"43280f",x"000000"),
(x"715b48",x"6b5643",x"5b4c3e",x"544538",x"4f4031",x"534132",x"4f3f30",x"4f3c2e",x"503e2f",x"5b4633",x"5a4533",x"5f4936",x"5b4734",x"614b36",x"614a36",x"624a36",x"644c38",x"604936",x"634c38",x"5f4b38",x"67503d",x"6a523e",x"654d39",x"654e39",x"664e39",x"6c523c",x"664e3a",x"69513d",x"695340",x"66503d",x"68503d",x"644e3d",x"574433",x"5d4734",x"67513d",x"68503b",x"6a523d",x"6a503a",x"654d37",x"6b513a",x"694e36",x"6c5139",x"674e39",x"6d543c",x"6a513c",x"735941",x"705740",x"6a503a",x"6e533b",x"674e38",x"674e38",x"634b35",x"6a513a",x"6c523b",x"644a36",x"634c38",x"664c38",x"6b513a",x"6f543c",x"6c523a",x"654d38",x"674e38",x"664d38",x"634b36",x"57402d",x"553f2a",x"5b4532",x"594332",x"634a36",x"604834",x"5f4834",x"604834",x"614b38",x"5f4a38",x"5f4937",x"5d4936",x"5a4533",x"574331",x"574332",x"564230",x"584434",x"594536",x"614d3d",x"614f3f",x"1d140b",x"1d140b",x"1c130a",x"1c130a",x"1c130a",x"1d140b",x"1d140b",x"20160c",x"21160c",x"21160c",x"23170d",x"25190e",x"201409",x"211509",x"2f2013",x"352517",x"382718",x"3a2919",x"3b2919",x"3b291a",x"412e1d",x"463220",x"493422",x"4a3523",x"4b3623",x"483422",x"4b3623",x"493422",x"4c3624",x"473320",x"4b3522",x"45311d",x"4d3722",x"4d3723",x"422e1d",x"46311f",x"46311e",x"483320",x"4a3421",x"493421",x"44301e",x"473220",x"47311f",x"412d1c",x"301e0c",x"34210d",x"45301e",x"46321f",x"4c3623",x"473220",x"45311f",x"483320",x"442f1e",x"493423",x"4e3926",x"513c28",x"634832",x"1b150e",x"251a10",x"24180e",x"23180e",x"22170d",x"22170d",x"23180d",x"281c10",x"2c1f12",x"2a1d11",x"281b10",x"261a0f",x"2e1f13",x"302114",x"2e1f13",x"2f2013",x"332315",x"342416",x"312113",x"27180a",x"2a1a0a",x"3a2717",x"3b2817",x"3a2819",x"3a2919",x"3e2c1b",x"3f2d1c",x"412e1d",x"432f1e",x"402e1d",x"422f1e",x"422f1e",x"473322",x"412f1e",x"3f2d1c",x"43301e",x"3b2919",x"3c2a1a",x"3c2b19",x"442f1d",x"45311f",x"3c2919",x"3c2a1a",x"3c2b1a",x"412d1c",x"3f2c1c",x"3d2b1b",x"362617",x"3c2a1a",x"3b291a",x"382819",x"342111",x"382310",x"21160c",x"2f2013",x"332416",x"342416",x"2f2114",x"342416",x"23170d",x"150e07",x"150e07",x"302214",x"302114",x"302215",x"332416",x"362617",x"2e2013",x"312214",x"332316",x"2e2013",x"312114",x"342416",x"2e1f13",x"2f2013",x"332315",x"392819",x"372618",x"352517",x"352516",x"352516",x"312214",x"322215",x"25170a",x"27180b",x"342315",x"372618",x"362517",x"382718",x"352516",x"3a2819",x"3b2919",x"3b2a1a",x"3b2a1a",x"3f2d1d",x"402e1d",x"3e2c1d",x"3d2c1c",x"3a291a",x"3b2a1a",x"382617",x"3a2919",x"382717",x"392717",x"3a2819",x"332315",x"362617",x"362516",x"382718",x"322215",x"322215",x"342415",x"342416",x"312214",x"2f2013",x"24170a",x"28190b",x"322214",x"2f2014",x"322315",x"322315",x"352516",x"372617",x"322315",x"352617",x"3b2a1a",x"3a291a",x"362618",x"352618",x"362718",x"322316",x"322416",x"2f2013",x"322315",x"2b1d11",x"2f2013",x"2f2013",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26190f",x"26190f",x"27190f",x"2e1c11",x"301d11",x"321e0f",x"382011",x"361f0f",x"371f0d",x"341d0d",x"341d0c",x"351d0d",x"341d0d",x"361e0d",x"361d0d",x"351d0c",x"321b0b",x"2f190b",x"311a0b",x"30190a",x"311a0b",x"301a0a",x"311a0b",x"2f180a",x"3a200e",x"371f0d",x"39210f",x"3a200e",x"351d0c",x"2f190a",x"291508",x"251208",x"2e180a",x"30190b",x"321b0b",x"351d0c",x"331c0c",x"371e0d",x"3a200e",x"3b210f",x"3c220f",x"3c220f",x"39200e",x"381f0e",x"3a210f",x"3d2310",x"3c2210",x"3d2310",x"3d2310",x"3b2210",x"39200f",x"3c220f",x"3e2310",x"402511",x"3b220f",x"402511",x"3e2311",x"3b210f",x"3b210f",x"371f0e",x"3b200e",x"3a200e",x"351d0d",x"39200f",x"3e2310",x"3d2310",x"39200e",x"3a210f",x"3f2410",x"3f2410",x"3c230f",x"351e0d",x"3a200e",x"361e0d",x"341d0d",x"361e0d",x"331c0d",x"321c0c",x"2b180b",x"2a180a",x"351d0d",x"331d0c",x"2f190b",x"301a0b",x"341c0c",x"231509",x"1d1208",x"201308",x"29180b",x"311c0b",x"36200c",x"3a230d",x"3e250e",x"3f2610",x"3b230f",x"3c230e",x"351f0c",x"371f0d",x"3b220e",x"3c220f",x"361f0d",x"331c0c",x"331c0d",x"2e1a0b",x"2e1a0b",x"331c0c",x"321c0c",x"311b0b",x"331c0c",x"341d0c",x"321c0c",x"321c0c",x"311b0c",x"2e1a0b",x"2d190b",x"331c0c",x"301b0b",x"301b0b",x"2e1a0b",x"2e190a",x"2d180a",x"2b160a",x"2c180a",x"2c180a",x"2a1709",x"2b170a",x"2f1a0b",x"351e0d",x"351d0d",x"371e0d",x"38200e",x"2e190a",x"2c1609",x"271308",x"2b1609",x"2f190b",x"301a0b",x"311a0b",x"311b0b",x"361e0d",x"361e0d",x"351d0d",x"3d220f",x"3c220f",x"3b210f",x"381f0e",x"3c220f",x"3b210f",x"3b2210",x"3a220f",x"3d2411",x"3d2411",x"3b210f",x"3c220f",x"361f0e",x"3f2411",x"422611",x"412511",x"3e2410",x"3e2310",x"3c220f",x"3d220f",x"3e230f",x"3c210e",x"3a200e",x"3c220f",x"3f2511",x"3d2410",x"3d230f",x"3d230f",x"3c220f",x"3f2410",x"3f250f",x"3d230f",x"3c220e",x"3e230f",x"3e240f",x"41270f",x"482b10",x"462a10",x"462a10",x"000000"),
(x"856a53",x"8c7058",x"58493b",x"57483b",x"524335",x"4f3f30",x"554333",x"534232",x"513e2e",x"594634",x"5e4734",x"5d4733",x"604835",x"5f4935",x"604833",x"5e4935",x"614936",x"634c38",x"66503d",x"644e3c",x"6b533f",x"674f3a",x"69503b",x"694e39",x"6b513a",x"6b523b",x"6a533e",x"6e553e",x"6d5541",x"715a45",x"6d5743",x"644d39",x"684f39",x"6f5741",x"715841",x"6d5440",x"69523d",x"674e3a",x"6c523c",x"6b523c",x"6a513a",x"6c513a",x"6c523b",x"6c5139",x"6d533d",x"72573d",x"6b513c",x"6e543e",x"6b513b",x"6e533b",x"674e38",x"6a513c",x"6c5139",x"6a4e37",x"6a4f38",x"694f3a",x"6b503a",x"6c513b",x"6f533a",x"6f533a",x"6c513a",x"70553d",x"6c523b",x"634b38",x"634a35",x"68503b",x"674f3b",x"604836",x"614936",x"604a35",x"654c37",x"644c37",x"634c38",x"604b38",x"5d4836",x"5f4937",x"574333",x"584532",x"54402f",x"544231",x"554232",x"5b4736",x"614e3e",x"614f3e",x"1d140b",x"1d130a",x"1d140b",x"1d140b",x"1e140b",x"20160c",x"20160c",x"20160c",x"23180d",x"23180d",x"24180e",x"25190e",x"2a1d11",x"322316",x"352517",x"3a2919",x"3d2b1b",x"3b291a",x"412d1c",x"44311f",x"453120",x"453120",x"473321",x"493422",x"4b3623",x"4e3824",x"483321",x"483320",x"493421",x"4a3422",x"473320",x"4b3522",x"4a3421",x"493420",x"463220",x"463220",x"473320",x"4c3623",x"4b3623",x"493421",x"4e3723",x"45311f",x"46321f",x"402c1b",x"46311f",x"4f3825",x"4b3422",x"4b3522",x"4b3522",x"46321f",x"4f3824",x"4e3824",x"483321",x"4a3523",x"4b3625",x"4e3926",x"674b32",x"1c150e",x"21180e",x"20160c",x"20160c",x"21160c",x"21170c",x"25190e",x"25190e",x"271b0f",x"2b1e11",x"2d1f13",x"2e2013",x"2a1d11",x"2f2114",x"342416",x"342416",x"322315",x"382718",x"362516",x"3c2918",x"3e2c1a",x"3d2a1a",x"412d1c",x"392819",x"3c2a1a",x"3f2c1c",x"44311f",x"402e1d",x"43301e",x"45311f",x"4a3522",x"473321",x"412f1e",x"432f1e",x"3e2b1b",x"3b291a",x"44301f",x"3f2d1c",x"412e1d",x"3a2919",x"3f2d1c",x"402d1c",x"3c2a1a",x"3f2c1c",x"442f1f",x"43301f",x"3e2c1c",x"432f1e",x"412e1d",x"392819",x"3a2819",x"473321",x"553d29",x"22170d",x"312214",x"302114",x"302114",x"362617",x"382818",x"22170d",x"150e07",x"150e07",x"322316",x"322316",x"332416",x"312215",x"322315",x"312215",x"352517",x"2f2113",x"322315",x"362517",x"322315",x"332315",x"372718",x"382818",x"382718",x"372718",x"322316",x"382718",x"3b2919",x"3a2819",x"342315",x"372617",x"3b2a1a",x"382618",x"3a2819",x"3b291a",x"382718",x"3c2a1b",x"3d2b1b",x"3e2b1b",x"3b2a1a",x"3d2b1b",x"3d2b1b",x"3f2d1d",x"3f2d1d",x"3d2b1b",x"392818",x"3a2919",x"3c2a1b",x"3a2819",x"3d2a1b",x"392818",x"332315",x"362617",x"372718",x"342516",x"3a2819",x"392819",x"382718",x"392819",x"382718",x"312214",x"2f2013",x"312214",x"3d2b1b",x"362517",x"362617",x"362617",x"342416",x"362617",x"3a2919",x"332416",x"382818",x"382819",x"382719",x"322316",x"332416",x"332316",x"332315",x"332416",x"322315",x"2b1e11",x"2e2013",x"2f2114",x"2f2114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"3f2411",x"442712",x"472812",x"442711",x"462912",x"462711",x"41240f",x"3e220e",x"412410",x"482913",x"4c2b14",x"4a2b13",x"4c2c14",x"462711",x"472711",x"42240f",x"3f220f",x"432510",x"452611",x"3e210e",x"472711",x"482912",x"482912",x"452812",x"432410",x"3f230e",x"3f220e",x"422510",x"472812",x"462712",x"452712",x"452711",x"4e2f17",x"4a2c15",x"492a14",x"412410",x"3f230f",x"432611",x"422511",x"402310",x"402410",x"422511",x"452712",x"472a14",x"462813",x"482914",x"472813",x"462812",x"422611",x"462813",x"432611",x"442611",x"422511",x"442711",x"412511",x"3e230f",x"40230f",x"412510",x"422511",x"442611",x"432611",x"432711",x"432612",x"452712",x"452712",x"472914",x"472813",x"482913",x"462813",x"472913",x"412511",x"422511",x"442611",x"402310",x"3a200e",x"361e0d",x"361e0d",x"361d0d",x"3e2310",x"412611",x"3e2310",x"412511",x"442713",x"2c1b0b",x"341d0d",x"39210f",x"3a210f",x"3f2410",x"402510",x"412510",x"442711",x"442711",x"432610",x"432510",x"3f230f",x"432611",x"422611",x"402510",x"3e2310",x"3f2410",x"39200e",x"351d0d",x"341c0c",x"371e0d",x"391f0e",x"341d0d",x"351d0c",x"39200e",x"3d230f",x"3c220f",x"3b210e",x"391f0d",x"391f0d",x"3c210f",x"422511",x"422511",x"3f2410",x"402410",x"482a15",x"452813",x"472914",x"3e2210",x"3b1f0e",x"422511",x"412511",x"3f2310",x"412410",x"412411",x"422410",x"432712",x"432612",x"432611",x"432712",x"462813",x"432612",x"412511",x"442712",x"412511",x"3d2310",x"402511",x"412511",x"3b210e",x"3f230f",x"3e2310",x"432711",x"3f2410",x"412511",x"3f2410",x"412511",x"3f2411",x"422611",x"432612",x"402511",x"3d2310",x"3f2411",x"3e2310",x"3d2310",x"3b210f",x"3d220f",x"3a200e",x"361d0d",x"361c0c",x"321c0b",x"301a0b",x"3a200e",x"412511",x"442711",x"432712",x"4a2b15",x"462813",x"442611",x"442711",x"432611",x"452811",x"492a13",x"442711",x"4a2a12",x"4f2f12",x"4f2f12",x"000000"),
(x"876b54",x"8a6d55",x"615244",x"57483b",x"554537",x"534232",x"524131",x"554332",x"544130",x"584331",x"5f4832",x"5d4734",x"5a4431",x"5d4632",x"5e4734",x"624c36",x"634c37",x"634c38",x"6a513c",x"68503c",x"654e3b",x"69513d",x"6b513a",x"684f3a",x"684f39",x"6b523a",x"6f543b",x"715741",x"725944",x"745c47",x"705743",x"705844",x"6f5743",x"725945",x"6f5742",x"6c5440",x"725942",x"6f5640",x"6a523b",x"6e5440",x"6f543e",x"654c38",x"6a5039",x"70543d",x"664d38",x"6a5139",x"6d523b",x"71563c",x"70543c",x"6f543d",x"70553e",x"6c523b",x"6f533b",x"6a503a",x"6e543c",x"6b5036",x"674e38",x"685038",x"6b5139",x"6e5239",x"6c533d",x"6c513b",x"6a4f38",x"684e39",x"6a503b",x"674e39",x"6a503b",x"654e38",x"674d39",x"6a5139",x"644c36",x"624b36",x"674e39",x"5f4b39",x"5c4737",x"5c4735",x"594534",x"574332",x"55412e",x"554231",x"564332",x"5b4939",x"645140",x"635040",x"1a1109",x"1e140b",x"191109",x"1d130a",x"1d140b",x"1e140b",x"20160c",x"20160c",x"20160c",x"23180e",x"281c10",x"281c10",x"2b1d11",x"312215",x"342416",x"3a2819",x"402d1c",x"3b2a1a",x"402e1c",x"463220",x"422f1e",x"412d1d",x"45311f",x"483321",x"46311f",x"473220",x"483320",x"493421",x"483320",x"4d3724",x"4a3522",x"4c3623",x"4e3824",x"493422",x"493421",x"46311f",x"463220",x"4b3623",x"4c3522",x"4d3724",x"493422",x"4b3623",x"4a3521",x"483220",x"4d3723",x"4f3824",x"4d3723",x"432f1d",x"4f3825",x"4e3824",x"4a3521",x"463220",x"4d3724",x"4b3623",x"473422",x"4d3826",x"5d442d",x"1c150e",x"21180e",x"20160c",x"23180d",x"23180e",x"23180e",x"281c10",x"251a0f",x"2b1e12",x"281c10",x"2f2013",x"2b1e11",x"2f2114",x"312214",x"352617",x"372718",x"382819",x"3a2819",x"3c2a19",x"3d2b1a",x"3e2b1a",x"432f1c",x"3f2d1b",x"432f1e",x"44301f",x"45311f",x"412f1e",x"453120",x"422e1d",x"45301f",x"463220",x"422e1d",x"45301f",x"432f1e",x"43301e",x"3b2919",x"432f1e",x"43301f",x"473220",x"453120",x"3f2d1c",x"3f2d1c",x"3f2c1b",x"3d2a1a",x"3f2d1c",x"432f1d",x"43301f",x"483421",x"473321",x"44311f",x"3f2c1e",x"4f3925",x"543c28",x"241a0f",x"302114",x"322315",x"382718",x"312315",x"342516",x"1e140b",x"150e07",x"150e07",x"312214",x"2f2013",x"352517",x"322315",x"342516",x"2e2013",x"382718",x"362617",x"382718",x"332416",x"372718",x"362618",x"322315",x"352517",x"352617",x"382718",x"39281a",x"3a2919",x"3d2b1b",x"3d2b1b",x"3b2919",x"3c2a1a",x"3a2919",x"3d2b1b",x"3a2819",x"3e2c1c",x"3e2c1b",x"3e2c1b",x"3d2b1b",x"3a2919",x"3b291a",x"3d2a1a",x"3e2b1b",x"3c2a1a",x"3b291a",x"3c2a1b",x"3d2b1b",x"3b2919",x"412e1d",x"3d2b1b",x"3f2c1c",x"3c2a1b",x"3a291a",x"382718",x"312214",x"352517",x"382718",x"3a2819",x"382719",x"372718",x"382819",x"322315",x"312214",x"392818",x"3c2a1a",x"382718",x"352516",x"3b2a1a",x"3a2819",x"392818",x"3a281a",x"342516",x"352517",x"382718",x"342416",x"312215",x"342417",x"342416",x"312215",x"312214",x"322315",x"322316",x"2e2013",x"2f2114",x"2f2114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"301a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"191008",x"1c1108",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"170f07",x"150e07",x"170f07",x"180f07",x"150e07",x"150e07",x"150e07",x"1d1108",x"29170a",x"1b150e",x"19130c",x"17110a",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1b1008",x"1b1008",x"1b1108",x"1b1108",x"1c1108",x"1b1008",x"1c1108",x"1b1008",x"1b1108",x"1b1008",x"1a1008",x"1b1008",x"191008",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1b110a",x"1c130b",x"1e150e",x"1f1710",x"201912",x"1f1911",x"1f1811",x"1d160f",x"1b1108",x"311c0d",x"3d2211",x"150e07",x"311c0d",x"251509",x"1c1108",x"29170a",x"150e07",x"321c0c",x"150e07",x"2a180b",x"150e07",x"190f08",x"150e07",x"2d190b",x"150e07",x"2e1a0b",x"2d190b",x"361c0c",x"321c0b",x"301a0b",x"3a200e",x"412511",x"442711",x"432712",x"4a2b15",x"462813",x"442611",x"442711",x"432611",x"452811",x"492a13",x"442711",x"4a2a12",x"4f2f12",x"4f2f12",x"000000"),
(x"866a54",x"846a53",x"5d4e40",x"57473a",x"504134",x"514234",x"513f30",x"533f2f",x"534030",x"554130",x"604934",x"604a36",x"634b36",x"654c38",x"604834",x"654d39",x"6a513c",x"6c543f",x"6a523d",x"6c523c",x"6b533c",x"6f563f",x"6f553f",x"715840",x"73573f",x"6a513b",x"6c533b",x"6f543c",x"725843",x"6d5743",x"715a45",x"715741",x"6e5541",x"6c5440",x"6e5742",x"6e5642",x"6d5541",x"6b533f",x"69523d",x"6a523d",x"674f3b",x"6b533c",x"6e543e",x"6f543c",x"6f543d",x"70553d",x"71553d",x"755a42",x"755b43",x"745a43",x"715841",x"715640",x"73583f",x"77593f",x"6f543c",x"74593f",x"70553c",x"6e543e",x"6d533b",x"6b513a",x"6b5139",x"6a513c",x"6e523b",x"6a503a",x"664e38",x"664e39",x"634c36",x"654c38",x"634c38",x"614a36",x"614a34",x"604833",x"5e4733",x"634d38",x"604a38",x"5a4737",x"5c4837",x"5a4533",x"5a4633",x"594534",x"5e4b39",x"614f3f",x"675645",x"655343",x"191109",x"191109",x"1a1109",x"1f150c",x"1f150c",x"1e150b",x"1e150b",x"20160c",x"22170d",x"21160d",x"291c10",x"281c10",x"2d1f12",x"302114",x"352516",x"3a2919",x"3c2a1a",x"3a2919",x"3d2b19",x"442f1e",x"3f2c1b",x"4a3522",x"493421",x"4a3422",x"473221",x"4c3623",x"483422",x"4d3826",x"513b28",x"4d3825",x"4c3724",x"503925",x"4a3523",x"503a27",x"4e3926",x"503b27",x"4c3725",x"4f3925",x"4c3623",x"4a3421",x"463120",x"4a3522",x"493421",x"493321",x"4b3521",x"483320",x"44301e",x"483320",x"46311f",x"46311f",x"45311d",x"4c3522",x"46311f",x"493523",x"4a3523",x"493524",x"634931",x"1b140e",x"22180f",x"22170d",x"24190f",x"251a0f",x"24190f",x"2a1d11",x"261b10",x"2b1e12",x"302215",x"322416",x"2d2013",x"302215",x"302214",x"352516",x"382718",x"3b2a1a",x"3a2819",x"3b2919",x"382718",x"3a2818",x"3f2c1b",x"3d2b1a",x"3f2c1b",x"3c2a1a",x"392817",x"432f1d",x"3f2d1c",x"432f1d",x"46311f",x"453220",x"4b3623",x"4a3522",x"443120",x"493423",x"493523",x"463321",x"43301f",x"473320",x"412f1e",x"463321",x"422f1f",x"423120",x"422f1f",x"412f1e",x"473321",x"43301e",x"412e1d",x"422f1f",x"453121",x"402d1e",x"483321",x"513a26",x"20170d",x"2f2113",x"2f2013",x"322315",x"312213",x"322315",x"21160d",x"150e07",x"150e07",x"2d2013",x"322316",x"342416",x"352517",x"362619",x"3b2a1b",x"3a2a1b",x"372719",x"352517",x"392819",x"3c2b1c",x"3e2d1d",x"3d2c1c",x"3b2a1b",x"3c2b1b",x"382819",x"352517",x"3d2a1b",x"3c2b1b",x"3a2819",x"392819",x"372617",x"382718",x"362617",x"362616",x"392718",x"382718",x"3b2919",x"3d2a1b",x"3a2819",x"3e2c1b",x"3e2c1c",x"3c2b1b",x"3d2b1c",x"43301f",x"412f1e",x"3f2d1d",x"3e2d1d",x"3c2b1c",x"412f1e",x"3c2a1b",x"3d2c1c",x"3f2d1d",x"42301f",x"3f2d1d",x"392819",x"3c2b1b",x"382819",x"372718",x"362617",x"39281a",x"372618",x"312214",x"342416",x"372617",x"372718",x"332415",x"322315",x"372617",x"372617",x"382718",x"372617",x"382718",x"392819",x"39281a",x"3b2a1b",x"352617",x"352517",x"372719",x"312216",x"382819",x"332416",x"302214",x"332416",x"332416",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c1108",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f08",x"1c150e",x"19130c",x"18110a",x"160e07",x"160f07",x"170f07",x"180f07",x"180f07",x"180f08",x"180f08",x"191008",x"191008",x"180f08",x"180f07",x"170f07",x"180f08",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"180f07",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1c1108",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"1c1108",x"1c1108",x"190f07",x"1a1008",x"1a1008",x"1b1109",x"1e150d",x"201810",x"211a12",x"231c14",x"231c15",x"211a13",x"201812",x"1a1008",x"251509",x"3e2414",x"150e07",x"150e07",x"150e07",x"2f1a0b",x"1a1008",x"27160a",x"170f07",x"150e07",x"150e07",x"42240f",x"1d1108",x"150e07",x"2a1b12",x"150e07",x"150e07",x"221309",x"221309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"846851",x"856a52",x"605144",x"57483b",x"534436",x"534234",x"4d3d2f",x"503d2f",x"4e3c2c",x"513d2d",x"483527",x"463524",x"594330",x"5b4430",x"654b37",x"644c36",x"644c38",x"654c3a",x"694e39",x"6a513b",x"71563f",x"6c533b",x"6b523c",x"6f543d",x"72573f",x"6b503a",x"6b513b",x"6b513a",x"6a513c",x"6c5440",x"6f5742",x"6f5743",x"705843",x"745a44",x"6b543f",x"6c533e",x"6d543e",x"6e5540",x"6b5440",x"6a513c",x"674f3b",x"634c3a",x"5b4330",x"54412f",x"6a503b",x"6e5239",x"725640",x"765a43",x"71563e",x"6c523d",x"6d513b",x"6f533c",x"775a41",x"72563d",x"70533b",x"74563d",x"6b523b",x"6b5039",x"70533c",x"694e36",x"654b33",x"664c35",x"6a503a",x"6a4f39",x"6a503a",x"6b503a",x"6a503a",x"624b37",x"644d3a",x"674e39",x"614831",x"5d4735",x"5d4935",x"5d4734",x"4f3d30",x"4b3b2c",x"544232",x"574534",x"5a4534",x"584432",x"574535",x"5b493a",x"685747",x"695747",x"191109",x"191109",x"191109",x"191109",x"1e140b",x"191109",x"1d140b",x"1c130a",x"1e140b",x"1f150c",x"271b10",x"2a1d11",x"2d1f12",x"342416",x"372718",x"352416",x"392819",x"3c2a1a",x"3c2a1a",x"3a2818",x"422f1d",x"3b2919",x"311f10",x"301e0c",x"3e2b1a",x"402d1c",x"412e1e",x"412f1e",x"493421",x"44301f",x"44301e",x"4c3724",x"4a3624",x"4a3523",x"473321",x"4e3824",x"4a3522",x"4a3422",x"4a3422",x"422f1c",x"3f2b1b",x"412e1d",x"432f1e",x"463120",x"453120",x"432f1e",x"44301f",x"412d1c",x"3f2d1c",x"45311f",x"43301e",x"3f2b1a",x"3e2c1b",x"422e1e",x"382616",x"312112",x"4f3824",x"1b140d",x"20160d",x"1e140b",x"22170d",x"1f150c",x"20160c",x"261b10",x"2a1d11",x"2e2014",x"291d11",x"2b1e12",x"2f2114",x"2e2013",x"2b1d11",x"342415",x"312114",x"342417",x"362618",x"3e2b1b",x"3a2818",x"3e2b1b",x"3c2a1a",x"342415",x"352516",x"382819",x"3c2a1a",x"392717",x"362616",x"3a2819",x"312010",x"2e1c0b",x"3d2a1a",x"3d2b1b",x"3b291a",x"3b2a1b",x"3a2919",x"3c2a1a",x"3a2919",x"3f2e1e",x"412f1e",x"412f1e",x"3f2d1c",x"43301f",x"402e1d",x"3e2b1b",x"3d2b1a",x"3e2b1a",x"3b2819",x"3b2a1a",x"3a291a",x"3f2d1d",x"493423",x"59402a",x"20170e",x"291c10",x"2a1d11",x"342517",x"312214",x"322214",x"1f150b",x"150e07",x"150e07",x"231609",x"2f2013",x"2d1f12",x"382719",x"322316",x"362517",x"372618",x"382718",x"3b2a1b",x"3c2b1b",x"3a2a1a",x"3a291a",x"3d2b1b",x"3e2d1c",x"392819",x"372617",x"352516",x"352416",x"3a2919",x"3a2819",x"3c2a1b",x"392819",x"3a2919",x"382718",x"362616",x"362617",x"3d2b1b",x"392819",x"3a2818",x"392818",x"322215",x"2d1d0e",x"28190a",x"3a2819",x"3e2b1b",x"402e1e",x"3d2b1c",x"392819",x"3a291a",x"3a2919",x"453220",x"3f2d1d",x"3d2c1c",x"3b2a1a",x"402e1d",x"3b2a1a",x"362517",x"3b291a",x"362516",x"352416",x"372617",x"382719",x"392819",x"382718",x"3c2a1b",x"382718",x"352516",x"352516",x"372718",x"332415",x"382617",x"332415",x"312114",x"2a1b0d",x"24170a",x"302113",x"352517",x"332416",x"322316",x"322315",x"2f2114",x"322315",x"332417",x"332417",x"332417",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1008",x"1a1008",x"1d1209",x"150e07",x"180f07",x"150e07",x"150e07",x"191008",x"150e07",x"150e07",x"180f08",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"1b1108",x"1d1208",x"150e07",x"180f08",x"191008",x"1d1108",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"170f07",x"1a1008",x"1a1008",x"170f07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"180f07",x"150e07",x"170f07",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"1a1008",x"1a1008",x"150e07",x"1a1008",x"150e07",x"150e07",x"26160a",x"26160a",x"25160a",x"241509",x"231409",x"211309",x"221309",x"231409",x"25150a",x"26160a",x"26160a",x"26160a",x"251509",x"231409",x"28170b",x"26160a",x"26160a",x"26160a",x"26160a",x"27170a",x"27170a",x"27170a",x"27170a",x"27170a",x"28170b",x"26160a",x"25150a",x"241509",x"241409",x"231409",x"27170a",x"25150a",x"25150a",x"25150a",x"28170b",x"26160a",x"26160a",x"27160a",x"26160a",x"28170a",x"27170a",x"29180b",x"28170b",x"29180b",x"2a190b",x"2a190b",x"29180b",x"28170b",x"28170b",x"28180b",x"26150a",x"27160a",x"28170a",x"28180b",x"27160a",x"251509",x"28170b",x"25150a",x"241509",x"231409",x"231409",x"251509",x"251509",x"231409",x"211308",x"28170b",x"26160a",x"241509",x"231409",x"231409",x"221409",x"23150b",x"251910",x"261c14",x"292018",x"281f18",x"261f18",x"261f18",x"1c1108",x"27170a",x"412614",x"150e07",x"150e07",x"150e07",x"2a170a",x"1b1008",x"29170a",x"150e07",x"150e07",x"150e07",x"331d0d",x"201208",x"150e07",x"281b11",x"150e07",x"150e07",x"2f1b0c",x"2f1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"866a53",x"866a51",x"5e4f41",x"594a3c",x"554537",x"554334",x"534131",x"544131",x"564232",x"55402e",x"503c2c",x"513d2c",x"513d2c",x"56402d",x"5c4431",x"614934",x"614835",x"654d39",x"654d38",x"644c37",x"664e3a",x"694e3a",x"6d523b",x"6b513c",x"6c513a",x"6e543d",x"694f38",x"664f39",x"705741",x"725842",x"6d5541",x"705742",x"735841",x"6e5541",x"6d5541",x"705741",x"70553f",x"705740",x"6e553f",x"6d543f",x"705844",x"6d543e",x"624b37",x"68503b",x"664f3b",x"68503c",x"69513c",x"6a5441",x"6c533f",x"6f5640",x"6b533e",x"71563e",x"70553e",x"69503b",x"6f543b",x"6f523b",x"72553c",x"73563c",x"6c5139",x"74573e",x"6f543c",x"70563e",x"6d523c",x"6d5138",x"70543d",x"6d543f",x"694f39",x"6b523c",x"69503b",x"664e38",x"664d39",x"614a36",x"614b37",x"614a36",x"5e4937",x"594635",x"534132",x"513e2f",x"524030",x"4f3d2f",x"534031",x"5c4c3d",x"675748",x"665546",x"160f07",x"150e07",x"150e07",x"191109",x"191109",x"191109",x"1d130a",x"1e140b",x"1e140b",x"21170d",x"20160c",x"2b1d12",x"2e2014",x"312215",x"362617",x"372718",x"3a2919",x"3a2919",x"3e2b1b",x"3d2b1b",x"422f1f",x"3f2c1a",x"3a2818",x"3c2919",x"362516",x"362516",x"372617",x"372617",x"3c2a1a",x"3e2b1b",x"3d2c1b",x"422f1e",x"432f1e",x"3f2c1c",x"432f1e",x"412e1d",x"45311f",x"453120",x"422e1d",x"4a3522",x"3e2c1c",x"473321",x"422f1e",x"493422",x"443120",x"453120",x"45311f",x"463120",x"463220",x"44301f",x"432f1e",x"422f1e",x"453120",x"402e1c",x"3f2d1c",x"3a291b",x"4c3623",x"1a130c",x"1e140c",x"1e140b",x"1c130a",x"1f150b",x"1f150b",x"23180d",x"291d11",x"291c11",x"291d11",x"2c1e12",x"2c1f12",x"2d1f13",x"312214",x"362617",x"312315",x"392819",x"372718",x"3a291a",x"3a291a",x"3c2b1b",x"3b291a",x"3c2a1b",x"3c2a1b",x"3a2919",x"3a2919",x"3b2a1a",x"3f2c1d",x"3b2918",x"3a2817",x"372617",x"362516",x"382617",x"352416",x"362516",x"362617",x"382819",x"372718",x"392819",x"3d2b1b",x"3a291a",x"402d1c",x"372618",x"3b2a1a",x"43301f",x"372618",x"402d1d",x"3a291a",x"412e1e",x"3d2b1c",x"3c2b1c",x"493624",x"58402b",x"1d140b",x"2c1e12",x"302114",x"322315",x"322315",x"332316",x"1c130a",x"150e07",x"150e07",x"2c1e12",x"2c1e11",x"2d1f11",x"2c1e12",x"312214",x"2f2013",x"332415",x"312215",x"372718",x"352517",x"362517",x"362618",x"352517",x"3d2b1b",x"3b2a1b",x"382718",x"3d2b1b",x"3d2c1c",x"3d2b1c",x"3e2b1c",x"3c2a1b",x"3a291a",x"3a291a",x"382718",x"392819",x"3a2919",x"392819",x"3f2c1c",x"402d1c",x"3b2a1a",x"382817",x"3a2919",x"332315",x"362516",x"352415",x"352416",x"362516",x"382818",x"3a2919",x"3c2a1a",x"372718",x"3b2a1a",x"362617",x"362618",x"3a2819",x"3b2a1a",x"3b2a1b",x"392819",x"3d2b1b",x"3a291a",x"3f2d1d",x"392819",x"3a291a",x"3a291a",x"3b2a1b",x"362617",x"392819",x"392819",x"392819",x"392819",x"382718",x"382719",x"352515",x"352516",x"2e1f13",x"2f2013",x"2f2012",x"2f2013",x"332315",x"2d2013",x"2f2114",x"332416",x"312214",x"332416",x"332416",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"24150a",x"201309",x"201309",x"24150a",x"1d1208",x"1d1108",x"201309",x"201309",x"201309",x"211409",x"201309",x"211409",x"231509",x"201309",x"1f1209",x"1f1208",x"211409",x"221309",x"251509",x"221409",x"241509",x"211309",x"201308",x"241509",x"231409",x"1f1208",x"201208",x"211309",x"1f1208",x"1d1108",x"1c1108",x"1c1108",x"150e07",x"150e07",x"1a1008",x"1e1208",x"1c1108",x"231509",x"1e1208",x"1a1008",x"211309",x"1c1108",x"201309",x"1f1208",x"1f1208",x"1d1108",x"150e07",x"1e1208",x"170f07",x"221409",x"211309",x"1f1209",x"221409",x"24150a",x"221409",x"221409",x"211409",x"1a1008",x"1d1208",x"150e07",x"150e07",x"150e07",x"27170a",x"27170a",x"27160a",x"26160a",x"241509",x"231409",x"241509",x"241509",x"241509",x"241509",x"25150a",x"231409",x"241509",x"241509",x"25150a",x"25150a",x"241509",x"241509",x"25160a",x"241509",x"241509",x"26160a",x"25150a",x"25160a",x"27170a",x"25160a",x"26160a",x"241509",x"25150a",x"241509",x"26160a",x"25160a",x"26160a",x"27170a",x"27170a",x"27170b",x"27170b",x"27170a",x"28170b",x"28180b",x"29180b",x"28170b",x"27170a",x"28170b",x"28180b",x"27170a",x"28180b",x"28170b",x"28170b",x"29180b",x"27160a",x"27160a",x"27170b",x"28170b",x"27160a",x"28170b",x"27170a",x"231409",x"231409",x"211308",x"261509",x"231409",x"261609",x"241509",x"261609",x"251509",x"231409",x"231409",x"221409",x"221309",x"211309",x"211409",x"23150b",x"23170f",x"261b12",x"261c14",x"271d16",x"221b15",x"1c1108",x"26160a",x"452815",x"150e07",x"150e07",x"150e07",x"2c190b",x"1c1108",x"261509",x"150e07",x"150e07",x"150e07",x"2c180b",x"201309",x"150e07",x"2b1c12",x"150e07",x"150e07",x"331d0d",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"866b54",x"876b54",x"5d4f42",x"5b4d3f",x"544437",x"534233",x"554232",x"574332",x"513f2d",x"55402f",x"584331",x"594431",x"624b36",x"624832",x"684f36",x"6b5139",x"6f543e",x"71563f",x"6b533e",x"6f533c",x"735841",x"735a44",x"765d45",x"725841",x"6b533d",x"6a513a",x"6b513c",x"553f2d",x"664c39",x"6e533d",x"6d543e",x"70553f",x"715741",x"70563f",x"745941",x"765b43",x"725740",x"735843",x"745a43",x"715740",x"6e543d",x"68503b",x"70563f",x"755b44",x"765b45",x"745942",x"775d46",x"7a5d45",x"7b604a",x"765c46",x"735944",x"725741",x"785c44",x"785c42",x"785c42",x"715740",x"6b513a",x"6b533d",x"6c513b",x"57412e",x"684e38",x"6c5038",x"6c523a",x"6f533c",x"70553e",x"6e543e",x"71563f",x"6d533d",x"69513c",x"6d543f",x"6e533d",x"69503b",x"614a35",x"614a36",x"664f3b",x"624d3b",x"5d4a39",x"5a4736",x"5a4635",x"594534",x"5c4838",x"5f4c3c",x"675647",x"675647",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181008",x"181008",x"170f07",x"181008",x"1d140b",x"24180e",x"281c10",x"2a1d11",x"2d1f13",x"2f2114",x"342517",x"372718",x"3a2a1b",x"39291a",x"3a2a1b",x"372616",x"322214",x"382718",x"3a291a",x"402e1d",x"3d2b1c",x"3d2c1c",x"3f2d1d",x"3e2c1d",x"3d2b1c",x"3f2c1c",x"422f1f",x"422f1f",x"433020",x"433020",x"3b2a1a",x"3d2b1b",x"372718",x"3b2919",x"2b1b0c",x"372517",x"3f2d1c",x"382718",x"3f2d1c",x"422f1e",x"3d2b1c",x"412e1e",x"422f1e",x"402d1d",x"412f1f",x"473322",x"443120",x"382717",x"3c2a1a",x"3e2c1d",x"412f1f",x"513b28",x"19130c",x"1b130b",x"1e150b",x"21170d",x"1e150b",x"20160c",x"20160d",x"2a1e12",x"2b1e13",x"2b1e12",x"2b1e12",x"2b1e11",x"2c1e12",x"2d1f13",x"24160a",x"302114",x"342517",x"342416",x"362618",x"3a291a",x"3d2b1c",x"3b2a1b",x"3b2a1b",x"352517",x"3a2a1b",x"3e2c1d",x"3d2c1d",x"3b2919",x"362616",x"382719",x"3b2a1b",x"3b2a1b",x"3a291a",x"443120",x"422f1e",x"402d1e",x"3a291a",x"3b2a1b",x"402d1d",x"3e2d1d",x"412f1f",x"443120",x"3c2b1b",x"3c2a1a",x"362617",x"382718",x"27180b",x"332315",x"382819",x"362517",x"3b2a1b",x"4b3725",x"5d432d",x"1e140b",x"2e2013",x"2d1f13",x"302215",x"302216",x"332417",x"150e07",x"150e07",x"150e07",x"362618",x"322316",x"352517",x"352517",x"382819",x"332417",x"392819",x"382818",x"39281a",x"3e2d1d",x"3e2d1d",x"433020",x"3b2a1a",x"3a291a",x"392819",x"352516",x"29190b",x"342416",x"392819",x"382718",x"3b291a",x"3b2a1b",x"3b2a1b",x"3b291a",x"3a291a",x"342517",x"42301f",x"3e2c1d",x"412f1f",x"3d2a1a",x"382616",x"3b291b",x"402d1d",x"412e1e",x"422f1e",x"412f1e",x"44311f",x"43301f",x"3f2d1d",x"402d1c",x"432f1f",x"402e1e",x"3e2d1d",x"3f2d1d",x"3c2b1b",x"372618",x"372718",x"3a2919",x"2b1b0c",x"332315",x"372718",x"382718",x"382718",x"3b2a1b",x"3a2919",x"3b291a",x"3f2d1d",x"3a291a",x"39291a",x"3c2b1c",x"3a291a",x"3b2919",x"382717",x"382718",x"382719",x"382719",x"332416",x"392819",x"382819",x"39291a",x"362618",x"362618",x"342416",x"372719",x"372719",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"24150a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"150e07",x"150e07",x"170f07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"180f08",x"191008",x"150e07",x"28180b",x"27170a",x"27170a",x"25160a",x"2a190b",x"191008",x"190f08",x"191008",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"190f08",x"190f07",x"1b1008",x"1c1108",x"1d1108",x"1d1208",x"1c1108",x"1e1208",x"1e1208",x"1f1208",x"1f1209",x"1f1208",x"201309",x"201309",x"1f1209",x"1f1309",x"1e1208",x"1f1309",x"201309",x"201409",x"201309",x"1f1309",x"201309",x"211409",x"211409",x"211409",x"211409",x"211409",x"211409",x"211409",x"211409",x"22140a",x"23150a",x"23150a",x"23150a",x"23150a",x"23150a",x"221409",x"221409",x"211309",x"1c1108",x"1e1208",x"1c1108",x"1c1008",x"1c1108",x"1a1007",x"1a1008",x"190f07",x"190f07",x"191008",x"191008",x"180f08",x"180f08",x"170f07",x"170f07",x"170f07",x"2c190b",x"201309",x"20140b",x"23180f",x"221810",x"221911",x"1d1710",x"1d1108",x"25160a",x"472916",x"150e07",x"150e07",x"150e07",x"301c0d",x"1d1208",x"2d1a0c",x"150e07",x"150e07",x"150e07",x"311c0c",x"1c1108",x"150e07",x"291b11",x"150e07",x"150e07",x"311b0c",x"311b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"7f6650",x"826750",x"5b4c3e",x"5a4a3c",x"574637",x"554435",x"564333",x"594532",x"58422d",x"58422f",x"5b4431",x"5b4532",x"5c4532",x"604733",x"654b33",x"634b36",x"69503b",x"6c523e",x"6c543e",x"6c523d",x"6d543e",x"745c46",x"715743",x"735943",x"705540",x"6e553e",x"6e543d",x"6b513a",x"70563e",x"715641",x"715740",x"6a513a",x"735841",x"6d543e",x"6f553e",x"71563f",x"755840",x"71573f",x"715740",x"745842",x"6e543d",x"6d533b",x"6f5641",x"6f553f",x"6b523e",x"6d533c",x"715740",x"735841",x"715741",x"755943",x"745b43",x"785c44",x"745941",x"785e46",x"70553f",x"72563e",x"735741",x"6e543d",x"725640",x"6b523c",x"71563f",x"70543d",x"6e543d",x"6b513a",x"745a41",x"6d533e",x"674e3a",x"6d533d",x"6f533d",x"6f553e",x"6b523c",x"6a503a",x"624b36",x"654e39",x"66503c",x"604c3b",x"5b4838",x"574434",x"524233",x"574535",x"584636",x"5a483a",x"655243",x"645142",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181008",x"191109",x"191109",x"1d140b",x"1f150b",x"261a0f",x"271b10",x"281c10",x"2c1e12",x"312215",x"2d2013",x"352518",x"342517",x"2f2013",x"302114",x"312215",x"322315",x"2f2014",x"332415",x"302214",x"302114",x"302114",x"332316",x"322316",x"352516",x"322315",x"362718",x"362618",x"382718",x"392819",x"352517",x"362617",x"352517",x"312215",x"352517",x"332416",x"362617",x"39281a",x"352517",x"352517",x"372718",x"392819",x"382819",x"3c2b1c",x"382819",x"2e2013",x"362617",x"3b291a",x"322316",x"412e1e",x"171009",x"150e07",x"181008",x"181008",x"1d140b",x"1d140b",x"20150b",x"20160c",x"21170d",x"25190f",x"281c10",x"25190e",x"271b10",x"2a1d11",x"291c11",x"291d11",x"2a1d11",x"2d1f12",x"281c10",x"312316",x"2d1f12",x"302114",x"2c1e12",x"2e2013",x"302214",x"352618",x"342517",x"2f2113",x"332315",x"312215",x"342417",x"312215",x"2e2013",x"312214",x"332416",x"312215",x"312215",x"312215",x"332314",x"322315",x"3a291a",x"322315",x"362617",x"372718",x"2f2114",x"362618",x"322315",x"312215",x"352517",x"2e2013",x"362619",x"433120",x"523b27",x"150e07",x"2a1d11",x"2c1e12",x"2e2013",x"302215",x"302214",x"150e07",x"150e07",x"150e07",x"312215",x"312215",x"2f2114",x"2e2013",x"2e2013",x"342416",x"2d1f13",x"372718",x"362616",x"3a2819",x"3b2a1b",x"382718",x"3a2819",x"392819",x"352517",x"3a2819",x"3b291a",x"392819",x"382818",x"3a2819",x"372618",x"3c2a1b",x"392819",x"362617",x"3c2a1b",x"3a2819",x"3f2d1d",x"402e1e",x"3f2d1d",x"362616",x"402d1c",x"382718",x"382719",x"3b291a",x"3a291a",x"3d2b1b",x"3a291a",x"3b291a",x"402d1c",x"402d1d",x"3e2b1a",x"3f2c1b",x"412f1e",x"3e2b1b",x"3d2a1b",x"3d2b1b",x"382718",x"3d2b1b",x"3b2a1a",x"3b291a",x"392818",x"3a2819",x"372618",x"3f2c1c",x"382718",x"3a2819",x"3a2919",x"3a2819",x"3d2b1c",x"3b2a1b",x"3a291a",x"352415",x"3f2c1c",x"3a2819",x"372618",x"352517",x"352517",x"332415",x"2f2114",x"312215",x"322215",x"3a281a",x"332314",x"312114",x"312114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"321c0d",x"3c2311",x"26150a",x"28160a",x"28160a",x"271509",x"211309",x"301b0c",x"321c0c",x"301b0c",x"321b0d",x"321c0c",x"341d0d",x"331c0d",x"321c0c",x"2c190b",x"2a180b",x"301c0c",x"341d0d",x"301b0b",x"301a0c",x"311b0c",x"331d0c",x"39200f",x"351e0d",x"361f0e",x"371f0e",x"331d0d",x"311b0c",x"321b0c",x"301a0c",x"331d0d",x"381f0e",x"311c0c",x"341d0d",x"371f0d",x"361e0d",x"311c0c",x"371f0e",x"361f0d",x"361e0e",x"351e0d",x"38200e",x"361f0e",x"371f0f",x"3c220f",x"371f0e",x"361f0e",x"37200e",x"321d0d",x"371f0e",x"331d0d",x"351e0e",x"38200f",x"36200e",x"341e0d",x"361f0e",x"38200e",x"371f0e",x"381f0f",x"341d0d",x"2f1b0c",x"361f0e",x"28180b",x"1a130c",x"18110a",x"19110a",x"180f08",x"180f08",x"191008",x"180f08",x"191008",x"191008",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1208",x"1d1208",x"1e1208",x"1d1208",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"1f1309",x"1f1309",x"1f1209",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1f1309",x"1e1208",x"1d1108",x"1d1108",x"1b1008",x"1a1007",x"1b1008",x"1a1008",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"1d1208",x"25150a",x"422613",x"150e07",x"150e07",x"150e07",x"321c0d",x"191008",x"261509",x"150e07",x"150e07",x"150e07",x"2f1a0b",x"180f08",x"150e07",x"24180f",x"150e07",x"150e07",x"2f1a0b",x"2f1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"876d55",x"896f58",x"5f5143",x"5e4f40",x"5b4a3b",x"5e4a38",x"5a4634",x"5b4533",x"634d38",x"654c38",x"69513b",x"664e3a",x"69503a",x"674e39",x"6a5039",x"6c523d",x"735840",x"715741",x"735a45",x"6f5743",x"745b46",x"725b47",x"6d5440",x"775d45",x"735943",x"785a40",x"76583d",x"735741",x"73573f",x"755a42",x"765a42",x"72563f",x"6f5640",x"755b42",x"6e5640",x"7b6347",x"7b6046",x"795d45",x"7a5d44",x"7a5c42",x"795d45",x"735840",x"775d45",x"7a5e46",x"7a5c43",x"6c523d",x"755840",x"765941",x"795d43",x"775d43",x"745840",x"715841",x"765d46",x"7d6149",x"745943",x"71573f",x"755a42",x"735943",x"765a43",x"735740",x"765b43",x"775a41",x"745941",x"755941",x"705640",x"705842",x"735c43",x"705b43",x"795f45",x"775d44",x"70563f",x"6b513c",x"6a533d",x"6d543f",x"6b533f",x"6c5642",x"65503e",x"5f4b3a",x"5e4a38",x"5b4737",x"5f4b38",x"5d4c3c",x"63503f",x"655342",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191109",x"191109",x"1e150b",x"191109",x"1e160c",x"20160d",x"23180e",x"251a0f",x"1e150b",x"1f150c",x"23180e",x"22170d",x"24190f",x"24190e",x"21160d",x"20160c",x"20160c",x"24190e",x"21170d",x"1d140b",x"1f150b",x"20160c",x"24190f",x"23180e",x"261a0f",x"261a0f",x"291c11",x"23180e",x"261a0f",x"251a0f",x"24190f",x"261a0f",x"21160d",x"291c10",x"24190e",x"241a0f",x"241a0f",x"291d12",x"281c11",x"251a0f",x"261a10",x"281c11",x"291d11",x"2f2115",x"271b10",x"3a2a1a",x"150e07",x"150e07",x"150e07",x"191109",x"191109",x"150e07",x"181008",x"191108",x"191109",x"191109",x"1e150b",x"191109",x"191109",x"191109",x"1e150b",x"1e140b",x"1e150c",x"1e140b",x"191109",x"1e140b",x"1e150b",x"1e150c",x"1e160c",x"20160d",x"1f160c",x"22170d",x"21170d",x"22180e",x"1e140b",x"241a0f",x"21170d",x"1e150b",x"23180e",x"20160c",x"23180d",x"24190e",x"24190e",x"20160c",x"23170d",x"22170d",x"2a1e12",x"21160c",x"24190e",x"21170d",x"23180e",x"20160c",x"24190e",x"261a0f",x"24190e",x"21160c",x"271b10",x"342517",x"4f3a25",x"191109",x"2a1f13",x"2f2215",x"2c1f13",x"2f2115",x"302215",x"150e07",x"150e07",x"150e07",x"332417",x"362618",x"322316",x"312214",x"332316",x"392819",x"392819",x"382718",x"332315",x"382717",x"362819",x"392819",x"3f2d1d",x"3a291a",x"3f2d1c",x"3a291a",x"3f2e1e",x"412e1e",x"3f2e1d",x"412e1d",x"3c2b1b",x"3e2c1c",x"3f2e1e",x"3c2d1d",x"3d2f1f",x"443222",x"412f1e",x"412f1e",x"443120",x"443120",x"3f2d1d",x"402f1f",x"402e1e",x"44311f",x"3f2c1c",x"412e1d",x"402d1c",x"422f1f",x"453220",x"3e2c1c",x"392717",x"3c2a19",x"3e2d1d",x"3e2c1c",x"43311f",x"3c2a1b",x"402e1d",x"3e2b1b",x"402e1e",x"402d1d",x"3d2c1c",x"3f2d1c",x"3e2c1c",x"3f2d1c",x"3c2b1b",x"3d2f1f",x"413221",x"463423",x"443220",x"3f2d1d",x"3f2d1e",x"443120",x"402e1d",x"423020",x"3c2b1c",x"392819",x"3d2b1b",x"322315",x"372718",x"332416",x"362718",x"372718",x"322314",x"322215",x"322215",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"361e0d",x"191008",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"1a120b",x"181009",x"191109",x"170f07",x"180f07",x"180f08",x"180f08",x"191008",x"180f08",x"180f08",x"190f08",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1b1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1d1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1b1008",x"191008",x"191008",x"191008",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"201508",x"251709",x"1d1208",x"25150a",x"452813",x"150e07",x"150e07",x"150e07",x"2e1a0b",x"1f1309",x"27170a",x"191008",x"150e07",x"150e07",x"351e0e",x"241509",x"150e07",x"261910",x"150e07",x"150e07",x"301b0c",x"301b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"8a6e55",x"886c54",x"57493b",x"554638",x"584738",x"544232",x"5d4836",x"5f4935",x"624d3a",x"644e39",x"644e39",x"69513b",x"6c533f",x"6a5440",x"705742",x"715a45",x"735a43",x"745b44",x"715843",x"765b46",x"715842",x"705845",x"745a45",x"745a44",x"735942",x"755940",x"6f543b",x"71563f",x"775a43",x"705640",x"735841",x"725740",x"755a41",x"755941",x"775a41",x"71563f",x"775c43",x"71553f",x"715740",x"775b41",x"67513c",x"755b43",x"775d44",x"755b44",x"775b43",x"7a5e45",x"775941",x"785e45",x"7a5d43",x"7a5f44",x"785c43",x"7c5f48",x"765b44",x"705540",x"725842",x"755a43",x"6f5640",x"745942",x"735841",x"71563f",x"775b42",x"72563f",x"725841",x"74573f",x"765c44",x"735943",x"725942",x"725740",x"725840",x"6e523b",x"725741",x"6b523c",x"6d5741",x"6a543f",x"6b5440",x"6a523f",x"6a533e",x"65503e",x"644f3d",x"5e4c3b",x"604c3d",x"5d4d3e",x"675545",x"675545",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181109",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1f13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"291d11",x"483422",x"181009",x"291c10",x"2e2114",x"291e12",x"191109",x"160f08",x"150e07",x"2d1a0b",x"150e07",x"352517",x"332416",x"332416",x"352618",x"39291b",x"362617",x"362718",x"3a281a",x"3c2a1b",x"3d2b1c",x"382718",x"3a2819",x"3b2919",x"3b2a1a",x"3d2b1b",x"382718",x"3a2919",x"3f2d1d",x"3d2b1b",x"3d2b1b",x"382719",x"412e1d",x"402e1d",x"412f1e",x"3e2b1c",x"3e2d1d",x"3b291a",x"42301f",x"453220",x"3d2f1e",x"3d2d1d",x"3f2d1d",x"3d2c1c",x"422f1f",x"412f1e",x"3e2c1d",x"453221",x"412e1e",x"42301f",x"45311f",x"44311f",x"402e1d",x"3e2c1c",x"432f1e",x"412e1d",x"3d2b1b",x"3f2c1c",x"3b291a",x"3d2b1b",x"42301f",x"3d2b1b",x"3b2a1a",x"3a281a",x"3a291a",x"3f2d1c",x"3a291a",x"3c2a1b",x"422f1f",x"3b291a",x"43301f",x"422f1f",x"3d2e1e",x"3e2d1d",x"3f2d1d",x"3c2b1b",x"3d2b1c",x"3b2a1a",x"372719",x"3c2c1c",x"382719",x"362618",x"392819",x"362618",x"322316",x"322316",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"301b0c",x"321c0c",x"3a210f",x"291609",x"150e07",x"180f08",x"170f07",x"1b1008",x"1c1108",x"1d1108",x"201208",x"1c1108",x"1c1108",x"170f07",x"170f07",x"1b1108",x"1c1108",x"1a1008",x"1d1208",x"1d1208",x"1e1208",x"1a1008",x"1a1008",x"1e1208",x"1d1108",x"1a1008",x"1b1008",x"180f08",x"1c1108",x"180f07",x"150e07",x"170f08",x"1a1008",x"201309",x"211309",x"1b1108",x"1a1008",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"170e08",x"1c1108",x"170f07",x"1b1108",x"170f07",x"170f07",x"1a1008",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"1c1108",x"150e07",x"191008",x"160f07",x"3b220f",x"19120b",x"181009",x"27160a",x"28170a",x"2a180a",x"2b180a",x"3d2311",x"311b0c",x"2b180b",x"2a180b",x"2c190a",x"2f1a0b",x"2c190b",x"2f1a0b",x"2e190b",x"2d190b",x"2c180b",x"321b0c",x"2d190b",x"29160a",x"2b180a",x"2c190b",x"301b0c",x"331c0c",x"321c0c",x"311b0c",x"301a0b",x"341d0d",x"321c0c",x"361f0e",x"331d0d",x"351f0e",x"341e0e",x"361f0e",x"331e0d",x"341e0d",x"2d190b",x"2e1a0b",x"321d0d",x"321d0e",x"2f1c0c",x"311c0c",x"351e0e",x"301c0c",x"321c0d",x"2f1c0d",x"311d0d",x"311c0d",x"331e0e",x"361f0f",x"36200e",x"351f0e",x"2f1b0c",x"331d0c",x"321c0c",x"2e1a0b",x"311c0c",x"331d0d",x"361f0e",x"351f0e",x"351e0e",x"341d0d",x"361f0e",x"361f0e",x"361f0f",x"341e0e",x"351f0e",x"341e0e",x"382110",x"341e0e",x"321d0d",x"361f0e",x"321d0d",x"2d190c",x"2d1a0c",x"321c0c",x"331c0c",x"341d0e",x"3d2310",x"412612",x"27180c",x"412412",x"150e07",x"150e07",x"150e07",x"2a170a",x"1d1108",x"29170a",x"180f08",x"150e07",x"150e07",x"311c0d",x"1d1108",x"150e07",x"261910",x"150e07",x"150e07",x"321c0c",x"321c0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"8b6d55",x"896e55",x"57493c",x"554436",x"564637",x"5d4939",x"5f4938",x"654f3c",x"654d3a",x"6a513c",x"6a533f",x"6b5440",x"725a46",x"715b46",x"735b47",x"765b47",x"715844",x"755d48",x"745b47",x"715843",x"725843",x"785e46",x"735842",x"765c45",x"755942",x"755a43",x"745841",x"765a42",x"6e553f",x"7c6148",x"775b43",x"73583f",x"795f47",x"7b6046",x"795e45",x"785c43",x"785c43",x"755940",x"73573f",x"7a5d44",x"785c43",x"795d42",x"7b5f46",x"785d44",x"7b6046",x"775a41",x"785b43",x"795c43",x"7a5d44",x"795d45",x"7d6147",x"73573f",x"7a5d45",x"775d44",x"745942",x"745a43",x"735842",x"725840",x"795e46",x"765a43",x"755b43",x"795f48",x"755841",x"745842",x"755b44",x"755b44",x"745a42",x"715640",x"6b523d",x"725741",x"6e5540",x"6e5640",x"6f553f",x"6d543e",x"6f5742",x"6b543e",x"6a533f",x"675342",x"665342",x"655140",x"614f41",x"625143",x"645343",x"655444",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2717",x"54453a",x"47372c",x"483b30",x"47382d",x"40342a",x"463428",x"463529",x"463427",x"45362a",x"4e3a2d",x"563925",x"4f3c2f",x"514034",x"4b392d",x"594436",x"543f31",x"584739",x"5c4334",x"5b4436",x"584132",x"584537",x"543f31",x"564336",x"534134",x"4b372a",x"503b2d",x"49372b",x"543f31",x"4b382b",x"503f32",x"4e382a",x"4f3d31",x"533d2f",x"594131",x"5a4030",x"5a402e",x"5a3c2a",x"553d2d",x"523e2f",x"563d2d",x"493528",x"483629",x"543c2c",x"533a2a",x"503a2b",x"5a402f",x"4f3b2d",x"48382d",x"483529",x"533c2f",x"46372c",x"4b3a2e",x"513a2b",x"573f2f",x"443125",x"483326",x"45352a",x"46382d",x"4a392d",x"523b2d",x"553d2f",x"523e30",x"4b3a2f",x"493a2e",x"473529",x"493528",x"4d3a2e",x"4e392c",x"4d3829",x"563f2f",x"563d2d",x"4f392b",x"513929",x"453124",x"553a28",x"4d3a2e",x"48382d",x"4a382d",x"4e3a2d",x"47372b",x"4f3b2e",x"4c382a",x"553f31",x"4e3b2e",x"4d3b2e",x"4d3a2d",x"4e3a2c",x"503c2e",x"5d4433",x"533f32",x"593f2f",x"563f30",x"593e2d",x"553c2b",x"483427",x"533c2d",x"4a3628",x"4b3627",x"413329",x"3e3228",x"43342a",x"513e31",x"46392e",x"473a30",x"4f3e32",x"4a3e34",x"533118",x"150e07",x"150e07",x"150e07",x"150e07",x"442711",x"191109",x"302215",x"302215",x"352517",x"332416",x"382718",x"342416",x"362618",x"39291a",x"3d2b1c",x"3c2a1b",x"3b2a1a",x"3c2a1b",x"3a2919",x"3c2a1a",x"412f1e",x"3f2d1c",x"422f1f",x"3d2b1c",x"402e1e",x"402d1c",x"402e1d",x"402e1e",x"433120",x"3f2d1d",x"3d2b1c",x"3e2c1c",x"412e1e",x"412e1d",x"412f1f",x"422f1e",x"3d2c1c",x"443120",x"443120",x"453220",x"43301f",x"3f2c1c",x"45311f",x"402d1d",x"453120",x"412f1f",x"422f1e",x"3f2d1c",x"43301f",x"3e2c1c",x"402d1c",x"3e2b1b",x"43301f",x"412e1e",x"402e1e",x"422f1e",x"473422",x"402d1c",x"3b2a1a",x"422f1f",x"433120",x"412f1e",x"3d2b1c",x"3c2a1b",x"3f2c1d",x"3d2b1b",x"43301f",x"3f2d1d",x"3c2b1b",x"3d2c1d",x"3a2a1a",x"3d2b1c",x"3e2c1c",x"372718",x"3e2b1b",x"362517",x"342517",x"332417",x"362618",x"312315",x"312315",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"160f07",x"2d190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"231409",x"25160a",x"25160a",x"241509",x"25150a",x"25160a",x"26160a",x"27160a",x"26160a",x"26160a",x"27170a",x"28170b",x"27170a",x"27170a",x"27160a",x"251509",x"27160a",x"28170a",x"28170b",x"2b190b",x"29170a",x"27170a",x"28170a",x"27160a",x"28170a",x"251509",x"241409",x"27160a",x"27160a",x"27160a",x"251509",x"27160a",x"26160a",x"27170a",x"27170a",x"28170b",x"26160a",x"28170b",x"28180b",x"28170b",x"27170a",x"29180b",x"2a190b",x"28170a",x"28170a",x"28170a",x"28170b",x"28170b",x"27170a",x"26160a",x"26160a",x"241509",x"26160a",x"28170a",x"26160a",x"261609",x"231409",x"261609",x"211308",x"241509",x"241409",x"25150a",x"26160a",x"26160a",x"251509",x"251509",x"241409",x"241509",x"241509",x"26160a",x"26160a",x"211409",x"1f1309",x"1f140b",x"1d130a",x"1e140d",x"21170f",x"20160c",x"27170c",x"3d2210",x"150e07",x"150e07",x"150e07",x"2a170a",x"1a1008",x"251509",x"1b1108",x"150e07",x"150e07",x"2e190b",x"221409",x"150e07",x"25190f",x"150e07",x"150e07",x"341e0d",x"341e0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"836851",x"876c54",x"534539",x"504234",x"584838",x"5e4b3c",x"65513f",x"67513e",x"6d5742",x"715842",x"6f5945",x"6d5844",x"765f4b",x"735b47",x"79634f",x"78614d",x"745d4a",x"735b46",x"745c48",x"715945",x"785c47",x"715742",x"705741",x"6d5440",x"6e5540",x"755a45",x"715740",x"775c44",x"775c44",x"735943",x"765b44",x"775b44",x"765c46",x"795e46",x"7a6047",x"7d6149",x"775c45",x"745b46",x"7c624a",x"7a5e46",x"7b6048",x"7d6148",x"715945",x"7d6047",x"7e6149",x"7c624a",x"7e644e",x"7b624b",x"7a604a",x"795e47",x"785c45",x"7a5d45",x"775a43",x"755942",x"6e553f",x"6c513d",x"70543e",x"745a43",x"765b43",x"765b43",x"755a43",x"765b43",x"765c43",x"765b45",x"755b43",x"775c44",x"765b44",x"785c43",x"775b42",x"735840",x"745941",x"735842",x"775d46",x"755c46",x"6f5640",x"6d5742",x"6b5541",x"725d4a",x"6d5a49",x"645241",x"604e40",x"5c4f42",x"695747",x"6d5a49",x"6d5a49",x"000000",x"000000",x"000000",x"472d1b",x"472d1b",x"4c3c31",x"493a2e",x"4f3e31",x"47382c",x"513c2e",x"4d3626",x"4e3524",x"523725",x"4f3727",x"483324",x"4e3727",x"553d2c",x"533a2a",x"523b2c",x"4d392b",x"593c2a",x"5a3f2d",x"5a4131",x"593e2d",x"5e4534",x"563b28",x"543c2c",x"573c2b",x"543e30",x"584232",x"5a3f2f",x"5c4333",x"573d2b",x"553d2d",x"533a2a",x"543e30",x"493325",x"573e2d",x"553b2b",x"5f422d",x"583a26",x"563723",x"5c3d27",x"583b26",x"4d3424",x"4e3523",x"533b29",x"543a29",x"4c3626",x"573c2a",x"553b29",x"5a3b28",x"553826",x"573b29",x"563b28",x"5c402e",x"5d412d",x"674732",x"503b2c",x"4f3c2d",x"4c382b",x"4b392d",x"4d392c",x"533a2a",x"573b29",x"513929",x"5b3e2b",x"523b2c",x"4e3a2c",x"543d2f",x"503828",x"4d3525",x"513625",x"4e3524",x"4f3624",x"543b2b",x"4d3628",x"593b28",x"543928",x"513727",x"513829",x"4d3728",x"483325",x"4b3323",x"4e382a",x"523928",x"553f30",x"543c2c",x"533d2f",x"533a2b",x"563e2e",x"573f30",x"593e2d",x"5a3f2c",x"563b2a",x"513b2c",x"5a3f2e",x"503a2d",x"4b3629",x"4c392b",x"4b3425",x"4c3222",x"4b3323",x"4e3829",x"3d2d22",x"473225",x"46352a",x"44362a",x"473426",x"4f3b2b",x"534033",x"4e2d15",x"150e07",x"150e07",x"150e07",x"150e07",x"472912",x"191109",x"332417",x"302215",x"372819",x"362617",x"342416",x"3c2b1b",x"362618",x"3a2819",x"372617",x"3a2919",x"3a2919",x"352516",x"352416",x"362617",x"3b291a",x"3a2819",x"3f2d1c",x"3e2c1c",x"3d2b1b",x"3e2c1c",x"3e2c1c",x"3e2c1c",x"402e1e",x"3d2c1c",x"422f1f",x"402e1d",x"422f1f",x"443120",x"3f2c1c",x"463321",x"483423",x"412e1e",x"43301f",x"42301f",x"433120",x"453220",x"412e1d",x"43301e",x"44301f",x"432f1d",x"412e1d",x"432f1e",x"44301e",x"3e2b1b",x"382718",x"3b2919",x"3e2b1c",x"3d2b1b",x"402e1d",x"3e2c1c",x"3e2c1c",x"3e2c1c",x"44301f",x"3c2a1b",x"3e2c1d",x"453220",x"412e1e",x"402e1d",x"422f1f",x"433020",x"412e1e",x"443120",x"412f1f",x"412e1e",x"3b2a1b",x"3f2d1d",x"3e2d1d",x"3e2c1c",x"382718",x"382718",x"342416",x"322315",x"322215",x"362517",x"362517",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c1108",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"27160a",x"26160a",x"24150a",x"25170a",x"27170b",x"28180b",x"27170a",x"27160a",x"26160a",x"27170a",x"27170a",x"27170a",x"26160a",x"241509",x"231409",x"25150a",x"27170a",x"27170a",x"27170a",x"26160a",x"27170a",x"25150a",x"27170a",x"26160a",x"25160a",x"251509",x"25160a",x"26160a",x"25160a",x"231409",x"241509",x"25150a",x"26160a",x"241509",x"26160a",x"25150a",x"26160a",x"28180b",x"28180b",x"28180b",x"28180b",x"28180b",x"28170b",x"26160a",x"25150a",x"25160a",x"25150a",x"26160a",x"27160a",x"29180b",x"2a190c",x"2a190c",x"2b1a0c",x"27160a",x"28180b",x"26160a",x"251509",x"231409",x"231409",x"25160a",x"25150a",x"25150a",x"25150a",x"26160a",x"231409",x"26160a",x"26160a",x"27160a",x"26160a",x"25150a",x"25160a",x"211409",x"21140c",x"22160d",x"22170f",x"241b13",x"231a12",x"241b14",x"27180d",x"3b200e",x"150e07",x"150e07",x"150e07",x"2b180a",x"1b1108",x"261609",x"1a1008",x"150e07",x"150e07",x"301c0d",x"1c1108",x"150e07",x"25180e",x"150e07",x"150e07",x"341d0d",x"341d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"7c644f",x"7b634d",x"564a40",x"574b3f",x"594b3f",x"5c4b3b",x"665242",x"6f5945",x"765d4a",x"775f4b",x"705945",x"725b49",x"745c49",x"77604b",x"785e4a",x"7b634e",x"79614e",x"7b614c",x"775e4a",x"765c47",x"745a44",x"7b614a",x"7b624b",x"80654c",x"7d634c",x"7c6149",x"7b614b",x"7a5f48",x"7b614b",x"7c614b",x"785d46",x"795d47",x"785e47",x"7c6149",x"795d47",x"755c47",x"715a46",x"745b46",x"765e4a",x"7d624a",x"7c614a",x"7d634c",x"7e644f",x"7d634d",x"79614c",x"7e644e",x"806751",x"826650",x"7c624b",x"7e634c",x"795e47",x"795d46",x"795d44",x"765941",x"7c5f46",x"80634b",x"795e46",x"785c44",x"816248",x"80634a",x"7c5f47",x"7d6149",x"7a5e45",x"7b5e45",x"785c44",x"795f49",x"785c46",x"765b43",x"6b513c",x"6e533e",x"725740",x"795d45",x"765d48",x"785e47",x"735b46",x"735943",x"6f5946",x"725d4b",x"6f5b4a",x"6d5a4a",x"625447",x"5e5144",x"836852",x"836952",x"836952",x"000000",x"000000",x"000000",x"452b1a",x"452b1a",x"534134",x"503a2b",x"543b2c",x"563f2f",x"4d3729",x"4d3728",x"4b3324",x"553827",x"593e2b",x"583e2d",x"573b28",x"4c3424",x"4c3223",x"573d2d",x"553928",x"5c3f2d",x"5a402f",x"5a3e2a",x"593a24",x"5d3f2a",x"583b28",x"513727",x"513625",x"543725",x"543a28",x"573b28",x"523725",x"4c3626",x"513929",x"4d3627",x"533826",x"4f3522",x"563827",x"60402b",x"61412a",x"603e27",x"5f3f28",x"5d3f2a",x"573d2a",x"593e2a",x"513929",x"4f3727",x"513524",x"4d3322",x"563925",x"61412c",x"593a26",x"5b3b26",x"5c3f29",x"573b27",x"5d412b",x"583c29",x"61422d",x"563d2b",x"503c2c",x"503b2d",x"523c2c",x"5b4231",x"573d2b",x"5a3e2c",x"5c3f2e",x"593f2e",x"543c2d",x"60432e",x"5d412e",x"553d2b",x"593c29",x"61412b",x"563b28",x"543c2a",x"4d3424",x"563b29",x"503626",x"543825",x"583d2b",x"543a29",x"593d2b",x"4f3627",x"503524",x"513828",x"4f3728",x"513727",x"563b2a",x"5b3e2c",x"583c2b",x"5b3f2c",x"5d3f2b",x"543827",x"543b2b",x"5e3c27",x"563a29",x"4c3324",x"513728",x"4e3728",x"4f3727",x"543a29",x"4b3324",x"453021",x"473223",x"482d1b",x"402a1b",x"3d291d",x"3b291d",x"453326",x"49372a",x"44362b",x"4d2c15",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2c14",x"150e07",x"312215",x"2f2114",x"352517",x"332316",x"342517",x"362618",x"3b291a",x"3c2a1b",x"392819",x"412e1d",x"3e2b1b",x"3e2b1b",x"412f1f",x"3d2b1b",x"44301e",x"3e2c1c",x"3c2b1c",x"3f2c1c",x"3f2d1c",x"3e2b1b",x"3e2c1c",x"3e2c1c",x"3c2b1b",x"3f2c1c",x"3c2a1a",x"3a2819",x"3c2a1b",x"412e1d",x"432f1e",x"43301f",x"402e1d",x"3e2c1c",x"44301f",x"3b291a",x"3e2c1c",x"3b2a1a",x"422f1e",x"43301f",x"412e1e",x"422e1d",x"402d1c",x"473220",x"432f1d",x"422f1d",x"412f1f",x"3f2c1c",x"3f2c1c",x"473221",x"453220",x"45311f",x"3f2d1c",x"3c2a1b",x"44301f",x"3d2b1b",x"3e2c1c",x"382718",x"3a291a",x"332316",x"382819",x"3a2819",x"3b291a",x"3c2a1b",x"402e1d",x"3d2b1c",x"382718",x"382718",x"3a2919",x"382718",x"3d2b1c",x"382819",x"342416",x"342416",x"332315",x"332316",x"332316",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"321d0d",x"180f08",x"181008",x"150e07",x"25170b",x"24160a",x"211409",x"1f1309",x"221409",x"1e1208",x"1e1208",x"1e1208",x"1b1108",x"1e1209",x"23150a",x"22150a",x"26170b",x"1c1108",x"191008",x"1d1209",x"211409",x"1f1309",x"1e1209",x"1f1309",x"1f1309",x"1b1108",x"1d1208",x"1c1108",x"1d1209",x"1f1309",x"180f08",x"1e1209",x"1e1209",x"191008",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"211409",x"180f07",x"211409",x"1d1108",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"1d1208",x"180f07",x"1a1008",x"160e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f08",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1d1208",x"1f1209",x"1f1309",x"1d1208",x"1f1208",x"1f1309",x"1f1309",x"1f1309",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1f1309",x"1d1208",x"1d1208",x"1f1209",x"1d1209",x"1e1209",x"1f1309",x"1f1309",x"1e1309",x"201409",x"201409",x"1f1309",x"1e1209",x"1d1208",x"1d1208",x"1d1108",x"1d1208",x"1d1108",x"1e1209",x"201409",x"1f1409",x"201309",x"1f1309",x"1f1309",x"1f1309",x"1d1208",x"1e1208",x"1e1209",x"1d1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"191008",x"180f08",x"180f08",x"170f07",x"180f08",x"170f07",x"170f07",x"170f07",x"170f07",x"241911",x"251b13",x"251c14",x"1d1208",x"27180c",x"3e230f",x"150e07",x"150e07",x"150e07",x"311d0d",x"1b1108",x"2d1a0b",x"1d1208",x"150e07",x"150e07",x"331d0d",x"1f1208",x"150e07",x"27180d",x"150e07",x"150e07",x"2f1b0b",x"2f1b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"765e4a",x"6b4b31",x"5e432c",x"593f2a",x"62472f",x"5a412b",x"674c34",x"6b5036",x"6b4f36",x"705238",x"715338",x"6f5138",x"6f5033",x"6f5035",x"674a2f",x"7a5a3f",x"735439",x"755539",x"76573a",x"77583a",x"725337",x"715136",x"745438",x"74563a",x"78583b",x"79593c",x"6e4f34",x"6d4e34",x"5f442c",x"6e4f35",x"75553a",x"79583c",x"7c5c3f",x"79583c",x"79583b",x"7c5c3d",x"805e41",x"7b5939",x"7a5739",x"705032",x"745437",x"846042",x"7e5b3e",x"785638",x"7b593b",x"7b593a",x"785738",x"7a573b",x"765539",x"7e5d3f",x"7b5b3e",x"745438",x"6f4f35",x"6f5035",x"715036",x"735438",x"77583a",x"7e5c40",x"7d5c40",x"7a593e",x"77573b",x"7f5e41",x"7c5c3f",x"725336",x"7c5a3b",x"745538",x"856345",x"7b5b3f",x"785a3d",x"73553a",x"715338",x"715339",x"6f5037",x"6e5138",x"6e5137",x"6a4d35",x"664b33",x"5e432c",x"533b26",x"60432c",x"664a30",x"705137",x"735338",x"77563b",x"000000",x"000000",x"000000",x"000000",x"442b1a",x"442b1a",x"544337",x"453326",x"4c392d",x"4f3829",x"4a3426",x"4d3120",x"4b301f",x"4e3321",x"533523",x"583a25",x"563b29",x"513626",x"4d3728",x"513929",x"543725",x"543826",x"553624",x"573824",x"573927",x"553928",x"523928",x"523929",x"4f3626",x"563927",x"5a3f2d",x"5c3d28",x"573b28",x"543928",x"4a3325",x"4c3323",x"473020",x"523726",x"573a26",x"593c28",x"5f402b",x"603f28",x"5a3b24",x"583a25",x"4e3523",x"4a3321",x"473020",x"503522",x"573a25",x"5a3b26",x"5b3c28",x"533725",x"4d3120",x"4e3323",x"4b3122",x"493224",x"4d3528",x"4e3527",x"4c3729",x"573c2c",x"443329",x"4b3528",x"4d382b",x"573d2d",x"5a3d2b",x"5c3e2b",x"593d2c",x"5e422e",x"583d2b",x"60422f",x"634532",x"60422e",x"61412b",x"5e3e28",x"5a3d2a",x"5d3f2c",x"5e3c27",x"563a28",x"573b28",x"593b27",x"543725",x"593b26",x"563925",x"563a27",x"593b28",x"583b27",x"573b28",x"4e3524",x"523725",x"543825",x"583c29",x"5c3e2b",x"593a26",x"603f2a",x"60412c",x"583b28",x"563b2b",x"533825",x"4f3422",x"432c1b",x"3f2a1d",x"402a1b",x"3b2515",x"432b1c",x"453023",x"3e2a1c",x"432c1d",x"3f2c20",x"452f20",x"3a281c",x"463327",x"453326",x"4e2e15",x"150e07",x"150e07",x"150e07",x"150e07",x"472812",x"191109",x"322316",x"332417",x"3a2a1b",x"3c2b1c",x"372718",x"3c2a1b",x"372719",x"3c2a1b",x"412e1e",x"3a291b",x"412f1f",x"402f1e",x"3c2a1b",x"402d1d",x"44301f",x"3c2a1b",x"3e2c1c",x"3b2a1b",x"412e1e",x"412e1d",x"3d2b1b",x"412f1e",x"3e2c1c",x"372617",x"372617",x"3c2b1a",x"3c2a1b",x"3e2b1c",x"3f2c1c",x"412e1d",x"422f1d",x"3f2d1d",x"3f2d1c",x"43301f",x"493523",x"473322",x"402d1d",x"463221",x"422f1e",x"453220",x"453220",x"433120",x"4d3825",x"483422",x"422f1f",x"443120",x"402e1d",x"463121",x"43301f",x"44311f",x"453120",x"412e1d",x"3c2a1b",x"3d2b1c",x"43301f",x"332214",x"3b2919",x"372618",x"392819",x"392819",x"372718",x"3e2c1c",x"3d2b1b",x"3f2d1d",x"3e2c1c",x"3e2c1d",x"3e2d1d",x"3c2b1c",x"372718",x"3a291a",x"392819",x"332416",x"392819",x"39291a",x"39291a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1008",x"1f1208",x"513118",x"563319",x"543319",x"513117",x"5b3519",x"5a361a",x"5a371c",x"59351a",x"553118",x"452511",x"45240f",x"3a1d0b",x"351d0c",x"361d0d",x"341c0c",x"311a0b",x"361d0d",x"3a200e",x"31190a",x"321a0b",x"371d0d",x"3e2210",x"3b210f",x"3d220f",x"412410",x"3a210f",x"402511",x"422611",x"462913",x"412511",x"3d2310",x"432712",x"442712",x"402410",x"3c220f",x"3e220f",x"3f2411",x"3e220f",x"3a200e",x"3b210f",x"3d220f",x"3d2310",x"442712",x"432712",x"3c2210",x"3f2411",x"412511",x"412611",x"432712",x"3d2311",x"422612",x"432812",x"412611",x"3c230f",x"3c220f",x"3a210e",x"3d230f",x"3c220f",x"3b210e",x"3b200e",x"3c200d",x"4b2b14",x"4f2d14",x"4c2a14",x"1a1008",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"191008",x"191008",x"191008",x"191008",x"190f07",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1e1209",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1c1208",x"1c1108",x"1c1208",x"1c1108",x"1c1108",x"1d1208",x"1d1209",x"1d1208",x"1c1108",x"1a1008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"190f07",x"1a1008",x"1c1108",x"190f07",x"190f07",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"180f08",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"251b13",x"1d1209",x"1d1209",x"27180c",x"381e0d",x"150e07",x"150e07",x"150e07",x"38210f",x"1f1309",x"2f1b0d",x"150e07",x"150e07",x"150e07",x"28160a",x"191008",x"150e07",x"26180e",x"150e07",x"150e07",x"2c190b",x"2c190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"211309",x"211309",x"1f1208",x"26160a",x"28170a",x"381f0e",x"3a200d",x"381f0d",x"3c210e",x"3e220f",x"40230f",x"41240f",x"412410",x"472712",x"442611",x"462712",x"4b2b14",x"492913",x"442611",x"351d0d",x"2f1b0c",x"402510",x"3f230f",x"3a1f0d",x"3e220f",x"422511",x"3d210f",x"402310",x"462913",x"462813",x"442712",x"442711",x"462813",x"442712",x"442712",x"3f2310",x"442612",x"452812",x"4c2c15",x"462813",x"381f0e",x"412612",x"4f2f17",x"4a2c15",x"4a2c15",x"482a15",x"482b15",x"452812",x"422611",x"412511",x"492a14",x"4d2e16",x"502f17",x"4b2c15",x"4b2c15",x"492a13",x"4b2c15",x"523017",x"4c2d15",x"472812",x"452712",x"472912",x"462712",x"402511",x"4a2a14",x"4a2b15",x"4c2c15",x"4c2c15",x"492a14",x"38200f",x"331d0d",x"2f1b0c",x"2d1a0c",x"41372e",x"150e07",x"6a4d35",x"664b33",x"5e432c",x"533b26",x"60432c",x"664a30",x"705137",x"735338",x"77563b",x"000000",x"000000",x"000000",x"000000",x"442b1a",x"442b1a",x"493a2f",x"4a3426",x"4a3426",x"503626",x"493123",x"483224",x"4d3424",x"473123",x"523623",x"583a26",x"563826",x"5a3924",x"533624",x"4e3323",x"4f3424",x"5b3a26",x"513422",x"513523",x"573a28",x"553828",x"533827",x"583e2d",x"4e3626",x"543a29",x"563b29",x"573927",x"543825",x"553a28",x"4e3625",x"543927",x"4e3424",x"4b301e",x"503725",x"543a28",x"4c301e",x"573926",x"553a29",x"573924",x"543726",x"553825",x"4a3222",x"533826",x"5e3d28",x"583a28",x"523828",x"5d3e2a",x"63422c",x"62432d",x"5a3b27",x"5e3f2b",x"543725",x"553929",x"60412d",x"5e3e29",x"61442f",x"634530",x"644530",x"654631",x"5e4432",x"5e4130",x"5a3f2d",x"5c402d",x"5c3f2b",x"5a402d",x"60402c",x"66442c",x"62412a",x"62422d",x"66442c",x"63412b",x"5d3e29",x"5a3b26",x"5c3c25",x"593a25",x"5b3a24",x"543928",x"5b3a23",x"573924",x"543825",x"613f28",x"513624",x"4f3421",x"523724",x"543724",x"563a27",x"5a3b26",x"583824",x"5d3b24",x"553621",x"553824",x"553723",x"4b311f",x"4c321f",x"482f20",x"472f1e",x"4a2e1d",x"472e1e",x"4a301e",x"472d1a",x"492d1a",x"372011",x"342216",x"392619",x"3c271a",x"412d20",x"402d21",x"4f2e17",x"150e07",x"150e07",x"150e07",x"150e07",x"442511",x"191109",x"2e2014",x"2d1f13",x"352618",x"38281a",x"3a291a",x"3c2b1c",x"3d2c1c",x"3f2d1d",x"423020",x"402e1e",x"3c2b1c",x"3c2b1c",x"433221",x"3f2d1e",x"3f2e1e",x"3f2d1e",x"3e2c1c",x"3d2b1b",x"3d2b1b",x"3b2919",x"392819",x"453220",x"412e1d",x"3f2d1d",x"402d1d",x"3d2c1d",x"3d2b1b",x"3a2819",x"352516",x"3d2b1b",x"453220",x"43311f",x"422f1f",x"422f1e",x"483422",x"4a3624",x"493523",x"453221",x"493523",x"4b3724",x"493524",x"4b3624",x"4b3725",x"4c3725",x"4e3a27",x"4c3725",x"483423",x"4b3725",x"44301f",x"412e1d",x"3f2d1c",x"3f2d1b",x"3d2b1b",x"422f1e",x"44311f",x"44311f",x"43301f",x"42301f",x"3d2b1b",x"3a2819",x"362617",x"3b291a",x"433120",x"402e1e",x"3a291a",x"392819",x"3f2d1d",x"3a2a1b",x"3a291a",x"3d2c1d",x"3d2c1c",x"3b2a1c",x"3f2d1e",x"3a2a1c",x"3a2a1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"3b210f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"28160a",x"170f07",x"1b1008",x"1f1208",x"1d1108",x"1f1208",x"180f07",x"160e07",x"190f07",x"170f07",x"170f07",x"170f07",x"180f07",x"170f07",x"180f07",x"1d1108",x"191008",x"1b1108",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1d1108",x"1b1008",x"1e1208",x"1b1108",x"1a1008",x"1f1308",x"1d1108",x"1b1008",x"231509",x"1a1008",x"1a1008",x"191008",x"1b1108",x"191008",x"180f07",x"180f07",x"1f1209",x"1f1309",x"1d1208",x"211409",x"180f07",x"1b1108",x"211409",x"201309",x"1c1108",x"201309",x"201309",x"1e1208",x"211409",x"1e1209",x"1f1309",x"211309",x"24150a",x"1c1108",x"22150a",x"22150a",x"24150a",x"211409",x"1d1208",x"201409",x"1b1108",x"1d1208",x"191008",x"180f08",x"1e1209",x"1f1309",x"1b1108",x"29180b",x"2f1c0d",x"36200f",x"3b2310",x"311c0d",x"2a180b",x"201309",x"201309",x"000000",x"1d1109",x"1d1109",x"26170c",x"3d220f",x"150e07",x"150e07",x"150e07",x"361f0f",x"180f08",x"2c1a0c",x"150e07",x"150e07",x"150e07",x"351f0e",x"150e07",x"150e07",x"2c1e15",x"150e07",x"150e07",x"2a170a",x"2a170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"27170a",x"26160a",x"29170a",x"331c0d",x"341d0d",x"2e190b",x"2b180a",x"2e1a0b",x"321c0c",x"351e0d",x"371f0e",x"38200e",x"341d0d",x"371f0e",x"351f0e",x"39210f",x"39210f",x"3a2110",x"331d0d",x"2e1a0c",x"361f0e",x"301b0c",x"331d0d",x"2f1a0c",x"341e0d",x"371f0e",x"331e0d",x"311d0d",x"3a2411",x"382210",x"321d0d",x"3d2411",x"37200f",x"37200f",x"38200f",x"2f1c0d",x"3a2110",x"3a2210",x"39210f",x"3c2511",x"37200e",x"392311",x"3c2512",x"3f2612",x"3c2512",x"3c2311",x"392612",x"382411",x"3b2411",x"38200e",x"3a210f",x"3b210f",x"381f0e",x"371e0d",x"351d0d",x"39200e",x"39200e",x"3a210f",x"39210f",x"39200f",x"371f0e",x"3a210f",x"3c2310",x"3f2411",x"39210f",x"351e0e",x"361f0e",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442c1b",x"442c1b",x"533d2e",x"453124",x"503829",x"483223",x"503624",x"513726",x"503524",x"513726",x"523523",x"4e3423",x"513928",x"523623",x"573622",x"513625",x"4f3626",x"523827",x"5c3b28",x"5d3c27",x"5b3c29",x"5d3d28",x"5a3b28",x"553726",x"4d3322",x"513627",x"563926",x"543726",x"593c29",x"5b3d27",x"5a3d2a",x"533827",x"533624",x"5c3e29",x"5c3d2a",x"5b3e2b",x"5b3e2b",x"5c402e",x"543b2b",x"563926",x"553622",x"503524",x"533826",x"553724",x"563825",x"5b3c27",x"513723",x"5b3e27",x"61402a",x"583c28",x"6a472f",x"5f3f29",x"573b28",x"5f412b",x"60412c",x"61432f",x"604330",x"5d4230",x"604732",x"5b4130",x"5f4431",x"674a34",x"664833",x"654832",x"61442f",x"5a422e",x"604730",x"60442e",x"63432d",x"5a3c27",x"63402b",x"593a26",x"593a26",x"553522",x"553622",x"593924",x"5d3b26",x"543824",x"5c3c25",x"593924",x"573926",x"4f3422",x"4d3422",x"523624",x"4c3424",x"513625",x"583a27",x"5c3c26",x"563823",x"5a3b26",x"5a3b26",x"523622",x"4e3424",x"462d1e",x"492f1d",x"432c1c",x"432b1b",x"4c2f1c",x"4f321e",x"4a2e1d",x"492f1d",x"452a18",x"462c1a",x"3e2719",x"3e2717",x"3e2a1e",x"3c2b1e",x"37271a",x"502f17",x"150e07",x"150e07",x"150e07",x"150e07",x"442511",x"191109",x"302114",x"342416",x"362618",x"382818",x"372718",x"3b291a",x"3d2b1b",x"382718",x"3d2b1b",x"3d2b1c",x"3d2b1b",x"3a2919",x"3c2a1b",x"44311f",x"3b291a",x"402e1d",x"3d2b1b",x"3b291a",x"3e2c1c",x"402e1d",x"3b2a1a",x"3e2c1c",x"453120",x"412e1d",x"382718",x"3a2819",x"382718",x"3a291a",x"392819",x"372718",x"402d1d",x"402d1c",x"412d1d",x"45311f",x"453120",x"402d1d",x"412e1d",x"43301e",x"44301f",x"422e1d",x"432f1e",x"443120",x"432f1e",x"422e1d",x"453120",x"473321",x"45311f",x"463220",x"412e1d",x"412e1d",x"44311f",x"43301f",x"3d2b1b",x"3e2c1c",x"3f2c1c",x"3f2c1c",x"3b291a",x"3a2819",x"3a2819",x"352517",x"342416",x"382718",x"392819",x"3b2a1a",x"372718",x"362618",x"3a291a",x"3d2b1c",x"3a2819",x"3f2c1c",x"3a2819",x"382718",x"352517",x"362617",x"362617",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f08",x"170f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"24160b",x"1d1108",x"1d1108",x"1f1208",x"201309",x"211309",x"251509",x"231409",x"24150a",x"231409",x"221409",x"231409",x"1d1208",x"201309",x"221409",x"231409",x"1e1209",x"1f1208",x"23150a",x"211409",x"1f1309",x"221409",x"231409",x"221409",x"211409",x"221409",x"25160b",x"23150a",x"221409",x"1f1309",x"24150a",x"25160a",x"211409",x"26170a",x"23150a",x"26160a",x"23150a",x"221409",x"221409",x"26160a",x"1f1208",x"1d1108",x"1f1209",x"1a1108",x"180f07",x"1c1108",x"180f08",x"1b1008",x"190f08",x"1c1108",x"201309",x"1b1108",x"1f1309",x"1f1309",x"231509",x"1f1309",x"201309",x"201309",x"1d1108",x"1f1208",x"1e1208",x"221409",x"231409",x"211409",x"231409",x"221409",x"1f1209",x"1f1209",x"2d1a0b",x"1c1108",x"1b1008",x"1a1008",x"1a1008",x"191008",x"191008",x"191008",x"000000",x"1d1208",x"1d1208",x"26170c",x"3c210f",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"1d1208",x"2a190b",x"150e07",x"150e07",x"150e07",x"331d0d",x"150e07",x"150e07",x"291e17",x"150e07",x"150e07",x"2d190b",x"2d190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2a190b",x"2c190b",x"37200f",x"321c0c",x"381f0d",x"351d0d",x"331c0c",x"351e0d",x"311b0c",x"321c0c",x"39200e",x"3b220f",x"351e0d",x"371f0e",x"3c220f",x"3f2410",x"361e0d",x"3c2310",x"3f2411",x"3b2210",x"402512",x"3c230f",x"39200e",x"3f2410",x"412511",x"432712",x"3a210f",x"351d0d",x"371e0d",x"3c2310",x"3a2210",x"3c2311",x"422712",x"402512",x"422712",x"422712",x"432813",x"3e2411",x"3c220f",x"442914",x"412814",x"472c16",x"432914",x"3f2511",x"392310",x"34200e",x"36210e",x"3f2410",x"39210f",x"3a210e",x"38200e",x"3e2310",x"3e2410",x"402511",x"432712",x"462914",x"432612",x"3e2310",x"3d2310",x"3e2310",x"422612",x"3f2511",x"412612",x"412612",x"442813",x"3e2310",x"3c230f",x"3c220f",x"3a210f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412919",x"412919",x"503b2c",x"4a3325",x"4b3627",x"503523",x"4f3524",x"4f3524",x"533623",x"563721",x"654029",x"563a27",x"5a3c28",x"5a3e2b",x"5c3a24",x"593c2a",x"5e412e",x"654631",x"67452d",x"67432c",x"61432f",x"5b3e2c",x"583c2c",x"5b3d2a",x"563b29",x"533929",x"573a28",x"583c29",x"5d3e29",x"543a29",x"5f412d",x"573b28",x"533623",x"5b3b26",x"593926",x"5f3f29",x"5c3e2a",x"5e402a",x"5b3d28",x"5d3e2a",x"62412c",x"62422e",x"613f29",x"61432e",x"5c3e2a",x"583a28",x"563a28",x"5d3e2b",x"5d3f2a",x"62422d",x"62422c",x"6d472e",x"61412c",x"60432e",x"62422c",x"644530",x"543b2a",x"583d2d",x"5d432f",x"684a31",x"704d33",x"65432b",x"5d4029",x"523b28",x"553a27",x"5f3f2b",x"593a26",x"563a27",x"5d3c29",x"623f2a",x"5c3d29",x"60402b",x"5e3d27",x"5f3d26",x"613e27",x"5a3b25",x"5c3b25",x"5b3b25",x"5d3d26",x"5a3b26",x"5c3c25",x"4e3422",x"4f3625",x"4f3726",x"4b3323",x"4e3423",x"523827",x"543826",x"523726",x"563a27",x"553723",x"523725",x"503422",x"422b1c",x"473020",x"3b281b",x"412b1c",x"412a1c",x"462e1e",x"563420",x"4d2e19",x"4f311b",x"492c18",x"442a1a",x"442b1a",x"362417",x"38261a",x"34271d",x"4e2d16",x"150e07",x"150e07",x"150e07",x"150e07",x"472711",x"1e150b",x"342416",x"382819",x"332416",x"372718",x"352517",x"3b2a1b",x"392819",x"392819",x"3f2d1c",x"3e2b1b",x"3f2d1d",x"362618",x"3c2b1c",x"402e1e",x"3c2b1b",x"422f1f",x"3d2b1b",x"402d1c",x"432f1e",x"362618",x"3a281a",x"3e2c1c",x"3f2d1d",x"443221",x"3c2b1c",x"3f2d1d",x"3e2c1c",x"4a3523",x"3a291a",x"3f2d1c",x"412d1d",x"422f1f",x"44311f",x"422f1e",x"3d2b1c",x"422f1e",x"453120",x"453120",x"422f1e",x"432f1f",x"453120",x"432f1e",x"473321",x"453120",x"443120",x"473422",x"443120",x"463220",x"483321",x"402d1c",x"412e1d",x"3b291a",x"402d1d",x"432f1e",x"3b2a1b",x"3c2b1c",x"3b2a1b",x"3d2b1c",x"3c2b1b",x"443120",x"3e2c1c",x"3e2c1c",x"3d2b1b",x"3d2b1c",x"3c2b1b",x"382819",x"3a291a",x"382819",x"3c2b1b",x"372718",x"322315",x"362618",x"3a291a",x"362617",x"362617",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26160a",x"25160a",x"231509",x"211309",x"321d0d",x"191008",x"150e07",x"150e07",x"1e1208",x"191008",x"1e1209",x"191008",x"170f07",x"1c1108",x"1b1108",x"150e07",x"180f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"1d1108",x"150e07",x"150e07",x"1f1309",x"1a1108",x"1d1209",x"181008",x"150e07",x"150e07",x"1b1108",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"27170a",x"1e1208",x"1f1209",x"1f1208",x"201309",x"221409",x"221409",x"231409",x"231509",x"24150a",x"25160a",x"231509",x"241509",x"231509",x"231409",x"231409",x"231509",x"25160a",x"25160a",x"25160a",x"221409",x"24150a",x"211309",x"231409",x"221409",x"211309",x"221409",x"231509",x"231409",x"241509",x"25160a",x"24150a",x"24150a",x"24150a",x"231409",x"231409",x"25160a",x"24150a",x"24160a",x"24150a",x"221409",x"231409",x"231509",x"24150a",x"24160a",x"221409",x"201208",x"24150a",x"25160a",x"26170a",x"27170b",x"28180b",x"28180b",x"28180b",x"28180b",x"28180b",x"25150a",x"231409",x"26170a",x"26180b",x"27180b",x"25160a",x"22150a",x"1f1309",x"1e1208",x"1f1309",x"1f1309",x"1d1208",x"1d1108",x"1d1208",x"1d1108",x"1c1108",x"1e130b",x"1d130b",x"1c130b",x"1c120b",x"1c120b",x"000000",x"1d1209",x"1d1209",x"28180c",x"402410",x"150e07",x"150e07",x"150e07",x"2c190b",x"150e07",x"2b190b",x"150e07",x"150e07",x"150e07",x"2f1b0d",x"150e07",x"150e07",x"2c2119",x"150e07",x"150e07",x"2c190a",x"2c190a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"180f07",x"301c0c",x"311c0d",x"38200f",x"371f0e",x"381f0e",x"3a200e",x"361e0d",x"2d190a",x"321c0c",x"2e190b",x"351d0d",x"3a210f",x"331d0d",x"2e1a0c",x"3a210f",x"38200e",x"3a220f",x"38200f",x"3c220f",x"3b2210",x"3b2210",x"3a210f",x"3a210f",x"3a210f",x"39200f",x"3d2310",x"3d2411",x"39210f",x"3c2310",x"402512",x"3e2511",x"3f2511",x"3b220f",x"3b220f",x"3d2310",x"3a210f",x"2f1c0c",x"2f1b0c",x"3d2310",x"412612",x"402512",x"422813",x"382310",x"3e2511",x"432612",x"3c220f",x"3f2411",x"422612",x"402411",x"402612",x"422712",x"3e2411",x"442813",x"3c2311",x"412712",x"3a210f",x"3b210f",x"3c220f",x"3e2411",x"3c2311",x"3f2511",x"422612",x"402512",x"402511",x"402511",x"3e2310",x"3f2410",x"3d2210",x"39200e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2516",x"3d2516",x"4b3b2f",x"523a2a",x"4d3627",x"453326",x"4c3223",x"503625",x"5e3d27",x"553a27",x"603f29",x"64442f",x"593c29",x"583924",x"5a3c26",x"63422c",x"62432e",x"65452f",x"61402c",x"63442f",x"63442f",x"5e422f",x"573d2c",x"5e3f2d",x"5d412e",x"4e3829",x"4c3628",x"503829",x"573c2b",x"593e2b",x"5f412d",x"593d2b",x"583c2a",x"634330",x"614431",x"5f412e",x"5b412f",x"60422e",x"62422d",x"61412a",x"69442d",x"64412b",x"5d3e2b",x"5c3f2d",x"65452f",x"61412c",x"61422e",x"66462f",x"5f422d",x"5f412c",x"5c402c",x"5d412e",x"5a3d2b",x"5a3c28",x"583b28",x"5a3d29",x"583d2b",x"5e402b",x"624430",x"634431",x"634731",x"604330",x"654631",x"64412b",x"61432f",x"60402c",x"593b28",x"6a462e",x"6c482f",x"5f3f29",x"563b29",x"5d3f2b",x"5d3f2a",x"593b27",x"583926",x"583825",x"5d3c26",x"643f26",x"593b27",x"593a25",x"513523",x"513624",x"4a3120",x"563723",x"4f3424",x"452f21",x"4c3424",x"4a3222",x"4e3525",x"5a3c28",x"563725",x"4c3220",x"553c2b",x"432d1f",x"3e2b1f",x"492f1d",x"412b1c",x"412817",x"462b19",x"472c1a",x"4b2f1c",x"4d301c",x"442a19",x"482c1a",x"482d1c",x"432919",x"442f21",x"37291e",x"482912",x"150e07",x"150e07",x"150e07",x"150e07",x"462812",x"1e140b",x"342416",x"362617",x"3a291a",x"3a2a1a",x"3d2b1b",x"3a291a",x"392819",x"43301f",x"43301f",x"402e1e",x"412e1d",x"443221",x"3d2b1c",x"433121",x"422f1f",x"3e2d1d",x"433020",x"3d2b1c",x"412e1e",x"3b2a1b",x"3d2b1c",x"3f2d1d",x"402e1e",x"443120",x"443120",x"44311f",x"473322",x"443120",x"412e1d",x"402d1d",x"45311f",x"463220",x"402e1e",x"463220",x"473321",x"473320",x"473321",x"503a27",x"473320",x"473321",x"473322",x"4a3624",x"483321",x"513b27",x"4a3523",x"4a3624",x"4c3825",x"453221",x"483422",x"422f1f",x"45311f",x"443120",x"453120",x"453220",x"3f2d1d",x"3f2d1d",x"423020",x"43301f",x"402e1e",x"3f2d1e",x"3f2d1c",x"422f1e",x"3f2d1c",x"402e1d",x"3c2a1b",x"3d2b1c",x"3f2d1d",x"3f2d1d",x"412e1d",x"372719",x"362618",x"3c2a1b",x"3c2b1b",x"3a291a",x"3a291a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26160a",x"26160a",x"25160a",x"211409",x"150e07",x"25160a",x"24150a",x"27170a",x"28180b",x"29180b",x"27160a",x"28180b",x"29180b",x"28180b",x"29180b",x"27170b",x"28180b",x"2d1b0c",x"2a190b",x"26160a",x"27170a",x"2a190b",x"29180b",x"27170a",x"28170b",x"221409",x"28180b",x"29190b",x"2b1a0c",x"2d1a0c",x"2c1a0c",x"29170b",x"2c1a0c",x"2d1a0c",x"28170b",x"2b1a0c",x"2e1b0d",x"2b190b",x"211409",x"24150a",x"27170b",x"211409",x"27170a",x"27160a",x"221409",x"28170b",x"26170a",x"28170b",x"1f1309",x"2a180b",x"24150a",x"24150a",x"28170a",x"26160a",x"26160a",x"2a180b",x"27170b",x"27170b",x"1f1309",x"29180b",x"26160a",x"231509",x"201309",x"28170a",x"251509",x"241509",x"231409",x"241509",x"221409",x"221409",x"351d0d",x"160e07",x"231409",x"231409",x"231409",x"231409",x"241509",x"25160a",x"26160a",x"27170a",x"27170b",x"27170a",x"26160a",x"25160a",x"25150a",x"26160a",x"26160a",x"25160a",x"24150a",x"25160a",x"26160a",x"25160a",x"241509",x"241509",x"231509",x"211309",x"211308",x"211309",x"211308",x"24150a",x"25160a",x"24150a",x"24150a",x"24150a",x"24150a",x"25160a",x"25160a",x"25160a",x"26160a",x"26160a",x"25160a",x"26160a",x"241509",x"25160a",x"26160a",x"27170b",x"26160a",x"27170b",x"27170b",x"26160a",x"26160b",x"24150a",x"25160a",x"25160a",x"25160a",x"24150a",x"24150a",x"24150a",x"25160a",x"25160a",x"24160a",x"211409",x"22150a",x"211409",x"211409",x"211409",x"201409",x"201409",x"201409",x"1e1209",x"1f140a",x"20160d",x"21180f",x"20170f",x"20160f",x"1e160f",x"1e160f",x"000000",x"1d1209",x"1d1209",x"28190c",x"3b210e",x"150e07",x"150e07",x"150e07",x"2e1a0c",x"150e07",x"2a180b",x"150e07",x"150e07",x"150e07",x"331d0d",x"150e07",x"150e07",x"27170a",x"150e07",x"160e07",x"321b0b",x"321b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"26150a",x"150e07",x"23150a",x"2b190c",x"2c190b",x"2f1a0c",x"28160a",x"301c0c",x"311d0d",x"321d0d",x"331d0d",x"37200e",x"2e1b0c",x"29180b",x"29180b",x"2e1a0b",x"2c190b",x"2b180b",x"2c180b",x"331d0d",x"361f0f",x"311d0d",x"2c190b",x"2f1b0c",x"2b190b",x"321c0d",x"301c0c",x"2c190b",x"311b0c",x"2c190b",x"25160a",x"2f1b0c",x"301b0c",x"29160a",x"201107",x"28170a",x"2f1a0b",x"301b0c",x"311c0d",x"311c0d",x"331d0d",x"2e1b0c",x"331d0d",x"311c0d",x"331d0e",x"331e0e",x"321d0d",x"321d0d",x"311c0d",x"331d0d",x"331e0e",x"3a2210",x"311d0d",x"311c0c",x"321d0d",x"2f1a0c",x"38210f",x"321c0c",x"37200f",x"37200e",x"361f0e",x"2e1a0b",x"331d0d",x"25160a",x"28170b",x"402511",x"150e07",x"3f2410",x"351e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2717",x"3f2717",x"463629",x"473224",x"4d3628",x"4d3627",x"462e1f",x"483021",x"4a3121",x"4d3323",x"543926",x"5b3d28",x"5f3d26",x"5b3b28",x"5d3c25",x"593b28",x"513829",x"5b3d2b",x"5b3d2b",x"60422e",x"6f4a32",x"5a3e2b",x"60412c",x"583b28",x"533929",x"503626",x"5c3f2c",x"583c29",x"5e3e2b",x"583a27",x"5f422f",x"664530",x"5c3d29",x"593926",x"573927",x"563a28",x"563827",x"533b2b",x"60402a",x"63412b",x"5f402c",x"593b27",x"593c29",x"5a3d2a",x"5f412d",x"5c4130",x"5b4131",x"583f2e",x"593e2c",x"573d2d",x"5c4130",x"523d2e",x"45362d",x"563e30",x"5b3f2d",x"5c3f2d",x"5c3f2d",x"5f4331",x"5c3e2b",x"583d2c",x"5f3f2a",x"5a3d29",x"64422b",x"5c3c26",x"62412c",x"5a3d29",x"5b3a24",x"5c3e2a",x"65442d",x"5b3d29",x"553a28",x"593b28",x"4e3424",x"523726",x"513624",x"523523",x"61412a",x"593a24",x"593b27",x"523624",x"4e3322",x"513523",x"4b3222",x"523725",x"573825",x"4c3322",x"563926",x"4d3523",x"493121",x"563622",x"533523",x"533826",x"483120",x"483223",x"452e1e",x"4d3423",x"462f1f",x"422b1c",x"462c1a",x"3c2617",x"4a2c18",x"4a2c1a",x"472b18",x"432817",x"3c2414",x"442c1c",x"342217",x"322820",x"462711",x"150e07",x"150e07",x"150e07",x"150e07",x"472812",x"191109",x"3a291a",x"3d2c1d",x"39281a",x"362517",x"392819",x"322315",x"3b291a",x"3d2c1c",x"402e1e",x"423120",x"3f2d1d",x"412f1f",x"3c2b1c",x"3a291a",x"392819",x"382718",x"392819",x"3a2819",x"382717",x"392717",x"382717",x"372718",x"382617",x"392819",x"44311f",x"412f1e",x"44301f",x"453220",x"3f2d1d",x"463221",x"43301f",x"483422",x"433120",x"493523",x"453220",x"463120",x"463220",x"422f1d",x"4a3422",x"483422",x"4a3523",x"4e3a26",x"4c3825",x"4b3725",x"4d3825",x"3f2c1c",x"432f1e",x"3f2d1c",x"3a2919",x"3f2c1b",x"3e2b1a",x"3e2a1a",x"402c1b",x"3c2a1a",x"392717",x"3b291a",x"3d2c1c",x"402e1d",x"3f2d1c",x"3f2d1d",x"473322",x"443120",x"453120",x"43301f",x"433120",x"433020",x"453220",x"3f2c1c",x"3c2a1b",x"382718",x"39281a",x"3a291a",x"3b2a1b",x"3b2a1b",x"3b2a1b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341d0c",x"39200e",x"432510",x"3c210f",x"3b210f",x"3a200e",x"3d220f",x"3d220f",x"3c220f",x"3a200e",x"3b210f",x"3a200f",x"3d230f",x"3d240f",x"3e2410",x"3d220f",x"3f2410",x"39200e",x"381f0e",x"361e0d",x"371f0d",x"381f0d",x"3c220f",x"3a200e",x"39200e",x"361e0d",x"39200e",x"3a200f",x"39200e",x"39200e",x"3a200e",x"371e0d",x"391f0d",x"361e0d",x"301a0b",x"341c0c",x"381e0d",x"371e0d",x"381e0d",x"371e0d",x"361d0d",x"351d0d",x"361e0d",x"351d0d",x"39200e",x"39200e",x"3c220f",x"402411",x"3e2310",x"371e0d",x"3b200e",x"3b200f",x"3c2310",x"3e2411",x"402510",x"3e240f",x"412511",x"402410",x"3a210f",x"3c220f",x"3e220f",x"3c210e",x"381f0d",x"391f0e",x"391f0d",x"412411",x"422611",x"412510",x"371e0d",x"381f0d",x"150e07",x"201308",x"201309",x"201309",x"211309",x"221409",x"231409",x"231409",x"231409",x"24150a",x"25160a",x"25160a",x"25150a",x"24150a",x"211309",x"201208",x"221409",x"231409",x"24150a",x"26160a",x"25160a",x"25160a",x"241509",x"221409",x"231409",x"25150a",x"25160a",x"26160a",x"231509",x"26160a",x"26160a",x"26160a",x"24150a",x"231509",x"231409",x"231409",x"241509",x"26160a",x"26170b",x"26160a",x"24150a",x"25160a",x"24150a",x"25160a",x"24150a",x"231409",x"231409",x"24150a",x"241509",x"241509",x"221409",x"1c1007",x"1d1108",x"221409",x"231409",x"231509",x"23150a",x"231509",x"211409",x"221409",x"221409",x"23150a",x"22150a",x"22150a",x"211409",x"201309",x"1e1208",x"1f1309",x"1e1209",x"1d1208",x"1e130b",x"1d130b",x"1e140d",x"1d140d",x"1c140c",x"1c140c",x"000000",x"1e1209",x"1e1209",x"2a190d",x"371e0d",x"150e07",x"201309",x"150e07",x"180f08",x"160e07",x"150e07",x"331d0d",x"150e07",x"221409",x"150e07",x"2f1b0c",x"150e07",x"1e1208",x"150e07",x"1c1108",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"38200f",x"28170a",x"3e2310",x"472914",x"432712",x"412410",x"3e220f",x"3d210e",x"412511",x"3f2410",x"3f2411",x"402410",x"422612",x"3f2310",x"412511",x"462813",x"432712",x"452813",x"3c210f",x"3c210e",x"3e230f",x"3f2410",x"3a210e",x"432611",x"422611",x"381f0e",x"371f0e",x"3d2210",x"3e2310",x"3f2410",x"432612",x"422612",x"492b15",x"412511",x"432612",x"3b210f",x"402310",x"472912",x"432612",x"412411",x"432712",x"462813",x"412511",x"412410",x"442611",x"462813",x"422611",x"462913",x"462813",x"412410",x"412511",x"442711",x"442712",x"472914",x"452712",x"422511",x"422511",x"3d210f",x"442611",x"311c0c",x"331c0c",x"1e1208",x"301b0c",x"150e07",x"3e2310",x"341d0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412918",x"412918",x"543f31",x"4b3425",x"503827",x"583a27",x"513625",x"4f3526",x"4b3222",x"493122",x"583824",x"583a27",x"5a3b25",x"634029",x"5e3e2b",x"624028",x"5b3b26",x"5a3d2a",x"5e412e",x"583d2b",x"61432f",x"5e402b",x"5d402e",x"593f2f",x"5e3f2a",x"60412d",x"5a3e2b",x"553825",x"533727",x"553a29",x"553b29",x"593c2a",x"563c2b",x"593e2c",x"593c2a",x"563b2a",x"5a402f",x"614534",x"563d2d",x"5c4332",x"5c4131",x"563b2a",x"5f4433",x"5f4332",x"5f422e",x"5e4230",x"5c402e",x"543b2b",x"503727",x"583925",x"5c3c29",x"5c3e2a",x"4f3828",x"5a3f2d",x"5d3f2b",x"5b3d2a",x"573b28",x"543623",x"5a3e2b",x"5b3d29",x"5e3e2a",x"603f28",x"593b26",x"5a3d2a",x"5b3d2b",x"573926",x"573a26",x"5b3f2d",x"62402b",x"583b29",x"4f3828",x"4c3323",x"583b28",x"523725",x"513623",x"5b3c26",x"553623",x"583622",x"503523",x"4c3221",x"503421",x"4d3322",x"4c3323",x"4d3321",x"513625",x"4c3424",x"533826",x"543825",x"5b3e2a",x"5f412e",x"503726",x"533726",x"4a3223",x"452f20",x"452d1e",x"3f291a",x"4a3021",x"51331f",x"462e1e",x"53341f",x"462b19",x"482c18",x"4a2c16",x"472b17",x"3b2516",x"52311c",x"3d281b",x"36291f",x"492b14",x"150e07",x"150e07",x"150e07",x"150e07",x"482913",x"231a10",x"3d2d1e",x"3d2c1d",x"38281a",x"3b2a1b",x"3e2d1d",x"3b2a1b",x"3e2d1d",x"402e1f",x"493523",x"423020",x"41301f",x"433120",x"412f1f",x"3e2c1c",x"402d1d",x"422f1f",x"3d2b1b",x"3c2a1b",x"3b2a1a",x"3b2b1b",x"443220",x"402f1e",x"3e2d1e",x"422f1f",x"463423",x"473323",x"473422",x"453221",x"4b3726",x"4a3624",x"463323",x"493625",x"4b3827",x"4f3b28",x"4e3926",x"493523",x"4f3a27",x"493624",x"4e3926",x"4f3a27",x"493523",x"4e3926",x"493523",x"493523",x"4d3826",x"422f1d",x"422e1d",x"3b291a",x"3e2a1a",x"3c2919",x"3d2b19",x"422f1d",x"402d1c",x"3d2b1b",x"3d2b1c",x"3e2c1c",x"422f1f",x"412f1f",x"402d1d",x"42301e",x"443120",x"4a3624",x"4a3523",x"4b3824",x"4d3926",x"493524",x"43301f",x"433120",x"3f2d1d",x"3c2a1b",x"3f2d1d",x"3f2d1e",x"3e2d1d",x"3c2b1c",x"3c2b1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"28170a",x"28170a",x"150e07",x"150e07",x"150e07",x"1d1208",x"211409",x"1c1108",x"1f1208",x"1d1208",x"150e07",x"150e07",x"1e1208",x"1d1108",x"1f1208",x"1f1209",x"201309",x"1f1209",x"25160a",x"24150a",x"26170b",x"23150a",x"211409",x"201309",x"221409",x"24150a",x"201309",x"221409",x"25160a",x"27170a",x"24150a",x"25160a",x"25150a",x"28170a",x"221409",x"211409",x"201309",x"221409",x"241509",x"23150a",x"221409",x"1d1208",x"24150a",x"231409",x"1d1208",x"1d1108",x"1d1208",x"1f1209",x"1c1108",x"1e1208",x"1c1108",x"180f07",x"150e07",x"150e07",x"150e07",x"180f08",x"23150a",x"1f1209",x"1f1208",x"191008",x"150e07",x"1e1209",x"1e1209",x"201309",x"1f1309",x"1d1208",x"24150a",x"1e1209",x"201309",x"381f0e",x"361d0d",x"231409",x"26160a",x"29170a",x"28170a",x"29170b",x"150e07",x"341d0d",x"341e0d",x"351e0e",x"361f0e",x"351f0e",x"331d0e",x"37200f",x"351e0e",x"361f0e",x"341d0d",x"331d0d",x"331d0d",x"341d0d",x"311c0c",x"301a0b",x"331c0c",x"311b0b",x"2d1a0b",x"301b0b",x"321c0c",x"301b0c",x"301b0b",x"311b0c",x"311b0c",x"351e0d",x"311b0c",x"321c0c",x"361e0d",x"351e0d",x"391f0e",x"361e0d",x"371f0e",x"341d0d",x"371f0e",x"38200e",x"361e0e",x"361e0d",x"321c0c",x"351e0d",x"351e0d",x"3a200f",x"371f0e",x"341d0d",x"321c0c",x"331c0c",x"331d0c",x"321c0c",x"351d0d",x"361e0e",x"38200e",x"371f0e",x"3a210f",x"39200f",x"331c0c",x"341d0d",x"371f0e",x"3b220f",x"39200f",x"321d0d",x"371f0d",x"361f0e",x"311c0c",x"371f0e",x"361e0d",x"3f2410",x"36200f",x"321d0f",x"24160c",x"24160c",x"000000",x"23160b",x"23160b",x"2a1a0d",x"361d0d",x"2e1a0b",x"150e07",x"150e07",x"1d1209",x"150e07",x"150e07",x"1e1209",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"2b190b",x"3f2511",x"341e0d",x"2d1a0b",x"3b2210",x"3d2411",x"3d2310",x"321c0d",x"2d190b",x"331c0c",x"361e0d",x"361e0d",x"321d0d",x"351e0d",x"351e0e",x"351f0e",x"361f0e",x"331d0d",x"331d0d",x"361e0d",x"341d0d",x"321c0d",x"351e0d",x"341d0d",x"351d0d",x"2f1a0b",x"2e190b",x"2b170a",x"311b0c",x"321c0c",x"351e0e",x"39200f",x"38200f",x"341d0d",x"331d0d",x"341e0d",x"361f0e",x"341d0d",x"311c0c",x"351f0e",x"331c0d",x"321c0c",x"371f0e",x"351d0d",x"361f0e",x"38210f",x"3c2311",x"3b2210",x"3d2410",x"38200f",x"371f0e",x"331c0c",x"371e0d",x"371f0e",x"3a210f",x"3e2310",x"412611",x"3e2310",x"3b210f",x"472711",x"2d190b",x"3f2310",x"422611",x"452712",x"150e07",x"412511",x"331c0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2818",x"3f2818",x"584335",x"573c2a",x"503827",x"563724",x"563a27",x"553926",x"553927",x"4f3421",x"5a3a24",x"5a3c27",x"563825",x"573c29",x"60402b",x"5e3e2a",x"61422d",x"5b3e2a",x"5e402c",x"563e2d",x"563c2c",x"5a3e2c",x"543a28",x"503726",x"593d2b",x"5f412c",x"5e412e",x"5b3e2b",x"573b2b",x"523828",x"503728",x"543d2d",x"5d412f",x"5e412d",x"5c3f2c",x"573d2c",x"5a3e2d",x"573d2d",x"533a29",x"4b3425",x"573b29",x"5b3d2b",x"513726",x"5c412f",x"593f2f",x"503728",x"4e3525",x"4a3629",x"503a2c",x"563f30",x"5e4535",x"5e4330",x"563e2d",x"573f30",x"563d2c",x"543827",x"5a3d2b",x"513625",x"4c3525",x"563927",x"5a3c27",x"573c2a",x"593d2c",x"593c2a",x"5f422f",x"654530",x"62432f",x"553c2a",x"5d3f2c",x"5c3f2a",x"503b2c",x"553a29",x"513727",x"4e3627",x"523725",x"473224",x"543a27",x"593b28",x"583a26",x"4f3728",x"553928",x"593a27",x"593b27",x"553826",x"543826",x"4e3626",x"4b3526",x"493325",x"4d3525",x"553827",x"5d3f2c",x"553c2c",x"523929",x"4f3727",x"4e3524",x"4f3626",x"573926",x"513523",x"4f3523",x"4d2f1c",x"492d1a",x"472c1b",x"422918",x"402716",x"4f311f",x"462d1c",x"432b1c",x"3e2d22",x"4b2b14",x"150e07",x"150e07",x"150e07",x"150e07",x"452712",x"231a11",x"3c2c1d",x"36271a",x"38291c",x"3e2d1e",x"3d2d1e",x"423121",x"412f1f",x"3f2d1d",x"412f20",x"453221",x"403020",x"412f1f",x"3a2b1b",x"412f1f",x"413020",x"433121",x"423121",x"412f20",x"3c2a1c",x"3e2d1f",x"3f2e1f",x"412f20",x"433122",x"463222",x"443323",x"4a3727",x"483624",x"493625",x"4a3726",x"473524",x"463422",x"463323",x"4b3826",x"412e1f",x"4a3624",x"4a3725",x"483523",x"503c29",x"4e3926",x"463321",x"4c3725",x"493523",x"4d3825",x"4a3421",x"43301e",x"422e1d",x"3b2919",x"412d1d",x"3c2a1a",x"3d2b1a",x"3a2819",x"3b2919",x"3e2c1c",x"3d2b1b",x"3f2d1d",x"3c2a1b",x"402d1d",x"3f2d1d",x"402e1d",x"412f1e",x"443121",x"463221",x"463320",x"493421",x"473321",x"422d1d",x"3e2b1c",x"39281a",x"3f2d1d",x"402f1e",x"3f2d1c",x"382818",x"3a2a1a",x"3b2a1b",x"3b2a1b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"28170a",x"28170a",x"26160a",x"26160a",x"160f07",x"2e1a0b",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"190f07",x"190f08",x"1f1309",x"150e07",x"211409",x"180f08",x"1f1309",x"1d1208",x"231509",x"201309",x"1e1208",x"1c1108",x"1d1208",x"1f1208",x"27160a",x"211309",x"231409",x"1f1309",x"1b1108",x"1f1309",x"221409",x"1b1108",x"201309",x"1e1208",x"1c1108",x"1f1208",x"1b1108",x"150e07",x"1d1208",x"23150a",x"1b1108",x"1b1108",x"1e1208",x"211409",x"201309",x"1d1108",x"25160a",x"1d1208",x"201309",x"150e07",x"1a1008",x"1a1008",x"201309",x"1d1208",x"150e07",x"1c1108",x"1a1008",x"1d1208",x"1f1209",x"1b1108",x"1e1208",x"1e1208",x"24150a",x"201309",x"29180b",x"3e230f",x"39200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"191008",x"191008",x"191008",x"180f08",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"180f08",x"190f08",x"190f08",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"171009",x"19120b",x"1b150e",x"1c150e",x"1e1711",x"1d160f",x"1b150e",x"1b150d",x"1b150d",x"000000",x"1d1108",x"201309",x"28180c",x"351e0d",x"3e291c",x"3e291c",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1209",x"1c1108",x"1c1108",x"000000",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0c",x"150e07",x"180f07",x"2b180b",x"2f1b0c",x"2d1a0c",x"341e0d",x"3c2210",x"3a200f",x"3d2310",x"3a2210",x"3f2411",x"3f2411",x"39200e",x"3f2410",x"3a210f",x"3a210f",x"3c220f",x"3a200f",x"371f0e",x"38200f",x"3c220f",x"39200f",x"3c2310",x"3f2411",x"3e2411",x"3b2210",x"3a210f",x"3e2310",x"3f2411",x"3c2310",x"3f2411",x"412612",x"3f2411",x"3f2410",x"3e2310",x"3c220f",x"3b210f",x"39200e",x"3c220f",x"39200e",x"3a210f",x"3e230f",x"371e0d",x"39200e",x"3e2310",x"3c2310",x"3f2410",x"3e2310",x"3e2410",x"3b2210",x"3b210f",x"3b210f",x"432712",x"3f2410",x"432712",x"432712",x"422612",x"412310",x"371e0d",x"391f0d",x"422410",x"150e07",x"2c190b",x"301a0b",x"2b180a",x"2a180a",x"452712",x"341d0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432918",x"432918",x"553e2f",x"5a4031",x"523828",x"543726",x"593b28",x"513725",x"472f1f",x"533827",x"523625",x"4b3222",x"493123",x"4c3528",x"543827",x"593c2a",x"5e4231",x"5f402d",x"604331",x"5a3e2d",x"563c2b",x"5a4334",x"5c3f2d",x"5c3f2b",x"593d2b",x"5c3f2c",x"553a27",x"5a3f2e",x"5e4331",x"5c3f2c",x"5c4231",x"513828",x"543b2a",x"553a28",x"5c3f2c",x"583b28",x"563a28",x"513624",x"583b28",x"5d3d29",x"523624",x"60412c",x"5f3f2b",x"563c29",x"5c3f2a",x"5a3e2c",x"543828",x"523b2c",x"543b2b",x"5a3d2b",x"5c3f2a",x"5e3f2c",x"5c3e2b",x"533826",x"593d2b",x"563b2b",x"593e2d",x"593d2c",x"583d2b",x"5d4333",x"5a3e2b",x"5a3b29",x"543927",x"573a29",x"593c29",x"5e422f",x"5a3e2b",x"5a4130",x"583f2f",x"593f2d",x"5d412f",x"563c2a",x"5a3d2b",x"553a27",x"5c3d27",x"4b3627",x"4e3524",x"4e3424",x"523624",x"4d3221",x"543624",x"513523",x"533523",x"4f3220",x"503423",x"563926",x"543927",x"553b2a",x"523a2b",x"4f3422",x"553928",x"5a3f2e",x"4d3526",x"573b29",x"543a29",x"4b3425",x"513625",x"523624",x"50321f",x"492e1d",x"492d1c",x"462a18",x"4e311e",x"472c1a",x"482e1c",x"472d1c",x"482e1d",x"412c1d",x"3f220e",x"150e07",x"150e07",x"150e07",x"150e07",x"472711",x"271e15",x"392b1d",x"3d2d1e",x"3f2e20",x"3e2e20",x"3f2e20",x"402f21",x"443223",x"483624",x"443324",x"453323",x"453323",x"433222",x"433223",x"453324",x"433222",x"443223",x"493726",x"423123",x"443324",x"493626",x"443221",x"423120",x"453322",x"443323",x"433223",x"433222",x"4a3626",x"493625",x"4b3827",x"4c3827",x"4d3928",x"4d3a28",x"483624",x"473423",x"4a3726",x"4f3b29",x"4b3827",x"503c2a",x"4e3a29",x"4f3a28",x"4a3726",x"483423",x"4b3624",x"463220",x"453220",x"422f1f",x"44311f",x"473220",x"4b3623",x"422f1e",x"453120",x"483423",x"402d1b",x"3f2d1a",x"412d1c",x"412f1e",x"3f2d1d",x"422f1e",x"473221",x"43301f",x"453221",x"493523",x"453220",x"4b3623",x"483420",x"412e1c",x"3e2c1c",x"3e2c1d",x"422f1e",x"402e1e",x"412e1e",x"422f1f",x"3c2b1c",x"3d2c1d",x"3d2c1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26160a",x"26160a",x"2c190b",x"331c0c",x"321b0b",x"331c0c",x"2d190b",x"321b0c",x"361e0d",x"3a200e",x"3a200e",x"3e220f",x"3c210e",x"3b210e",x"3d220f",x"3c220f",x"381f0d",x"381f0e",x"371e0d",x"381f0d",x"381e0d",x"3b200e",x"3b210e",x"3d220e",x"3c220f",x"3b210f",x"381f0d",x"3d220f",x"3b210f",x"3f2310",x"422611",x"402511",x"452813",x"452812",x"412511",x"442813",x"452813",x"422611",x"3f2410",x"3e2310",x"3d220f",x"3a200e",x"3c210f",x"3d220f",x"412510",x"422611",x"402410",x"3e220f",x"3f2310",x"422611",x"3f2410",x"412410",x"3b200f",x"3a200e",x"39200d",x"391f0d",x"3a200e",x"3c210e",x"3c210f",x"39200e",x"3d220f",x"3d220f",x"3d220f",x"41240f",x"462711",x"442711",x"3b210e",x"3b200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"191008",x"190f08",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"190f08",x"180f08",x"190f08",x"191008",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"191008",x"180f08",x"180f08",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"170f07",x"180f08",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"17110a",x"19130c",x"1c150e",x"1d1610",x"1f1811",x"1f1811",x"1e1711",x"1f1811",x"1d160f",x"1d160f",x"000000",x"1c1108",x"1e1208",x"342114",x"492913",x"423024",x"423024",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1f1208",x"331d0d",x"150e07",x"211409",x"301b0c",x"321c0d",x"2d1a0b",x"29180b",x"3a200f",x"3a210f",x"361f0e",x"351e0e",x"371f0e",x"371f0e",x"38200e",x"3b220f",x"3b210f",x"391f0e",x"371f0e",x"3c2310",x"37200f",x"361f0e",x"39210f",x"38210f",x"3a210f",x"361f0e",x"3c2210",x"38200f",x"371f0e",x"3a210f",x"361f0e",x"39200f",x"412612",x"3b2210",x"3f2512",x"3e2411",x"3c2310",x"39200f",x"3a210f",x"3d2311",x"3d2411",x"3c2310",x"3f2411",x"3e2411",x"3a2210",x"412712",x"3c2311",x"39200f",x"3b210f",x"3a200e",x"371f0e",x"38200f",x"311c0d",x"3d2310",x"3e2411",x"3c230f",x"3f2410",x"3f2511",x"422612",x"3c220f",x"402410",x"3e220f",x"3e220f",x"1d1108",x"371f0e",x"38200e",x"3a210f",x"311c0c",x"3c210f",x"371f0e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2617",x"3e2617",x"4c382a",x"4e382a",x"4d3628",x"4a3022",x"462c1e",x"533523",x"533726",x"533420",x"503321",x"563a29",x"553826",x"573b29",x"593f2e",x"5c3e2d",x"573c2b",x"5b3d2a",x"5d4332",x"5a3f2d",x"573d2c",x"5a3f2d",x"573c2a",x"543b2b",x"583b2a",x"5a3c29",x"5b3e2b",x"583c2a",x"583a27",x"5c3f2d",x"543a2a",x"553a2a",x"563b2a",x"573a27",x"513523",x"563621",x"5c3b25",x"5c3b25",x"603e27",x"5c3a23",x"573824",x"5b3b27",x"5a3a24",x"563824",x"5b3c27",x"513422",x"513726",x"523725",x"533b2c",x"5f412c",x"5f422d",x"64442d",x"5a3f2c",x"5b3e2c",x"5b3f2d",x"5e3e2a",x"5a402d",x"61412c",x"63422c",x"64422c",x"60422f",x"694934",x"62432e",x"624532",x"5a4131",x"5b4130",x"573c2a",x"5c3f2e",x"563d2c",x"5c3f2c",x"5f412d",x"5a3b27",x"5c3f2d",x"5c3d29",x"553b2a",x"5d3e29",x"523727",x"573927",x"503523",x"543622",x"583824",x"563724",x"563723",x"563722",x"573824",x"5c3b26",x"523624",x"523522",x"4c3627",x"533a29",x"583c2a",x"553a29",x"5d412f",x"553c2c",x"543b2d",x"4a3324",x"4c3222",x"503524",x"4b3120",x"4b2c19",x"4e311f",x"462915",x"3f2514",x"3e2515",x"3e2413",x"482d1c",x"3f2517",x"3d291d",x"3f220e",x"150e07",x"150e07",x"150e07",x"150e07",x"3f230f",x"221a13",x"3c2c1d",x"402e20",x"423021",x"3c2b1e",x"402f20",x"433122",x"3e2d1e",x"413021",x"3f2f20",x"3f2f21",x"413122",x"433122",x"3f2f20",x"433122",x"483626",x"443323",x"433223",x"413123",x"483626",x"473423",x"453221",x"402f20",x"3d2c1d",x"453223",x"3f2d20",x"412f21",x"433121",x"423121",x"453322",x"453322",x"473523",x"473423",x"402e1f",x"493523",x"4b3725",x"4c3725",x"453221",x"473524",x"453322",x"443222",x"493624",x"453321",x"433120",x"42301f",x"422f1e",x"45301f",x"443120",x"463321",x"44301f",x"43301f",x"422f1e",x"47311f",x"452f1d",x"3b2919",x"3e2b1a",x"432f1e",x"3c2919",x"3c2919",x"412e1d",x"432f1e",x"412e1d",x"463220",x"483421",x"44301e",x"442f1d",x"412f1d",x"3e2c1c",x"3f2c1c",x"3d2b1b",x"3a2a1a",x"3e2b1b",x"3a2819",x"3f2d1d",x"3b2b1c",x"3b2b1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29170a",x"29170a",x"150e07",x"150e07",x"150e07",x"180f07",x"191008",x"1d1108",x"180f08",x"190f08",x"201309",x"1d1208",x"1c1108",x"191008",x"22140a",x"211409",x"1e1209",x"221409",x"1f1209",x"25160a",x"211409",x"221409",x"25160a",x"26160a",x"26170a",x"211409",x"24160a",x"241509",x"201309",x"231409",x"1f1209",x"24150a",x"231509",x"201309",x"1b1108",x"26160a",x"201309",x"150e07",x"1c1108",x"1a1008",x"1d1108",x"1f1308",x"1c1108",x"1d1208",x"170f07",x"190f08",x"221409",x"221409",x"1e1208",x"27160a",x"231409",x"1c1108",x"1f1208",x"1e1208",x"211309",x"1f1209",x"1f1208",x"231409",x"231409",x"261609",x"26160a",x"211409",x"25160a",x"201309",x"211309",x"291609",x"432611",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"191008",x"1a1008",x"191008",x"191008",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"190f08",x"180f08",x"180f08",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f08",x"180f08",x"180f08",x"180f08",x"180f08",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"17110a",x"1a130c",x"1c160f",x"1e1710",x"201913",x"201a13",x"201913",x"201912",x"1e1811",x"150e07",x"150e07",x"150e07",x"1e1209",x"352115",x"4c2b14",x"4b2d19",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"190f08",x"190f08",x"180f07",x"190f07",x"190f07",x"1a1107",x"1a1007",x"191007",x"180f07",x"180f07",x"170f07",x"170f07",x"160f07",x"160f07",x"170f07",x"170f07",x"201408",x"261809",x"281909",x"2c1a0a",x"351e0c",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"191008",x"311c0c",x"150e07",x"1e1208",x"331d0d",x"311c0c",x"331d0d",x"180f08",x"3f2411",x"432712",x"3f2410",x"3e220f",x"442712",x"452813",x"452813",x"452713",x"432611",x"432611",x"412511",x"432712",x"412511",x"3d2310",x"422611",x"432712",x"442712",x"432511",x"3f220f",x"3e230f",x"3f2310",x"412410",x"412410",x"3e220f",x"3f230f",x"412310",x"3f2410",x"442712",x"412511",x"412511",x"452712",x"442712",x"432511",x"3d220f",x"3f2310",x"462813",x"412511",x"452813",x"412511",x"432611",x"432711",x"462812",x"452711",x"3f2310",x"422611",x"432712",x"492a14",x"442712",x"4a2b15",x"4b2d15",x"492a14",x"452813",x"442712",x"422511",x"150e07",x"2b190b",x"3b220f",x"3a210f",x"38200f",x"331d0d",x"3b200e",x"321c0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2516",x"3e2516",x"4c382b",x"4d392d",x"503626",x"4f3424",x"503525",x"533827",x"5b3b27",x"593c2b",x"5b3a24",x"573824",x"5c3d29",x"5e402d",x"5f4331",x"5b3c28",x"614430",x"5d412e",x"5d4231",x"5d3d29",x"614330",x"533a27",x"523828",x"543622",x"553926",x"5e402b",x"61412b",x"60402a",x"573b29",x"62432f",x"65442e",x"533927",x"5f402c",x"593f2f",x"5a3d29",x"523929",x"64432c",x"61402a",x"60402b",x"624029",x"593a25",x"593c28",x"5b3b27",x"5a3d2b",x"533928",x"593d2c",x"503624",x"523828",x"5a3d2c",x"543c2d",x"593c2a",x"573927",x"5b3e2c",x"5f412c",x"62432f",x"62432f",x"62432e",x"5a3e2d",x"533b2b",x"543929",x"5b3e2b",x"62432c",x"5f3f29",x"65442f",x"603f2b",x"573c2a",x"563e2e",x"513d2e",x"644530",x"593f2d",x"60412d",x"62402b",x"5e3e2a",x"65412a",x"5d3d28",x"5d3e29",x"5d3a23",x"5e3d26",x"543622",x"543621",x"533523",x"573824",x"563722",x"563823",x"5a3c26",x"573724",x"4e3423",x"463022",x"4e3527",x"473022",x"493225",x"4c3020",x"533928",x"553d2f",x"4f3525",x"503828",x"50382a",x"4a3120",x"4e3322",x"482d1b",x"4e2c17",x"482a18",x"432817",x"422615",x"3e2313",x"402515",x"3e2618",x"3e291c",x"3f220e",x"150e07",x"150e07",x"150e07",x"150e07",x"40230f",x"1f1912",x"38291c",x"36281b",x"35271b",x"36271a",x"35261a",x"35261a",x"37281c",x"3a2b1e",x"35271b",x"3b2b1e",x"392b1e",x"37291d",x"37291d",x"392a1e",x"392b1f",x"392a1c",x"3e2e21",x"402f22",x"413021",x"3c2c1d",x"37291c",x"3b2c1d",x"433120",x"3f2d1f",x"423020",x"463221",x"453121",x"473222",x"493623",x"4f3927",x"4a3523",x"473322",x"4a3624",x"463321",x"443120",x"432f1f",x"412f1e",x"473322",x"433020",x"433121",x"433121",x"432f20",x"3e2d1d",x"3b291a",x"3c2b1c",x"3f2c1c",x"3e2c1c",x"382819",x"3b291a",x"382718",x"3d2b1b",x"352516",x"372616",x"352416",x"362516",x"362517",x"362516",x"352517",x"3a2819",x"382718",x"3b291a",x"392719",x"3a2918",x"3e2b19",x"402d1b",x"362517",x"372617",x"322315",x"302114",x"322316",x"352517",x"322215",x"322316",x"332417",x"332417",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29170a",x"231409",x"221409",x"231409",x"150e07",x"180f08",x"1b1108",x"1a1008",x"170f07",x"180f08",x"28170a",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1d1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1209",x"201409",x"1f1309",x"1f1209",x"201309",x"1f1309",x"1e1208",x"1d1208",x"1e1209",x"1e1209",x"1e1208",x"1e1209",x"1e1208",x"1e1208",x"1e1209",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1f1309",x"1c1108",x"1b1108",x"1c1108",x"1a1008",x"190f08",x"190f08",x"180f07",x"1b1008",x"180f07",x"180f07",x"170f07",x"170f07",x"180f07",x"180f08",x"1a1008",x"1b1108",x"180f07",x"170f07",x"170f07",x"160f07",x"170e07",x"160e07",x"150e07",x"191008",x"180f08",x"180f08",x"170f08",x"170f08",x"191008",x"160e08",x"160e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1008",x"170f08",x"150e07",x"160e07",x"150e07",x"150e07",x"191008",x"160e07",x"160e07",x"1a1008",x"170f07",x"170f07",x"1a1008",x"170f07",x"150e07",x"170f07",x"1c1108",x"170f07",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"180f08",x"1c1108",x"1c1108",x"150e07",x"1a1008",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"190f08",x"190f08",x"180f07",x"190f07",x"190f07",x"1a1107",x"1a1007",x"191007",x"180f07",x"180f07",x"170f07",x"170f07",x"160f07",x"160f07",x"170f07",x"170f07",x"201408",x"261809",x"281909",x"2c1a0a",x"351e0c",x"351e0c",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1d1208",x"27170a",x"150e07",x"191008",x"301c0d",x"351f0f",x"321d0e",x"3b2210",x"3c2311",x"3e2411",x"331d0d",x"321c0d",x"331c0d",x"351e0e",x"3a2210",x"361f0e",x"38200e",x"38200e",x"361f0e",x"331c0d",x"311b0c",x"301b0c",x"311b0c",x"321b0c",x"331b0b",x"311b0b",x"331c0c",x"331c0c",x"301b0c",x"361e0d",x"351d0d",x"381f0e",x"38200e",x"38200e",x"351d0d",x"3d220f",x"37200f",x"39210f",x"3a210f",x"3a2110",x"3c2310",x"3d2411",x"3e2310",x"38200f",x"3b220f",x"3c210f",x"3b210f",x"38200e",x"3c2310",x"3d2410",x"39210f",x"361f0e",x"371f0e",x"331d0d",x"3a210f",x"3c2311",x"341f0e",x"3a2110",x"3e2410",x"402512",x"3e2411",x"3c2310",x"150e07",x"27170a",x"38200f",x"341d0d",x"381f0e",x"2e1a0b",x"3f2310",x"351d0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a2315",x"3a2315",x"533b2b",x"553b2a",x"5a3e2d",x"5e3e2a",x"61402b",x"603f2a",x"5f402c",x"5d3c27",x"553521",x"5a3a27",x"5b3c27",x"603f2a",x"664633",x"5e422f",x"5f402c",x"593a28",x"5e402d",x"63432e",x"64442f",x"60412e",x"563d2c",x"5b3f2c",x"573b28",x"65432c",x"65452f",x"5f3e2a",x"60402e",x"5d402d",x"5a3d2b",x"593c28",x"5a3d2b",x"583c29",x"5c3e2b",x"5c3c28",x"573927",x"543929",x"503524",x"4c3526",x"563724",x"4e3322",x"4b3324",x"523829",x"573c2b",x"583e2d",x"573d2d",x"573d2c",x"573c2c",x"5e422e",x"573c2b",x"583e2d",x"573c2a",x"5c3d28",x"563a27",x"61402a",x"5e3d27",x"5b3c28",x"5d3e2b",x"573b29",x"553724",x"63412b",x"5f402d",x"5f412d",x"634330",x"5e4332",x"5e4432",x"5f422e",x"5f3e28",x"5d3e29",x"573927",x"563928",x"5b3e2b",x"66432c",x"62402a",x"5f3d28",x"5d3d26",x"634128",x"684228",x"5e3c26",x"563622",x"563722",x"4e3321",x"543623",x"583823",x"5a3b26",x"543827",x"553825",x"5b3c28",x"573723",x"543825",x"553b2a",x"513420",x"543a2a",x"513828",x"593d2a",x"543b2a",x"4d3627",x"4b3121",x"4d321f",x"50321d",x"4c2f1a",x"4b2e1c",x"50301b",x"4d2e1a",x"472b1a",x"422a1b",x"432b1c",x"3f210e",x"150e07",x"150e07",x"150e07",x"150e07",x"40230f",x"1c160f",x"1f1710",x"1f1811",x"1f1811",x"1f1811",x"1f1811",x"1f1811",x"1e1711",x"201811",x"211912",x"221b14",x"231c14",x"251d16",x"241d15",x"251d16",x"221c15",x"221b15",x"221b14",x"211a14",x"211b14",x"1f1811",x"1e1711",x"1f1912",x"1d1610",x"1d160f",x"1d1610",x"1d1610",x"1c150f",x"1b150e",x"1b150e",x"1b140d",x"1b150e",x"19120c",x"19120b",x"19120b",x"1b150e",x"1b140d",x"1b140d",x"1d1710",x"1f1811",x"1d1710",x"1d1610",x"1c150e",x"19130c",x"19120b",x"171009",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"181008",x"191109",x"191109",x"191109",x"191109",x"191109",x"191109",x"191109",x"191109",x"191109",x"1b1108",x"1b1209",x"1e140a",x"211509",x"211509",x"1c1208",x"1b1208",x"181008",x"181008",x"181008",x"191008",x"181008",x"191109",x"1a120b",x"1a120b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"231409",x"150e07",x"180f08",x"1b1108",x"1a1008",x"170f07",x"180f08",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1d1208",x"1d1208",x"1e1209",x"1e1208",x"1e1208",x"1f1209",x"1f1309",x"201309",x"201309",x"201309",x"1f1209",x"1e1208",x"1f1209",x"201309",x"201309",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1e1208",x"1e1209",x"1f1209",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1f1209",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"191008",x"180f08",x"180f07",x"180f07",x"180f07",x"180f08",x"190f08",x"180f07",x"180f07",x"180f08",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f07",x"190f08",x"191008",x"191008",x"191008",x"191008",x"191008",x"191008",x"1b1008",x"1a1007",x"1a1007",x"191007",x"191007",x"160f07",x"150e07",x"160e07",x"160f07",x"170f07",x"191007",x"1f1408",x"1e1308",x"261809",x"211508",x"1f1408",x"27170a",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1d1208",x"29180b",x"150e07",x"150e07",x"211309",x"28160a",x"241509",x"2b180b",x"3c2310",x"381f0e",x"371e0e",x"3b210f",x"3d2310",x"412611",x"3d2310",x"371f0e",x"381f0e",x"381f0e",x"3a210f",x"3a210f",x"381f0e",x"371f0d",x"3a200e",x"381f0e",x"3c210f",x"351d0d",x"321c0c",x"321c0c",x"311b0b",x"321b0b",x"3b210e",x"3b200e",x"3d2210",x"371f0e",x"3a210f",x"3b210f",x"3b220f",x"3f2410",x"3c220f",x"3f230f",x"371e0d",x"371e0d",x"351d0d",x"371e0d",x"3b210f",x"432612",x"3f2511",x"3f2411",x"412511",x"3b210f",x"3c210f",x"3a200e",x"402410",x"371f0e",x"3c220f",x"3a210f",x"39200f",x"3b220f",x"422511",x"412511",x"422611",x"3d220f",x"462812",x"150e07",x"2e1a0b",x"331d0d",x"341d0d",x"2c190b",x"3d220f",x"361e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"392215",x"392215",x"563d2c",x"5f4432",x"6d4a33",x"62412c",x"5f3e29",x"5f3d28",x"5e3f2b",x"563825",x"5c3b25",x"5b3823",x"5b3b25",x"5f402b",x"60422f",x"5f402c",x"644430",x"644734",x"694b36",x"654632",x"60412d",x"583a28",x"513726",x"553624",x"5c3c28",x"523521",x"533623",x"5a3b28",x"5b3d29",x"613f2a",x"69432b",x"60402a",x"5a3d2a",x"5c3e2a",x"583c2b",x"573b28",x"563b29",x"553a29",x"61422f",x"553725",x"563c2a",x"5e3f2b",x"5a3c29",x"513727",x"4f3525",x"513422",x"563a29",x"573b29",x"563c2c",x"5c3e2c",x"573d2d",x"513a2b",x"5a3e2b",x"5d412d",x"5e4331",x"5b3f2d",x"61412c",x"5c4130",x"4c3525",x"553a29",x"553c2c",x"573c2b",x"5c3e2a",x"60412d",x"5f422f",x"583e2d",x"5f422f",x"593d2a",x"5a3f2d",x"5a3c2a",x"5e412e",x"5c3d29",x"593b28",x"64402a",x"5f3e27",x"5c3b24",x"593823",x"643f28",x"563622",x"5c3b24",x"54331f",x"4f311d",x"4d311f",x"533521",x"4b2f1e",x"523521",x"523523",x"513524",x"5f3c27",x"583a26",x"563724",x"492f1f",x"4b3222",x"523725",x"5d3e2b",x"5b3a27",x"4c3324",x"4a3224",x"4a3223",x"462e1e",x"4b2f1d",x"412817",x"482a15",x"50311d",x"55351d",x"4e311b",x"4e321d",x"442d1d",x"40230e",x"150e07",x"150e07",x"150e07",x"150e07",x"3c210e",x"19130c",x"21180f",x"211810",x"21180f",x"20170f",x"21180f",x"21180f",x"20160d",x"1f160d",x"1f160d",x"20180f",x"251b12",x"241a12",x"261c13",x"241b12",x"241a12",x"241b13",x"231a11",x"271e15",x"251b12",x"241b11",x"261b12",x"1f170e",x"1f170e",x"21180f",x"231910",x"22190f",x"22180f",x"231a10",x"231a10",x"241a11",x"241a11",x"241a10",x"241a10",x"241a11",x"261c13",x"271d14",x"2a2016",x"291f16",x"281d14",x"261c13",x"251a11",x"231910",x"24190f",x"241a10",x"20160c",x"23180e",x"23180d",x"20160c",x"23180e",x"21170d",x"24180e",x"20160c",x"22170d",x"21170c",x"20160c",x"21160c",x"22170d",x"1f150b",x"1f150b",x"20160c",x"21160c",x"22170d",x"24190d",x"261a0d",x"261a0d",x"23180d",x"23180d",x"23180d",x"21170d",x"21160d",x"20160c",x"20150c",x"20150c",x"20150c",x"20150c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1c1108",x"1d1108",x"1e1209",x"201309",x"1f1309",x"201309",x"1f1309",x"1f1208",x"1e1208",x"1f1208",x"1e1208",x"1f1209",x"1f1209",x"1f1309",x"1e1208",x"1e1208",x"1e1208",x"1e1209",x"1d1108",x"1e1209",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1d1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1a1008",x"1a1008",x"191008",x"191008",x"180f07",x"180f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f08",x"191008",x"191008",x"191008",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"190f08",x"191008",x"191008",x"1a1008",x"1b1008",x"1a1007",x"191007",x"191007",x"170e07",x"180f07",x"170f07",x"160f07",x"170f07",x"180f07",x"181007",x"1c1208",x"221608",x"231608",x"261809",x"231608",x"1f1408",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1a1008",x"251509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"341f0e",x"39210f",x"361e0d",x"39200f",x"3e2310",x"3d2310",x"3b210f",x"3c2310",x"3d2310",x"39200e",x"3a210f",x"39200f",x"3a200f",x"381f0e",x"39200e",x"3c220f",x"3b2210",x"37200e",x"311c0c",x"331c0c",x"351d0d",x"3b210f",x"3e2310",x"3c220f",x"402511",x"3c2310",x"3d2310",x"3e2310",x"3f2410",x"3e2410",x"3a210f",x"402411",x"3e2311",x"432713",x"39210f",x"402511",x"3f2411",x"3f2410",x"402410",x"3f2310",x"3f2410",x"3d220f",x"3e2310",x"3e2310",x"3f2410",x"402511",x"39210f",x"3c2210",x"3a200e",x"3c210f",x"3a200e",x"3c210f",x"3f2411",x"462813",x"432612",x"402310",x"150e07",x"160e07",x"170f07",x"1a1008",x"201309",x"3d220f",x"351f0e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422817",x"422817",x"503c2f",x"573d2d",x"66442e",x"5f3d26",x"5f3d27",x"654129",x"67452d",x"634128",x"63422b",x"613f27",x"67452d",x"69452e",x"684731",x"614533",x"694a36",x"5e3f2a",x"6a4d3b",x"6a4a35",x"664530",x"61422c",x"69432a",x"603e28",x"63432d",x"614028",x"5c3e2b",x"5a3e2d",x"5e3d28",x"643f27",x"5e3c27",x"65422c",x"62412d",x"5d3d29",x"5a3c28",x"5a3d2a",x"583b29",x"5b3e2a",x"5b3c28",x"60412d",x"5e3f2a",x"65432c",x"5c3d28",x"563b2b",x"583e2f",x"5a3f2f",x"644430",x"64432e",x"63442f",x"604330",x"583e2d",x"593f2d",x"593e2d",x"5f3f2a",x"61402a",x"573b27",x"5f3e2a",x"5d3f2b",x"63432f",x"563a26",x"61412c",x"613f29",x"583a26",x"5a3c28",x"5c3e2a",x"5f3c25",x"593a27",x"63432f",x"5f3f2a",x"64422b",x"61412c",x"61412b",x"603e28",x"5e3e29",x"5c3924",x"5c3a25",x"5f3d27",x"633d23",x"603b23",x"573520",x"563825",x"4a3122",x"462e21",x"4c301e",x"492e1d",x"4a3020",x"53331e",x"523520",x"583823",x"563621",x"573824",x"543725",x"5a3d29",x"5d3c27",x"563621",x"573824",x"4f321f",x"4c3424",x"482f1f",x"513320",x"4d2f1d",x"53321b",x"4e301c",x"472a15",x"482b17",x"472d1c",x"422917",x"492f1f",x"452611",x"150e07",x"150e07",x"150e07",x"150e07",x"40230f",x"150e07",x"1e150b",x"20160c",x"1d140b",x"1e140b",x"20160c",x"1d140b",x"20160c",x"20160c",x"1d140b",x"20160c",x"1d140b",x"1f160d",x"21180e",x"20160c",x"22170e",x"23180e",x"231910",x"23190f",x"22170e",x"1f160d",x"21180e",x"23180f",x"23180e",x"21170e",x"21180e",x"23180f",x"261b10",x"261a11",x"251a11",x"21170d",x"24190f",x"22170d",x"21170d",x"20160c",x"251a0f",x"21170e",x"21180e",x"24190f",x"241a0f",x"241a0f",x"24190f",x"25190e",x"22170d",x"23180d",x"23180d",x"20160c",x"21160c",x"21160d",x"20150c",x"21170d",x"21160c",x"20160c",x"20160c",x"24180e",x"23180e",x"20150c",x"20160c",x"21160d",x"21170d",x"22170d",x"22170d",x"22170d",x"24180d",x"271b0f",x"25190d",x"21170c",x"21170c",x"20160c",x"23170d",x"20160c",x"20160c",x"20160c",x"20150c",x"20150b",x"20150b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f08",x"191008",x"1a1108",x"1c1108",x"1c1108",x"1d1208",x"1d1208",x"1e1209",x"1f1209",x"1f1209",x"1f1309",x"1f1309",x"1f1209",x"201309",x"201309",x"201309",x"201309",x"1f1309",x"1f1209",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1f1309",x"1f1209",x"1d1108",x"1d1108",x"1a0f07",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1d1208",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"191008",x"180f08",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"180f08",x"180f08",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1108",x"1b1008",x"191007",x"181007",x"191007",x"170e07",x"160f07",x"150e07",x"170f07",x"170f07",x"1b1108",x"1d1308",x"211508",x"261809",x"251709",x"261809",x"261809",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"150e07",x"150e07",x"432611",x"3b210e",x"3c230f",x"321d0d",x"341e0d",x"341d0d",x"371f0e",x"3c230f",x"3a210f",x"361f0e",x"361f0e",x"351e0e",x"341d0d",x"341d0d",x"351e0d",x"341d0d",x"341d0d",x"321c0c",x"351e0e",x"361f0e",x"39200f",x"361f0e",x"3b2210",x"39210f",x"39210f",x"3e2411",x"3a210f",x"3a210f",x"361f0e",x"361f0e",x"3a2210",x"3b2210",x"361f0f",x"3a210f",x"371f0e",x"3a200f",x"351d0d",x"381f0e",x"38200e",x"3c210f",x"3b220f",x"3a220f",x"3a210f",x"3e2411",x"3a2210",x"3c2311",x"422612",x"3d2310",x"3b2210",x"3d2310",x"3c2310",x"39200f",x"39200f",x"3c230f",x"3d2210",x"3c2310",x"3f2411",x"462914",x"4d2d16",x"3f2411",x"4b2c15",x"412612",x"351e0e",x"150e07",x"3b200e",x"3a210f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402716",x"402716",x"573c2b",x"563d2d",x"593b27",x"603b24",x"5d3c27",x"5e3c26",x"5f3e27",x"62412b",x"674228",x"603c25",x"613f28",x"5b3e2a",x"5b3e29",x"5d412f",x"5c402e",x"5a3c28",x"634531",x"5e3e28",x"64442e",x"644632",x"5f402d",x"644029",x"614029",x"5e3f2b",x"5a3e2b",x"563927",x"5c3c27",x"60412c",x"664734",x"634430",x"654835",x"5c402d",x"634431",x"5c3f2d",x"5d4232",x"5d402f",x"5e4333",x"604533",x"6b4b38",x"654530",x"6a4a34",x"6b4a35",x"694a35",x"6b4b36",x"6d4b36",x"6a4832",x"654734",x"684732",x"684934",x"61432e",x"634531",x"634633",x"63432f",x"61432e",x"5f3f2c",x"5c3e2c",x"583d2b",x"5a3d2b",x"5e3d27",x"5e412f",x"5c402d",x"5e422f",x"614431",x"674731",x"694934",x"6a4a34",x"644530",x"68452d",x"69452d",x"63412b",x"63402a",x"5e3f2b",x"5f3e28",x"5d3c27",x"603e27",x"613e27",x"613e27",x"624129",x"5a3c27",x"613f29",x"5c3a22",x"563621",x"503322",x"4a3221",x"5f3e28",x"513423",x"563825",x"5a3a26",x"573823",x"543827",x"563622",x"5b3923",x"5a3a26",x"523724",x"4f321f",x"4c3220",x"4a2f1d",x"4e301d",x"4f301c",x"4a2c19",x"51321c",x"53321c",x"4a2a16",x"4a2e1c",x"452b19",x"412919",x"482912",x"150e07",x"150e07",x"150e07",x"150e07",x"3e220f",x"150e07",x"1c130a",x"1e150c",x"1e140b",x"1e140b",x"1e150b",x"1f150c",x"1e140b",x"20160c",x"1e140b",x"1e140b",x"1e140b",x"1d140b",x"20160c",x"20160c",x"20150c",x"20160c",x"23180e",x"23180d",x"23180d",x"20160c",x"20160c",x"21160c",x"23180d",x"20150c",x"1f150b",x"1c1209",x"1f150b",x"1f150b",x"23180d",x"21170d",x"22170d",x"21170d",x"1e140b",x"21170d",x"21160d",x"21160d",x"21170d",x"22170d",x"23180e",x"20150c",x"24180e",x"23180e",x"23180e",x"23180d",x"20150c",x"20160c",x"20150c",x"23180d",x"23180e",x"23180d",x"20160c",x"20160c",x"23180d",x"23180e",x"20160c",x"20150c",x"1f150b",x"1c1209",x"1f150b",x"1f150b",x"23180d",x"24190f",x"23180d",x"20160b",x"20150b",x"22170d",x"22160d",x"21160d",x"21170d",x"22170d",x"21160c",x"20150c",x"21160d",x"21160c",x"21160c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1b1008",x"1b1108",x"1d1108",x"1d1208",x"1e1208",x"1f1309",x"201309",x"211409",x"221409",x"221409",x"221409",x"211409",x"201309",x"211409",x"211409",x"201409",x"1f1309",x"201309",x"1f1209",x"1f1309",x"1f1309",x"201309",x"201409",x"1f1309",x"201309",x"201409",x"201309",x"1e1208",x"201309",x"1f1309",x"1d1108",x"1e1208",x"1e1209",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"191008",x"191008",x"1b1108",x"180f08",x"180f08",x"180f07",x"191008",x"180f08",x"180f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1108",x"1a1108",x"1a1008",x"181007",x"170f07",x"180f07",x"170f07",x"181007",x"180f07",x"181007",x"191007",x"201508",x"231608",x"281909",x"281909",x"2a1b0a",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"231509",x"150e07",x"180f08",x"27160a",x"2a180b",x"201309",x"341d0c",x"361e0d",x"3c210f",x"3a200e",x"3c210f",x"391f0e",x"381e0d",x"371f0d",x"361e0d",x"391f0e",x"391f0e",x"3b210e",x"391f0e",x"391f0e",x"391f0d",x"2d1608",x"2a1408",x"2d1608",x"331b0b",x"371e0c",x"371e0d",x"371e0d",x"3a200d",x"381f0d",x"3a200e",x"3d220f",x"3e2310",x"3e2310",x"3d230f",x"3b210e",x"3d220f",x"3e230f",x"402410",x"3d220f",x"3f2410",x"402410",x"432611",x"442711",x"452812",x"432712",x"472913",x"442813",x"472913",x"452812",x"4b2b15",x"452813",x"462813",x"452813",x"472a14",x"4a2c15",x"432712",x"3f2310",x"3e220f",x"412411",x"452814",x"3f2410",x"150e07",x"412511",x"180f07",x"39200f",x"150e07",x"3d220f",x"3b220f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412716",x"412716",x"563a2a",x"5a3d2a",x"5e3e28",x"644028",x"654128",x"603b24",x"603c23",x"654128",x"64422c",x"5f3c24",x"5e3c25",x"573823",x"593924",x"563c2c",x"593c2a",x"5e4332",x"614736",x"583d2d",x"5e422f",x"583c29",x"5a3d2a",x"5d3e2a",x"543623",x"5a3d2b",x"5a3d2a",x"573c2a",x"614431",x"593b28",x"5a3e2c",x"5c402e",x"593d2d",x"543724",x"583b29",x"573825",x"573a27",x"543724",x"593a26",x"513222",x"452d21",x"492e22",x"503525",x"563927",x"5d402d",x"5c4030",x"5d412f",x"5c412f",x"604231",x"60412d",x"61422d",x"5c3d2a",x"5e4231",x"5c3e2a",x"5b3f2c",x"60412e",x"573d2c",x"543c2c",x"5c4230",x"5c402e",x"5d412f",x"5e4230",x"5d402e",x"5e402b",x"5f412e",x"5f4330",x"624430",x"61412c",x"60402a",x"61432d",x"61432d",x"644531",x"654530",x"67452e",x"603f2a",x"5d3d28",x"5b3a26",x"5d3924",x"644026",x"583621",x"543522",x"50321d",x"523420",x"503422",x"533624",x"543825",x"553825",x"543724",x"523624",x"523523",x"4e3220",x"4f3524",x"543621",x"5a3925",x"5e3c25",x"523520",x"51331f",x"422b1b",x"493020",x"4e301d",x"492d1a",x"4c2d18",x"4c2f1b",x"56341b",x"452915",x"4a2b18",x"432a1a",x"4a3120",x"452712",x"150e07",x"150e07",x"150e07",x"150e07",x"3f220f",x"150e07",x"1d140b",x"1c130a",x"1f150b",x"1d140b",x"1d140b",x"1e140b",x"20160c",x"1e140b",x"1d140b",x"20160c",x"1e140b",x"1d140b",x"20160c",x"1f150b",x"1f150b",x"21170d",x"20160c",x"21170d",x"24190f",x"21170d",x"24190f",x"21170d",x"24190e",x"22180e",x"22180e",x"21170d",x"21160c",x"22170d",x"24190f",x"24190f",x"21170d",x"20160c",x"20160c",x"1f150b",x"1f150b",x"20150c",x"20150c",x"21160d",x"20160c",x"20160c",x"23180d",x"23180d",x"23180e",x"23180d",x"23180d",x"1f150b",x"1f150b",x"24190e",x"23180e",x"24190e",x"21170d",x"21170d",x"24190e",x"24190e",x"24190e",x"251a0f",x"22180e",x"21170d",x"21160c",x"22170d",x"1e150c",x"22170d",x"21160d",x"20160c",x"20160c",x"1f150b",x"21160c",x"20150c",x"20150c",x"21160d",x"20160c",x"20160c",x"1d140b",x"20160c",x"20160c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"190f07",x"190f07",x"170f07",x"180f07",x"160e07",x"160f07",x"170f07",x"180f07",x"191008",x"1a1008",x"1a1008",x"1c1108",x"1c1108",x"1d1208",x"1e1209",x"201309",x"201309",x"211409",x"211409",x"211409",x"221409",x"211409",x"221409",x"211409",x"22140a",x"22150a",x"22150a",x"201409",x"1f1309",x"1e1208",x"1f1208",x"211409",x"1f1209",x"1f1309",x"211309",x"201309",x"25160a",x"211409",x"211409",x"221409",x"201309",x"24150a",x"201309",x"1f1309",x"1f1309",x"1e1209",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"201309",x"1b1108",x"1b1108",x"201309",x"1d1108",x"1b1108",x"1b1108",x"1a1008",x"1b1108",x"1a1008",x"1b1108",x"1f1309",x"1b1108",x"1d1108",x"1b1008",x"180f08",x"180f07",x"1a1008",x"180f07",x"180f07",x"180f07",x"1a1008",x"1a1008",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"191008",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160e07",x"170e07",x"190f07",x"1d1108",x"160f07",x"160f07",x"170f07",x"160f07",x"160f07",x"170f07",x"191008",x"170f07",x"191008",x"191008",x"160f07",x"160f07",x"160e07",x"1f1208",x"1b1108",x"160e07",x"160e07",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"190f08",x"150e07",x"150e07",x"160e07",x"1c1108",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1b1008",x"1b1108",x"190f08",x"191007",x"191007",x"180f07",x"180f07",x"1b1107",x"1b1108",x"1c1208",x"211409",x"201408",x"211508",x"2e1c0a",x"2b1a09",x"281809",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"201309",x"29180b",x"150e07",x"27160a",x"2e1a0c",x"2e1a0c",x"2c190b",x"28160a",x"2e1a0b",x"331c0d",x"371f0e",x"371f0e",x"371f0e",x"321d0d",x"3b2311",x"3b2210",x"3d2411",x"3f2512",x"38210f",x"3e2411",x"2d1a0c",x"3e2411",x"37200f",x"3c2311",x"3c2310",x"3b2310",x"3a2210",x"3f2511",x"3e2410",x"38200e",x"38200f",x"38200e",x"371f0e",x"381f0e",x"38200f",x"3a2210",x"37200f",x"3a220f",x"3b2210",x"412713",x"3f2512",x"3e2411",x"3e2410",x"3a2210",x"3a220f",x"3e2410",x"3a220f",x"412612",x"412612",x"3e2411",x"39200e",x"3c2210",x"422712",x"3d2310",x"3b210f",x"3f2512",x"3f2411",x"432712",x"3e2411",x"3e2411",x"3c2310",x"39200f",x"321c0c",x"2f1a0b",x"351e0d",x"351d0d",x"402310",x"150e07",x"442712",x"3c2310",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402616",x"402616",x"563c2c",x"66432c",x"61412b",x"603f2a",x"644127",x"6b4327",x"69432b",x"71472d",x"644129",x"623f28",x"644027",x"633f27",x"61412b",x"573a27",x"553b2a",x"5e4230",x"634532",x"644531",x"644532",x"5d4130",x"5a3d2c",x"604331",x"583d2c",x"5a3c29",x"5d3e2a",x"5c3c27",x"60432f",x"5a3e2c",x"624430",x"65452f",x"65432d",x"62432d",x"62422d",x"634530",x"624430",x"5f422e",x"62432f",x"6a4c37",x"6a4b36",x"644531",x"664530",x"6a4630",x"6b4830",x"6c4b35",x"6a4a35",x"644733",x"5f412e",x"654430",x"61412c",x"60422e",x"694830",x"64442f",x"644632",x"5d402c",x"5b3f2b",x"60432f",x"5c402d",x"5e4331",x"634633",x"61432e",x"62432f",x"60422e",x"5f412e",x"65442f",x"61422d",x"60402d",x"5c3f2d",x"62432e",x"61412a",x"583825",x"5e3f28",x"64432c",x"603f2b",x"60412b",x"62412a",x"63422a",x"64412a",x"613e28",x"543826",x"543523",x"533523",x"4f311f",x"51331e",x"503524",x"513421",x"523523",x"4e3320",x"4f3321",x"4b3121",x"472d1c",x"4e3220",x"573824",x"5a3924",x"513522",x"4f331f",x"462e1e",x"452d1d",x"472e1e",x"4a2e1c",x"4a2f1d",x"56341c",x"4d2f19",x"4c301c",x"50331f",x"4b2f1d",x"4e3220",x"4a2a12",x"150e07",x"150e07",x"150e07",x"150e07",x"412410",x"150e07",x"1f150b",x"1d140b",x"1f150b",x"1d140b",x"20150c",x"1f150b",x"1f150b",x"1f150b",x"1f150b",x"1f150b",x"1d130a",x"1f150b",x"20150c",x"20150b",x"1f150b",x"22170d",x"20160c",x"23180d",x"21160d",x"24180e",x"21160d",x"21160d",x"23180e",x"23180d",x"23170d",x"23180d",x"1f150b",x"1f150b",x"20160c",x"20150c",x"1f150b",x"1f150c",x"21160c",x"20160c",x"1f150b",x"22170d",x"20150c",x"1f150b",x"1f150b",x"21160c",x"21160c",x"21170c",x"1f150b",x"1f150b",x"22170d",x"22170d",x"22170d",x"22170d",x"23180d",x"23180d",x"23180e",x"24180e",x"24180e",x"23180e",x"23180d",x"23180d",x"23170d",x"20160c",x"1f150b",x"1f150c",x"20160c",x"20150c",x"1f150b",x"1f150c",x"1f150b",x"20160c",x"1f150b",x"20150c",x"20150c",x"1c130a",x"1f150b",x"1f150b",x"1f150b",x"1e140b",x"1e140b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341d0d",x"341d0d",x"150e07",x"201309",x"1a1008",x"170f07",x"1b1108",x"1a1108",x"1a1008",x"1c1108",x"1d1208",x"1d1209",x"1d1208",x"1f1309",x"201309",x"201309",x"221409",x"211409",x"22150a",x"221409",x"211309",x"211409",x"27170b",x"23150a",x"231409",x"23150a",x"221509",x"221509",x"22150a",x"22150a",x"27170b",x"231509",x"201309",x"1f1208",x"25150a",x"241509",x"26160a",x"27170a",x"27170a",x"27170b",x"29180b",x"26160a",x"27170a",x"241409",x"231409",x"25160a",x"28170b",x"25160a",x"26170b",x"26160b",x"24160a",x"1d1208",x"201309",x"24150a",x"23150a",x"24150a",x"26160a",x"24150a",x"24150a",x"26160a",x"211409",x"25160a",x"25160a",x"28180b",x"25160a",x"26160a",x"25160a",x"24150a",x"27170b",x"26160a",x"23150a",x"201309",x"1b1108",x"1b1108",x"231509",x"24150a",x"221409",x"24150a",x"1e1208",x"1a1008",x"191008",x"1c1108",x"1e1208",x"1f1309",x"201309",x"201309",x"29180b",x"25160a",x"221409",x"1f1309",x"1c1108",x"201309",x"201309",x"201309",x"201309",x"1e1209",x"27170b",x"22150a",x"201309",x"27170b",x"25160a",x"221409",x"211409",x"1f1309",x"27160a",x"201309",x"1d1108",x"1b1108",x"1d1208",x"1e1209",x"23150a",x"28180b",x"27170b",x"27170b",x"221409",x"1a1008",x"211409",x"26160a",x"1a1008",x"1c1108",x"150e07",x"191008",x"191008",x"1b1008",x"150e07",x"211409",x"1f1208",x"201309",x"191008",x"150e07",x"1f1309",x"1f1309",x"1c1108",x"211409",x"25160a",x"201309",x"221409",x"150e07",x"201309",x"1f1209",x"1e1209",x"29180b",x"211409",x"25160a",x"26160a",x"191008",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"241609",x"1e1208",x"231509",x"201308",x"1d1208",x"1b1108",x"1a1108",x"25160a",x"211409",x"231509",x"1b1108",x"23150a",x"28180a",x"36200d",x"2e1c0a",x"2c1a0a",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2f1a0c",x"150e07",x"221409",x"1d1108",x"211409",x"231409",x"231409",x"221409",x"211309",x"201208",x"231409",x"231409",x"211309",x"241509",x"241509",x"201309",x"251509",x"201309",x"251509",x"231509",x"28170a",x"221409",x"26160a",x"26160a",x"24150a",x"2e1b0d",x"301c0d",x"2d1b0d",x"2a190b",x"25150a",x"2a180b",x"27170b",x"25160a",x"2a190c",x"26160a",x"29180b",x"2c190c",x"25160a",x"26160a",x"2b190c",x"27170b",x"2c1a0c",x"2a180b",x"27160a",x"2a180b",x"25160a",x"2b190c",x"2d1a0c",x"301c0d",x"27170b",x"2f1b0d",x"28180b",x"2d1a0c",x"2b190b",x"2b190b",x"2b190b",x"2a190b",x"2d1a0c",x"311c0d",x"2e1b0d",x"27160a",x"211309",x"27160a",x"29170a",x"2c190b",x"3c210f",x"150e07",x"452712",x"3b2210",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432917",x"432917",x"533a2a",x"573b2a",x"583926",x"5f402d",x"5d3e2a",x"5f3c25",x"5d3c24",x"603d25",x"5e3b25",x"5a3b28",x"573b28",x"503624",x"593c2a",x"543928",x"503625",x"563a28",x"583d2b",x"5a3c2b",x"5d4231",x"5a4030",x"593f2d",x"543928",x"5c3f2e",x"5a4131",x"60412f",x"583c2b",x"5d4030",x"563d2e",x"583f2f",x"5c4231",x"584132",x"5d402e",x"5c4030",x"594030",x"583f30",x"594131",x"5b412f",x"614331",x"634836",x"654733",x"6a4e3b",x"6a4e3b",x"73513b",x"714f38",x"6d4c36",x"6c4c38",x"6a4b37",x"674b3a",x"6b4c38",x"6d4e38",x"694c39",x"674a35",x"684b38",x"644735",x"614634",x"5d4332",x"614632",x"644734",x"674833",x"5f4332",x"66452f",x"634734",x"644632",x"684733",x"644631",x"674530",x"604635",x"684934",x"654732",x"634430",x"644431",x"664632",x"684530",x"64442f",x"68452f",x"6c492f",x"5c3e29",x"573825",x"573824",x"563723",x"543522",x"4f3321",x"513625",x"533522",x"523523",x"543826",x"513523",x"422d1e",x"4e3422",x"4e3321",x"503320",x"462c1d",x"4e301d",x"4c301c",x"432b1b",x"442b1b",x"472d1d",x"412a1c",x"3a2518",x"472d1c",x"4f2f18",x"502f18",x"4e2f18",x"432a19",x"422917",x"3c271a",x"4b2913",x"150e07",x"150e07",x"150e07",x"150e07",x"432611",x"150e07",x"1d140b",x"1d130a",x"20160c",x"20160c",x"1f150b",x"1f150c",x"1f150b",x"1f150b",x"1f150b",x"1f150b",x"1c130a",x"1f150c",x"21160c",x"1f140b",x"22170d",x"22170d",x"22170d",x"21160d",x"24180e",x"24190f",x"21160d",x"20160c",x"23180e",x"23180d",x"20160d",x"20160c",x"23170d",x"21170c",x"1f150b",x"1f150b",x"1f150b",x"21160c",x"20150c",x"1f150b",x"1d140b",x"23180e",x"1f150b",x"1f150c",x"21160c",x"23180d",x"24180e",x"21160c",x"21160c",x"22170d",x"21160c",x"23170d",x"24180e",x"22170d",x"22170d",x"23180e",x"24180e",x"24190f",x"24180e",x"23180d",x"21160d",x"23180d",x"20160d",x"23180e",x"25190e",x"21170c",x"21160c",x"21160c",x"21170d",x"1f150b",x"20150c",x"1f150b",x"20160c",x"20160c",x"1f150b",x"1f150c",x"1f150b",x"1f150b",x"1f150b",x"1e150b",x"1e150b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"331e0e",x"331e0e",x"2f1b0d",x"2d1b0c",x"2c1a0c",x"23140a",x"201309",x"24160a",x"24150a",x"1b1108",x"1d1208",x"1d1208",x"1f1309",x"1e1209",x"211409",x"27170a",x"2b1a0c",x"29180b",x"2d1a0c",x"2d1b0d",x"2b190b",x"2f1c0d",x"2c1a0c",x"2d1b0c",x"2b190b",x"2c190c",x"27170b",x"24150a",x"2d1a0c",x"2c1a0c",x"311d0d",x"2a180b",x"29170a",x"231409",x"29170a",x"29180b",x"28170a",x"301b0c",x"2d1a0c",x"311c0d",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"2f1b0d",x"2f1b0c",x"2d1a0b",x"2e1a0c",x"29180b",x"2e1b0c",x"2e1b0c",x"2e1b0c",x"2a170b",x"26160a",x"2e1a0c",x"2d1a0c",x"27170a",x"2f1b0c",x"2c190c",x"29170b",x"29170b",x"29180b",x"2b190b",x"2b180b",x"2d1a0c",x"2e1a0c",x"2b190b",x"2f1b0c",x"2d1a0c",x"2d1a0c",x"2d1a0b",x"2b190b",x"28160a",x"231509",x"28160a",x"27160a",x"2c190b",x"2b180b",x"28160a",x"29170a",x"26160a",x"241509",x"28160a",x"241409",x"251509",x"261509",x"251509",x"201309",x"221409",x"241509",x"27160a",x"251509",x"241409",x"29170a",x"26160a",x"26160a",x"26160a",x"2d1a0b",x"2e1b0c",x"2f1b0d",x"2e1b0d",x"2c1a0c",x"331e0e",x"2f1b0d",x"2c1a0c",x"29180b",x"301c0d",x"2c1a0c",x"2d1a0c",x"2d1a0c",x"29180b",x"2f1b0c",x"2d1a0c",x"2d1a0c",x"321d0d",x"2f1b0d",x"301d0d",x"2d1a0b",x"2d1a0c",x"2e1b0c",x"27170a",x"2a190b",x"29190b",x"27170b",x"27170b",x"1c1108",x"150e07",x"29180b",x"211409",x"301c0d",x"23150a",x"2a190b",x"2b190c",x"28180b",x"2c1a0c",x"251509",x"28170a",x"27160a",x"2b180b",x"26160a",x"25160a",x"2b190b",x"2e1a0c",x"311c0c",x"29180b",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"211409",x"27170a",x"221509",x"29190b",x"241509",x"2a180a",x"2c1a0b",x"29180b",x"2a180a",x"301c0c",x"2b190b",x"2d1a0b",x"2b1a0b",x"301c0b",x"38210d",x"38200e",x"2f1c0a",x"301d0b",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"170f07",x"321d0d",x"150e07",x"351e0d",x"351d0d",x"331c0c",x"371e0d",x"351d0c",x"331b0b",x"351d0c",x"341c0b",x"361d0c",x"371d0c",x"341c0c",x"361d0c",x"3c200e",x"3a200e",x"3c210f",x"3e230f",x"3d220f",x"3e2310",x"3f2310",x"432612",x"422611",x"402410",x"412511",x"442712",x"432612",x"462913",x"452813",x"422612",x"442713",x"442713",x"442913",x"472a14",x"3f2411",x"412511",x"3f2410",x"3d220f",x"381f0d",x"3f2410",x"432611",x"402410",x"3c210e",x"3b200e",x"3b200e",x"3a1f0e",x"3b200e",x"3e220f",x"412410",x"442712",x"472a14",x"482a14",x"492b15",x"472a15",x"442712",x"3e2210",x"402310",x"432611",x"492b15",x"472914",x"492b15",x"402511",x"452813",x"442713",x"472914",x"432712",x"150e07",x"422511",x"37200f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442815",x"442815",x"5c402d",x"5a3d2a",x"5f412f",x"66442e",x"634028",x"634029",x"633f27",x"5c3a26",x"5d3e2a",x"593824",x"543624",x"503726",x"553724",x"593a27",x"583824",x"5b3b27",x"593f2e",x"5d3e2a",x"604230",x"5d412f",x"573e2d",x"543c2d",x"563b2b",x"53392a",x"563929",x"523627",x"553a29",x"573c2c",x"51392a",x"594030",x"5d4332",x"5d4332",x"5f4536",x"5a3e2d",x"5e4331",x"5c412f",x"654734",x"664733",x"634836",x"62442f",x"6a4d3b",x"684b38",x"634836",x"6b4b35",x"694832",x"654936",x"654733",x"614431",x"694a35",x"6b4b36",x"674630",x"644733",x"664a38",x"614736",x"5f4332",x"594131",x"664834",x"614634",x"644635",x"5b4131",x"583f2f",x"5f4332",x"614331",x"5a3f2f",x"5c402f",x"664632",x"654733",x"6b4a34",x"6a4932",x"664631",x"66432d",x"62432f",x"62422e",x"613f29",x"6a4630",x"69452c",x"68472f",x"61402b",x"624029",x"5f3f29",x"5e3f2a",x"5c3d29",x"593c29",x"5b3d28",x"5d3e29",x"61422b",x"5a3c27",x"523824",x"443022",x"4d3522",x"4c3321",x"523521",x"4f3422",x"4e321f",x"513523",x"472d1b",x"422c1c",x"472e1d",x"472e1d",x"4a2e18",x"59371e",x"5d3a20",x"52331d",x"4a2c18",x"412a1c",x"472f1f",x"4d2c14",x"150e07",x"150e07",x"150e07",x"150e07",x"432510",x"150e07",x"22170d",x"20160c",x"24180e",x"21170d",x"21170d",x"23180d",x"21160d",x"21160d",x"1f150b",x"20150c",x"20160c",x"22170d",x"20160c",x"24190e",x"24180e",x"261a0f",x"20160c",x"22170d",x"23180e",x"21160d",x"24190f",x"281c10",x"23180e",x"23180e",x"251a0f",x"22170d",x"22170d",x"22170d",x"21160c",x"21160c",x"23180d",x"23180d",x"291c11",x"23180e",x"261a0f",x"24190e",x"271b10",x"20160c",x"23180e",x"23180e",x"23180d",x"22170d",x"251a0f",x"22170d",x"25190e",x"24190e",x"271b10",x"23180d",x"22170d",x"22170d",x"23180e",x"2b1e12",x"271b10",x"281c10",x"261a0f",x"25190f",x"23180e",x"24180e",x"24190e",x"1f150b",x"23180d",x"21160c",x"23180d",x"23180d",x"22170d",x"23180e",x"24180e",x"261a10",x"271b10",x"20160c",x"21160d",x"20160c",x"21160c",x"20160c",x"20160c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200f",x"38200f",x"3a2110",x"2f1c0d",x"2e1b0c",x"341d0e",x"2c1a0b",x"2c1a0b",x"1a1108",x"1a1008",x"1b1108",x"1d1108",x"1f1309",x"241509",x"261509",x"281709",x"27160a",x"29170a",x"29170a",x"2d190b",x"301b0c",x"331d0e",x"341f0e",x"341f0e",x"331e0e",x"331d0d",x"29170a",x"28170a",x"2c190b",x"311d0d",x"331d0e",x"2f1c0d",x"301c0d",x"2e1b0c",x"2f1b0c",x"331e0e",x"341e0e",x"351f0e",x"38210f",x"382110",x"382211",x"372110",x"3a2311",x"3e2512",x"382210",x"3b2311",x"36200f",x"331d0e",x"341e0e",x"361f0f",x"38210f",x"38210f",x"341f0f",x"37210f",x"331e0e",x"331e0e",x"37200f",x"361f0f",x"301b0c",x"2f1b0c",x"2f1b0c",x"29180b",x"341e0e",x"311c0d",x"311c0c",x"301b0c",x"2d190b",x"2f1a0b",x"2e1a0b",x"311c0c",x"321c0d",x"331d0c",x"2a180a",x"321c0c",x"301b0c",x"301b0b",x"2c190b",x"2e1a0b",x"2c180b",x"2a170a",x"281509",x"281609",x"261509",x"271609",x"2a170a",x"28160a",x"2b180a",x"261509",x"29170a",x"29170a",x"2e1a0b",x"301b0c",x"2f1b0c",x"2d1a0b",x"2d1a0c",x"321c0d",x"311c0d",x"321c0d",x"2f1b0c",x"341e0e",x"321d0d",x"341e0e",x"321d0d",x"321d0d",x"301c0d",x"361f0f",x"311d0e",x"341e0e",x"331d0d",x"331d0d",x"301b0c",x"2f1a0c",x"321c0c",x"351e0d",x"341d0d",x"321c0c",x"2e190b",x"2f1a0b",x"2e190b",x"2b180a",x"2c180b",x"2b180b",x"2a180b",x"2c1a0c",x"211409",x"1c1108",x"150e07",x"29180b",x"27160a",x"29170a",x"2d190b",x"341e0e",x"2c1a0c",x"39210f",x"38210f",x"311c0d",x"341e0e",x"351e0e",x"2e1b0d",x"321d0d",x"38200f",x"38210f",x"341f0f",x"180f08",x"191008",x"1a1108",x"1c1108",x"29190c",x"2d1b0c",x"2a180b",x"321d0d",x"301c0d",x"2e1b0c",x"331e0e",x"321d0d",x"35200f",x"331e0e",x"351f0e",x"351f0f",x"321d0d",x"3b220f",x"3d240e",x"40260f",x"422711",x"311e0b",x"2b1a09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"191008",x"2f1b0c",x"150e07",x"321d0e",x"2b190c",x"26160a",x"25150a",x"27160a",x"26160a",x"29180b",x"2d1a0b",x"2b190b",x"321c0d",x"2e1b0c",x"301c0c",x"2d1a0b",x"2d1a0b",x"29180b",x"2b190b",x"29180b",x"29170b",x"2e1a0b",x"2e1b0c",x"2d190b",x"27160a",x"2c190b",x"311c0d",x"29180b",x"301c0d",x"2e1a0c",x"2c190b",x"2f1c0d",x"2d1a0c",x"301c0d",x"2d1a0c",x"2e1b0c",x"2e1a0b",x"2d190b",x"2d190b",x"2c190b",x"301b0c",x"2c190b",x"2f1b0c",x"311c0d",x"341e0d",x"341e0e",x"311c0d",x"361f0e",x"311c0c",x"351e0d",x"39210f",x"37200f",x"321d0d",x"341d0d",x"311b0c",x"301b0c",x"301b0c",x"36200f",x"38210f",x"3a2210",x"361f0e",x"301b0c",x"331d0d",x"311d0d",x"321d0d",x"311c0d",x"432612",x"150e07",x"472913",x"3d2411",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472a17",x"472a17",x"553d2c",x"634734",x"64412b",x"65442e",x"68442d",x"714a2e",x"6e472d",x"6f4a2f",x"654229",x"5b3c26",x"5e3d28",x"5e3d28",x"66432c",x"5e412e",x"60412e",x"63432d",x"694731",x"664630",x"684630",x"66452f",x"65442e",x"614533",x"60412d",x"5d3f2a",x"5e402d",x"674732",x"64422d",x"66422c",x"61412a",x"60412d",x"603e29",x"5e3f2a",x"5b3e2b",x"5c3e2a",x"533827",x"513726",x"543827",x"5b3d29",x"583a27",x"583b29",x"5b3d29",x"5b3b25",x"64432d",x"67452f",x"67462f",x"5d3f2b",x"5a3d2a",x"63432e",x"67452f",x"65432e",x"5f412d",x"5c3e2c",x"5d3f2d",x"5f3f2d",x"5f402d",x"60402b",x"624532",x"5f412e",x"614534",x"654632",x"664530",x"65442f",x"6a4934",x"664632",x"694731",x"694834",x"674630",x"68452f",x"66442d",x"6a4731",x"654634",x"613f2b",x"66432b",x"6c4730",x"6c4831",x"66432d",x"62402a",x"593c29",x"60402a",x"62422c",x"623f27",x"573925",x"593a26",x"5a3b26",x"583824",x"5a3923",x"5a3b26",x"503523",x"483020",x"4a3223",x"432c1c",x"493121",x"4e311e",x"4f3320",x"4b311e",x"5a3a23",x"4f3320",x"472d1c",x"482f1d",x"422916",x"4c2e1a",x"51311a",x"4f301b",x"482f1e",x"442b19",x"412c1f",x"4b2b13",x"150e07",x"150e07",x"150e07",x"150e07",x"381d0c",x"150e07",x"21170d",x"24190e",x"24190f",x"21170d",x"1e140b",x"22170d",x"1f150b",x"20150c",x"21160c",x"22170d",x"23180d",x"20160c",x"21160c",x"26190e",x"25190e",x"2b1d11",x"23180d",x"23180d",x"281c10",x"22170d",x"24180e",x"1c1208",x"1d1309",x"21160c",x"21170d",x"281c10",x"24190e",x"261a0f",x"281b10",x"291c10",x"25190f",x"2a1d11",x"24190e",x"261a0f",x"2a1d12",x"261a0f",x"251a0f",x"281b10",x"24180e",x"281b10",x"261a0e",x"271b0f",x"25190f",x"25190e",x"23170d",x"271b0f",x"281c10",x"271b10",x"281c10",x"21160c",x"23180d",x"25190e",x"26190f",x"1c1208",x"1f140a",x"271b0f",x"291c10",x"281c10",x"22170d",x"281b10",x"24190e",x"251a0f",x"251a0f",x"24190e",x"21160d",x"2a1d11",x"24190f",x"24190e",x"251a0f",x"22170d",x"271b0f",x"22170d",x"1f150b",x"20160c",x"20160c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"37200f",x"37200f",x"36200e",x"2f1c0c",x"37200e",x"311d0c",x"311c0b",x"180f07",x"190f08",x"1a1008",x"1b1108",x"26160a",x"27170a",x"311d0c",x"321d0c",x"301c0d",x"2e1a0c",x"321d0d",x"311b0c",x"341e0e",x"341e0e",x"351f0e",x"331d0e",x"351f0e",x"331d0d",x"321c0c",x"2f1a0c",x"331d0d",x"36200f",x"3b2211",x"361f0f",x"341d0d",x"341e0d",x"36200e",x"321d0d",x"341e0e",x"351f0e",x"341e0e",x"321c0d",x"361e0e",x"361f0e",x"392110",x"361f0e",x"37200f",x"351f0e",x"38200f",x"351e0e",x"361e0e",x"38210f",x"3b2210",x"3c2311",x"3d2411",x"3e2512",x"3a2210",x"3a2210",x"37200f",x"38200f",x"392110",x"38200f",x"38200f",x"3a2210",x"3d2411",x"3b2311",x"3a2311",x"3a2311",x"3c2411",x"392210",x"392110",x"38200f",x"3c2311",x"3b2210",x"311c0d",x"2f1b0c",x"3c2210",x"38210f",x"39210f",x"39210f",x"39210f",x"38200f",x"341e0d",x"351e0d",x"351e0d",x"361e0d",x"371f0e",x"361f0e",x"361f0e",x"341e0e",x"331d0d",x"2d1a0c",x"341e0e",x"321d0d",x"351e0e",x"321d0d",x"301c0c",x"311c0d",x"2f1b0c",x"341d0d",x"361e0d",x"351e0d",x"351f0e",x"37200f",x"321d0d",x"351e0e",x"361f0e",x"351f0e",x"38210f",x"331e0d",x"38200f",x"2f1b0c",x"331c0c",x"301a0c",x"321c0c",x"351e0d",x"351e0d",x"341d0d",x"371f0e",x"3a200f",x"38200f",x"38210f",x"38200e",x"331d0d",x"341e0e",x"321d0d",x"331f0d",x"301c0c",x"301c0d",x"201408",x"27160a",x"28170a",x"331d0d",x"2f1c0d",x"301d0d",x"3a2110",x"311c0d",x"351e0d",x"351e0e",x"351e0e",x"361f0e",x"371f0e",x"402511",x"351e0e",x"341d0d",x"160f07",x"170f07",x"180f07",x"191008",x"201309",x"2d1a0c",x"2f1b0c",x"2c190b",x"2e1b0c",x"311d0e",x"37200f",x"3b2311",x"3d2411",x"392210",x"3c2411",x"38200f",x"3a2110",x"3d2411",x"402610",x"472b11",x"472b12",x"3f260e",x"311d0b",x"301c0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1b1108",x"2a180b",x"150e07",x"2e1b0c",x"351e0e",x"2d190b",x"2f1a0b",x"331c0c",x"351d0d",x"381f0e",x"2f1a0b",x"331c0c",x"321c0c",x"341d0d",x"351d0d",x"331d0d",x"341e0d",x"351e0e",x"37200f",x"38210f",x"341e0d",x"3a210f",x"371f0e",x"351e0d",x"361f0d",x"341d0d",x"361e0d",x"301a0b",x"351d0d",x"38200e",x"361e0e",x"361f0e",x"321c0d",x"351e0d",x"321c0c",x"3a210f",x"371f0e",x"321c0c",x"341d0d",x"311c0c",x"351d0d",x"341d0d",x"351e0d",x"361f0e",x"38200e",x"39200e",x"321c0d",x"351d0d",x"361e0d",x"311b0b",x"311b0c",x"351d0d",x"361e0d",x"321c0c",x"311b0c",x"331c0c",x"321c0c",x"371f0e",x"38200f",x"331d0d",x"331c0d",x"341d0d",x"311c0c",x"321c0c",x"2e190b",x"2f190b",x"381e0d",x"150e07",x"3e220f",x"37200f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472b17",x"472b17",x"5c4331",x"563b29",x"61412d",x"69452d",x"6c472f",x"6d472d",x"6b452d",x"65412a",x"613e27",x"61412a",x"61412b",x"61422d",x"674630",x"694c38",x"5e3f2c",x"664630",x"65442f",x"654531",x"674731",x"63422a",x"5a3b26",x"5b3b28",x"553928",x"553927",x"5f402d",x"62422f",x"634330",x"5b3f2d",x"614230",x"5d4130",x"5e4230",x"5f412e",x"5d3e2b",x"5c4332",x"59402f",x"564031",x"614531",x"624431",x"573e2e",x"563e2f",x"563d2d",x"5b3f2d",x"583d2d",x"563b2b",x"5b3f2d",x"5d402d",x"573e2d",x"593e2c",x"5c4231",x"604532",x"644734",x"624836",x"5e4333",x"614634",x"634534",x"624432",x"624432",x"684836",x"644532",x"634532",x"654734",x"654734",x"654734",x"62432e",x"5d3f2c",x"624331",x"5e402f",x"5c412f",x"5b3f2d",x"5f412f",x"5b4131",x"604332",x"61422e",x"644531",x"644633",x"60432f",x"5e3f2c",x"5a3c29",x"563a29",x"553928",x"4d3121",x"533625",x"523626",x"503321",x"563927",x"563826",x"543623",x"533521",x"4f3221",x"4d3424",x"503524",x"4d3321",x"513623",x"563521",x"553621",x"54331d",x"4d301b",x"4d2f1b",x"4d321f",x"492c18",x"50331e",x"59361c",x"452b17",x"472e1d",x"4c2f1d",x"4c3323",x"4a2812",x"150e07",x"150e07",x"150e07",x"150e07",x"3c1f0d",x"150e07",x"23180e",x"2c1e12",x"261a0f",x"25190e",x"20160c",x"23180d",x"24190e",x"21170d",x"23170d",x"20150c",x"22170d",x"271b0f",x"25190e",x"291c10",x"251a0f",x"251a0f",x"281c10",x"25190e",x"2a1d11",x"23180d",x"291b0f",x"271a0f",x"261a0f",x"25190e",x"291c10",x"291c10",x"2d1f12",x"2a1d11",x"251a0f",x"2b1e12",x"291c10",x"291d11",x"291d11",x"261a0f",x"261a0f",x"281c10",x"2a1d11",x"2d1f12",x"2e2013",x"2c1e12",x"2a1d11",x"2c1e11",x"2c1e11",x"291c11",x"2c1e12",x"2b1d11",x"251a0f",x"291c10",x"2e2013",x"2c1e12",x"2c1e12",x"2a1d11",x"22170d",x"281c10",x"2d2013",x"281b10",x"291c10",x"22170d",x"271b10",x"2a1d11",x"251a0f",x"251a0f",x"291c10",x"291d11",x"291d11",x"2a1d11",x"2a1d11",x"25190e",x"20150c",x"23180e",x"24190e",x"21170c",x"1d140b",x"24180d",x"24180d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"37200e",x"37200e",x"331c0d",x"351d0d",x"2e1a0b",x"341d0d",x"2e1a0b",x"1e1208",x"191008",x"1a1008",x"211309",x"271609",x"311d0c",x"311d0b",x"2d1a0b",x"311c0c",x"2e1a0b",x"2d190b",x"331c0d",x"2d190b",x"2d190b",x"311b0c",x"2f1a0b",x"2e1a0b",x"2f1a0b",x"2e1a0b",x"2e190b",x"311b0c",x"311c0c",x"311c0d",x"361e0e",x"311c0c",x"311b0c",x"2e1a0b",x"2e190b",x"2b170a",x"2f190b",x"2f1a0b",x"311b0c",x"311b0c",x"361d0d",x"351d0d",x"351e0d",x"37200f",x"38210f",x"37200e",x"3b2210",x"38200f",x"371f0e",x"361f0e",x"3a210f",x"36200e",x"351f0e",x"3a2210",x"3a2110",x"38200f",x"3d2411",x"3c2311",x"37200f",x"361f0f",x"3e2411",x"392210",x"3d2411",x"38210f",x"3c2310",x"3c2311",x"38210f",x"3a2210",x"3a2210",x"3b2210",x"3d2411",x"38200f",x"361f0e",x"361f0f",x"361f0e",x"39210f",x"39210f",x"331d0c",x"311b0b",x"2f190b",x"2f1a0b",x"2f1a0b",x"341d0d",x"311b0c",x"311b0c",x"321c0c",x"311b0c",x"321c0c",x"311c0d",x"341e0e",x"331d0e",x"38200f",x"361f0e",x"341e0e",x"351e0e",x"341d0d",x"321c0c",x"361e0d",x"341d0d",x"311b0c",x"2f1a0b",x"331d0d",x"311c0c",x"351e0e",x"361f0e",x"371f0e",x"321c0c",x"311c0c",x"301b0c",x"311c0c",x"311c0c",x"2f1a0c",x"361e0e",x"371f0d",x"371f0e",x"361f0d",x"301b0c",x"331d0d",x"361e0e",x"351d0d",x"351d0d",x"341d0c",x"331d0c",x"2f1b0b",x"2b1a0b",x"281709",x"231509",x"150e07",x"27160a",x"2c190b",x"321c0d",x"321d0d",x"341d0c",x"2d190b",x"2f1a0b",x"311b0c",x"2f1a0b",x"2c170a",x"2d190a",x"301a0b",x"351c0c",x"341d0c",x"160e07",x"170f07",x"170f07",x"1d1208",x"2e1b0c",x"2c1a0c",x"2e1b0c",x"341e0e",x"301c0d",x"301c0c",x"331c0d",x"361f0e",x"341e0e",x"3a210f",x"39220f",x"37200e",x"3c2310",x"402711",x"442912",x"4a2d13",x"4a2c13",x"36210b",x"36200b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"331d0d",x"150e07",x"231409",x"2e190b",x"180f07",x"321c0c",x"381e0d",x"371d0c",x"341c0c",x"351c0c",x"361d0c",x"361d0c",x"381e0d",x"3a200d",x"3c210f",x"412511",x"412511",x"452813",x"432712",x"452813",x"432713",x"3c2311",x"412612",x"3f2410",x"422611",x"402411",x"3e230f",x"3e220f",x"3f230f",x"3e220f",x"432511",x"422611",x"422511",x"3f2310",x"402410",x"402410",x"3f2310",x"3a200e",x"3c210f",x"3b200e",x"3c210f",x"3e220f",x"442712",x"442711",x"412511",x"422611",x"412411",x"462812",x"402410",x"422611",x"3f2310",x"402310",x"3d210f",x"3d210f",x"3e220f",x"3d210f",x"422611",x"452813",x"422712",x"432612",x"3e220f",x"3b200e",x"150e07",x"39200e",x"231409",x"321c0c",x"150e07",x"412410",x"39210f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452916",x"452916",x"513c2d",x"533828",x"573a27",x"61412c",x"5f3e28",x"66422c",x"674229",x"68442b",x"613f28",x"614029",x"60412c",x"614431",x"62432e",x"5b3e2c",x"5d402e",x"604330",x"61412d",x"61422d",x"60412c",x"573b29",x"5c3e2c",x"5d3d2b",x"583a28",x"533728",x"553827",x"583a28",x"5a3b2a",x"583e2f",x"583a29",x"563d2d",x"593d2c",x"593d2a",x"5f412d",x"60422d",x"593d2a",x"543d2d",x"553f30",x"5a3f2d",x"583f2d",x"573d2c",x"4d382a",x"573e2d",x"563d2d",x"583e2d",x"573c2a",x"503829",x"513a2b",x"583e2d",x"5a4030",x"5b4131",x"604431",x"624533",x"573f30",x"5b4130",x"5e4332",x"5a3f2f",x"634633",x"654835",x"684a36",x"674a36",x"674631",x"674833",x"664631",x"694834",x"674735",x"674835",x"674733",x"654532",x"664835",x"684936",x"654734",x"634330",x"64432d",x"674733",x"664630",x"5f412c",x"634531",x"573d2c",x"5a3e2c",x"5f412f",x"5b3f2d",x"60412e",x"5f402c",x"5e3d29",x"5b3b26",x"593b28",x"523524",x"503423",x"4f3321",x"482f1e",x"452e1f",x"472f20",x"4c311f",x"58341e",x"56341f",x"50311d",x"4a2e1d",x"342118",x"321f15",x"3c2516",x"442917",x"452917",x"462c1a",x"412a1b",x"3f2718",x"442f20",x"492912",x"150e07",x"150e07",x"150e07",x"150e07",x"3b1f0d",x"150e07",x"23180d",x"24190e",x"22170d",x"281c10",x"23180d",x"23180d",x"261a0f",x"23180e",x"251a0f",x"251a0f",x"291c11",x"25190e",x"24180e",x"271b10",x"291c10",x"25190e",x"291c11",x"261a0f",x"2b1e12",x"2d1f12",x"2a1d11",x"2d1f12",x"291c10",x"2a1d11",x"2b1d11",x"251a0f",x"2d1f12",x"2e2013",x"2b1e12",x"2d2013",x"291c11",x"281b10",x"2a1d11",x"24190e",x"271b10",x"2a1d11",x"2a1d11",x"281b10",x"291c10",x"2d2013",x"2d1f12",x"2d1f13",x"291c11",x"281c10",x"2d1f12",x"291d11",x"2b1e12",x"2c1e12",x"2b1e12",x"2b1e12",x"291d11",x"291c10",x"2a1d11",x"2b1d11",x"2b1d11",x"2c1e12",x"291c10",x"291c10",x"2b1d11",x"291c10",x"291c11",x"2d2013",x"271b10",x"24190e",x"281c10",x"271b10",x"291c11",x"2a1d11",x"281c10",x"25190e",x"23180e",x"291d11",x"23180d",x"24190e",x"24190e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351e0d",x"351e0d",x"351d0d",x"2d1a0b",x"2f1b0c",x"311c0c",x"191007",x"180f07",x"190f08",x"1c1208",x"221408",x"2e1b0b",x"331d0c",x"321d0c",x"3a220d",x"321d0c",x"311c0c",x"2f1b0c",x"2f1b0c",x"331d0d",x"321c0d",x"331c0d",x"301b0c",x"321c0c",x"331c0c",x"2f1a0b",x"321c0d",x"311c0c",x"341d0e",x"3a2210",x"351f0e",x"371f0e",x"301b0c",x"321c0c",x"331c0d",x"321c0c",x"341d0d",x"351e0d",x"351e0e",x"321c0c",x"2e1a0b",x"301a0b",x"311b0c",x"321c0c",x"311b0c",x"301a0b",x"331c0c",x"331c0c",x"321c0c",x"2e1a0b",x"301b0c",x"2e1a0b",x"221107",x"241208",x"2d190b",x"331c0c",x"321c0c",x"331c0d",x"351e0d",x"321c0d",x"331d0d",x"341e0d",x"361f0e",x"38200f",x"38210f",x"3a2210",x"38210f",x"3a2210",x"38210f",x"37200f",x"38200e",x"2e1a0b",x"351e0d",x"341d0d",x"361f0d",x"3a210f",x"321c0c",x"2f190b",x"331c0c",x"2e190b",x"2c180a",x"271509",x"2d180a",x"2d180a",x"2f190b",x"2d180a",x"2e190b",x"2d190b",x"2f1b0c",x"2f1b0c",x"341e0e",x"37200f",x"321d0d",x"341e0e",x"38210f",x"38200f",x"341e0e",x"341e0d",x"341e0e",x"321c0d",x"331c0d",x"341d0d",x"331d0d",x"351e0d",x"331d0d",x"341e0d",x"2f1b0c",x"301b0c",x"301b0c",x"321c0d",x"2e190b",x"2d190b",x"2f1a0b",x"311b0c",x"38200e",x"381f0e",x"38200e",x"351f0e",x"371f0e",x"3c230f",x"361f0d",x"311c0c",x"3a220e",x"2b190a",x"2e1b0b",x"2d1b0a",x"251609",x"1d1208",x"27160a",x"2e1a0b",x"38210f",x"351f0d",x"3c2310",x"371f0e",x"331c0c",x"331c0d",x"341d0d",x"361e0d",x"361e0d",x"38200e",x"3b220f",x"160e07",x"160e07",x"160f07",x"170f07",x"1f1208",x"261509",x"2b180a",x"2c190b",x"2d190b",x"2f1a0c",x"311b0c",x"2d190b",x"2f1b0b",x"251408",x"241107",x"2f190b",x"331d0c",x"3a210e",x"3f250f",x"422710",x"492c11",x"40280d",x"39240b",x"36210b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"351e0e",x"150e07",x"150e07",x"3b1f0d",x"3f2310",x"3d2310",x"3d220f",x"391f0e",x"3b210f",x"3b210e",x"381f0e",x"371e0d",x"321c0c",x"341c0c",x"351d0d",x"361f0e",x"371f0e",x"361e0e",x"351d0d",x"351e0d",x"351e0d",x"351f0e",x"37200f",x"371f0e",x"381f0e",x"341d0d",x"331c0c",x"301b0b",x"391f0e",x"371e0d",x"351d0d",x"321b0c",x"321c0b",x"321b0c",x"351d0d",x"351d0d",x"331c0c",x"321b0c",x"351d0d",x"371f0d",x"341d0d",x"371e0e",x"3b210f",x"381f0e",x"38200f",x"39200e",x"3b210f",x"3a200f",x"3c210f",x"2f1b0c",x"3c210f",x"39200e",x"381f0e",x"3c220f",x"3f2411",x"422612",x"3e2411",x"3f2411",x"3d230f",x"3b210f",x"402511",x"472913",x"412411",x"432510",x"2d190b",x"2d1a0b",x"150e07",x"3e220f",x"38200e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482b18",x"482b18",x"513b2c",x"583c2b",x"5a3f2e",x"65432d",x"5b3b25",x"634029",x"644028",x"5d3d26",x"593a26",x"563b2a",x"4e3526",x"543a2b",x"583e2d",x"4d3527",x"4e3526",x"573f2f",x"543929",x"543929",x"5a3a26",x"543828",x"5e3d29",x"633f28",x"603e27",x"5d3b26",x"5d3e2b",x"623f29",x"5c3c27",x"5f3f2d",x"543927",x"5b3d2b",x"583b2b",x"573a28",x"583c2b",x"5b3e2c",x"553a29",x"543b2b",x"563a28",x"563b28",x"5c3f2c",x"5a3f2e",x"584030",x"573c2b",x"523a2a",x"573c2b",x"4f392c",x"533b2b",x"513b2c",x"4f3a2b",x"4b382c",x"503c2f",x"563d2d",x"5b4231",x"574234",x"594132",x"5b4536",x"5e4433",x"614533",x"634634",x"654a38",x"684a38",x"614735",x"664937",x"654936",x"654733",x"624330",x"644531",x"624532",x"674a37",x"61402d",x"684632",x"704e39",x"6a4933",x"6c4832",x"674732",x"654734",x"5a3c2a",x"5b4130",x"5d4433",x"5b4131",x"614534",x"5b4130",x"5d3d2a",x"573b29",x"553827",x"583926",x"5a3b27",x"573724",x"5a3a26",x"513522",x"4f3321",x"4e321f",x"513524",x"4c3221",x"583723",x"4f3220",x"583722",x"50311d",x"472c19",x"452c1d",x"422919",x"392415",x"3d2415",x"402a1c",x"482e1d",x"3d2719",x"4b3222",x"4c2b14",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200e",x"150e07",x"251a0f",x"23180e",x"251a0f",x"271b10",x"2d1f13",x"24190f",x"271b10",x"24190f",x"261a0f",x"271b10",x"281c11",x"2d2014",x"2c1f13",x"2a1d11",x"2c1f13",x"2e2013",x"291c11",x"25190e",x"2f2114",x"281c10",x"281b10",x"291c10",x"261a0f",x"281c10",x"2a1d11",x"291c10",x"271a0f",x"291c10",x"312214",x"291c10",x"291c10",x"291c10",x"291c10",x"291c11",x"2b1d11",x"2c1f13",x"2d1f13",x"312316",x"2b1e12",x"2c1f13",x"2e2013",x"2d1f13",x"302215",x"2d2014",x"302215",x"2c1e12",x"2e2114",x"302114",x"2b1e12",x"2a1d11",x"2d2013",x"2c1f12",x"2a1d11",x"2b1d11",x"281c10",x"281c10",x"261a0f",x"291c10",x"271a0f",x"281b0f",x"2a1d11",x"2b1e11",x"2b1d11",x"2b1d11",x"2b1d11",x"291d11",x"251a0f",x"271b10",x"2a1e12",x"271b10",x"24190f",x"2a1d11",x"24180e",x"271b0f",x"271b0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0b",x"311c0b",x"2c180a",x"271609",x"29160a",x"261509",x"180f07",x"170f07",x"1c1107",x"201408",x"26160a",x"2b190b",x"2f1b0b",x"37210d",x"36200d",x"2f1b0c",x"331d0d",x"2f1b0c",x"2f1a0c",x"2f1b0c",x"2e1a0b",x"311b0c",x"301b0c",x"311b0c",x"361f0e",x"38200f",x"341e0e",x"341f0e",x"341e0e",x"331d0d",x"321c0d",x"351e0d",x"331d0d",x"301b0c",x"311b0c",x"331c0c",x"2f1b0c",x"2e1a0b",x"2e190b",x"2d190b",x"311b0c",x"301b0c",x"341d0d",x"301a0c",x"331d0d",x"311d0d",x"361f0e",x"311c0c",x"311b0c",x"331c0d",x"2e1a0b",x"2c190b",x"2d190b",x"2d190b",x"2a180b",x"2d190b",x"2a180a",x"2c190b",x"311b0c",x"321c0d",x"301c0c",x"311c0d",x"301c0c",x"2f1b0c",x"2e1a0c",x"2d190b",x"2c190b",x"331c0c",x"311b0c",x"311c0d",x"2d190b",x"2a170a",x"2d190b",x"2c190b",x"2d190b",x"2e190b",x"2e190a",x"301a0b",x"331d0d",x"311c0d",x"2d1a0b",x"28170a",x"2c190b",x"2f1a0c",x"2d190b",x"2c190b",x"2a180b",x"2c190b",x"2b190b",x"2b190b",x"2e1a0b",x"2e1a0c",x"2d190b",x"2e1a0c",x"301c0c",x"341e0e",x"331d0d",x"2b190b",x"2c190b",x"2e1a0b",x"2b180a",x"2d190a",x"311b0c",x"301b0c",x"2b180a",x"2d180a",x"29170a",x"28160a",x"2d190b",x"28170a",x"2a170a",x"2f1a0b",x"321c0c",x"2c190b",x"2f1a0c",x"321c0c",x"331d0d",x"2a180b",x"361f0d",x"361e0e",x"331d0d",x"39210e",x"39210d",x"3d240e",x"2f1d0b",x"2a190a",x"221509",x"221509",x"351f0d",x"311d0d",x"321e0c",x"2e1b0b",x"351e0d",x"311c0d",x"321d0d",x"2e1b0c",x"29170a",x"361e0d",x"351d0d",x"331c0c",x"341d0c",x"160e07",x"180f07",x"170f07",x"1f1209",x"201309",x"27170a",x"2d1a0c",x"26160a",x"2d1a0b",x"2c190b",x"331d0c",x"2f1b0b",x"301c0b",x"2e1a0b",x"2d190b",x"321c0c",x"301b0b",x"351e0c",x"3f250d",x"41270e",x"472b10",x"3c250b",x"3b250b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"311d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301c0c",x"341d0c",x"381f0d",x"39200e",x"3d220f",x"381f0e",x"391f0d",x"371e0d",x"3a200e",x"3b210f",x"3c230f",x"351e0d",x"311b0c",x"351e0d",x"381f0f",x"341d0d",x"361e0e",x"371f0e",x"371f0e",x"3a200f",x"3a210f",x"381f0e",x"3a200f",x"39200e",x"3d220f",x"3d220f",x"3b210f",x"3a200f",x"3a200e",x"3d2310",x"412511",x"412511",x"3f2410",x"3e2310",x"3b210f",x"422612",x"402511",x"3d2310",x"3a210f",x"3d220f",x"39200e",x"3a200e",x"371f0e",x"2a170a",x"351e0d",x"3c220f",x"3d2310",x"3a220f",x"3f2411",x"3b2411",x"412612",x"422612",x"3f2411",x"3e2310",x"3b210f",x"412511",x"150e07",x"150e07",x"150e07",x"180f07",x"1e1208",x"3f2310",x"2e190b",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2e19",x"4b2e19",x"574031",x"523725",x"5f422d",x"63432b",x"674227",x"67432a",x"654128",x"61412b",x"603d26",x"5b3c29",x"593c2a",x"5c402e",x"5c3f2d",x"5c3f2e",x"593c2b",x"5e402d",x"61422d",x"5f3c27",x"583a28",x"5c3d29",x"613f29",x"5e402b",x"64412a",x"593d2a",x"563a29",x"5e3f2b",x"61402d",x"61412f",x"5a3d2c",x"583f2f",x"543c2d",x"5b3d2b",x"604330",x"5f412d",x"593d2c",x"5b4030",x"5d3e2b",x"563d2d",x"5b3e2b",x"5d4231",x"5d412f",x"5e4332",x"5b4232",x"593d2b",x"5c4333",x"5c412f",x"5d4333",x"563e2d",x"5a402f",x"5b3f2d",x"593e2d",x"5e4231",x"5e4331",x"5d4433",x"634837",x"614330",x"644938",x"6b4e3b",x"694c38",x"6b4d3b",x"674835",x"5e4434",x"604230",x"644735",x"614735",x"5f4533",x"594131",x"664a38",x"644532",x"654733",x"6e4e39",x"684933",x"6c4932",x"644632",x"674a36",x"5a4131",x"5a4232",x"523a28",x"5d412f",x"5b4332",x"5b4230",x"553827",x"523a2b",x"583f2f",x"563b2b",x"593d2d",x"60402d",x"60402b",x"5e3e28",x"5a3d29",x"583d29",x"533b27",x"513624",x"543825",x"593a26",x"5a3b25",x"533724",x"523320",x"472d1d",x"442b1a",x"492f1d",x"472c1b",x"452b1b",x"4d301d",x"452f1f",x"4a3322",x"553218",x"150e07",x"150e07",x"150e07",x"150e07",x"3f230f",x"150e07",x"1c1208",x"21160c",x"22170d",x"23180e",x"24190e",x"281b10",x"22170d",x"23180d",x"25190f",x"2c1f13",x"24190e",x"23180e",x"2a1d11",x"2a1d11",x"25190e",x"291c10",x"26190e",x"271a0f",x"2b1e11",x"2c1e12",x"2e2013",x"281b10",x"2a1d11",x"2a1d11",x"281b0f",x"271a0f",x"2f2014",x"281c10",x"2a1c11",x"281b0f",x"271b0f",x"23170c",x"211508",x"281b10",x"2b1d11",x"2b1e12",x"2c1f12",x"2c1e12",x"291c11",x"2e2013",x"312316",x"2e2013",x"302215",x"342516",x"2c1f13",x"2a1d11",x"2c1e12",x"2c1f12",x"2b1d11",x"281b10",x"291c11",x"2c1e12",x"2a1d11",x"2a1d11",x"2c1e12",x"24180e",x"281b0f",x"2a1d11",x"271b10",x"2a1d11",x"271a0f",x"291c10",x"22170c",x"1f140a",x"1f1308",x"281b10",x"271b10",x"291c11",x"261a0f",x"22170d",x"271b10",x"23180d",x"271b10",x"251a0f",x"251a0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0c",x"311c0c",x"341d0d",x"2d190b",x"2e1a0b",x"2b180b",x"170f07",x"181008",x"1b1108",x"201408",x"2e1b0a",x"301c0c",x"39220e",x"37210e",x"321d0d",x"2e1b0b",x"2e1a0b",x"2e1a0b",x"2f1a0c",x"2a180b",x"2a180b",x"2a180b",x"311c0d",x"331c0d",x"311c0d",x"321d0d",x"321f0e",x"2f1c0d",x"321d0e",x"2d1a0c",x"311c0d",x"311b0c",x"2e1b0c",x"2f1c0d",x"321d0d",x"2d1a0b",x"2b170a",x"2c180a",x"2a170a",x"2a170a",x"2d190b",x"321d0d",x"341e0e",x"311c0c",x"301c0d",x"311d0e",x"311e0e",x"311d0d",x"2e1b0c",x"321c0d",x"321d0d",x"2f1b0c",x"2f1b0c",x"2e1a0b",x"301b0c",x"2f1b0c",x"2e1a0c",x"2d190b",x"301b0c",x"2f1c0d",x"321e0e",x"331f0f",x"301c0d",x"2e1b0c",x"2e1a0c",x"2e1a0b",x"2d190b",x"2e1a0b",x"2f1a0c",x"2d190b",x"2f1b0c",x"2b180b",x"2c190b",x"2f1b0b",x"2e1a0b",x"2c190b",x"2c190b",x"2e1a0c",x"331d0d",x"2d1a0b",x"2c190b",x"29170a",x"29170a",x"2d1a0b",x"2a180b",x"29170a",x"2b180a",x"2b180a",x"26160a",x"29180b",x"311c0d",x"2b180a",x"2d190b",x"2b190b",x"2b180b",x"2a180b",x"28170a",x"26160a",x"2b190b",x"2f1b0c",x"2c190b",x"2b180b",x"2d190b",x"2f1b0c",x"321c0c",x"2e1a0b",x"2e1a0b",x"2d190b",x"2d190b",x"2f1b0c",x"311d0d",x"2a180b",x"2f1a0c",x"2e1a0c",x"321d0d",x"301c0d",x"321d0c",x"311c0c",x"301c0c",x"321c0c",x"2f1b0b",x"321d0b",x"361f0c",x"2c1a0a",x"301d0c",x"34200c",x"2b1b0a",x"251809",x"33200d",x"321e0c",x"301d0d",x"321e0c",x"2c1a0b",x"2a180b",x"2f1b0c",x"2e1b0c",x"2f1b0c",x"2d1a0b",x"2b180a",x"311b0b",x"1a1007",x"1e1308",x"160e07",x"170f07",x"180f07",x"1f1209",x"27170a",x"2e1c0d",x"29190c",x"29180b",x"2b1a0b",x"301c0c",x"2e1b0c",x"311c0d",x"301b0c",x"2e1a0b",x"331c0d",x"311c0c",x"3b230e",x"452a10",x"492c0f",x"42290e",x"3d250c",x"3f270c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"392110",x"150e07",x"231409",x"2f1b0c",x"331d0d",x"2f1b0c",x"2e1a0b",x"331c0c",x"371e0d",x"3a200e",x"3b210f",x"391f0d",x"3a200e",x"361d0d",x"391f0d",x"371e0d",x"341c0c",x"341d0d",x"381f0e",x"3c220f",x"371f0e",x"311c0d",x"321c0c",x"371f0e",x"381f0d",x"341c0c",x"361e0d",x"371f0e",x"3c210f",x"3b220f",x"3c220f",x"402411",x"3c210f",x"361d0d",x"341c0c",x"371e0d",x"351d0d",x"341c0c",x"371e0d",x"3b210f",x"3b210f",x"3d220f",x"3c220f",x"3d2310",x"3f2410",x"3a1f0e",x"341c0c",x"371e0d",x"361e0d",x"381f0e",x"3d2310",x"3d2210",x"3a210f",x"3b210f",x"3e2310",x"412511",x"3b210f",x"3e2310",x"402511",x"3c210f",x"381e0d",x"3c210e",x"150e07",x"2f1a0c",x"371f0e",x"351f0e",x"311c0d",x"381f0c",x"341d0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462915",x"462915",x"4e3b2e",x"563f30",x"543927",x"5e402d",x"5d3b26",x"603f2a",x"67432c",x"65432d",x"63432f",x"63432e",x"604330",x"674631",x"5d402c",x"553a28",x"634532",x"583c28",x"573a28",x"5c3c29",x"5f3e2a",x"63402b",x"634028",x"603f29",x"5c3c28",x"5b3b27",x"573b29",x"5d3d2a",x"5d412f",x"5f4231",x"5b3d2d",x"593e2d",x"533b2d",x"563f30",x"584031",x"5c412f",x"5b4232",x"614331",x"5f412f",x"593e2d",x"5a4130",x"553c2c",x"5b4231",x"573c2c",x"5a3e2e",x"5a3e2d",x"5f402d",x"5b3e2c",x"553b2a",x"5b3f2e",x"583e2d",x"573c2a",x"51382a",x"594031",x"583e2e",x"584132",x"574032",x"5a4131",x"5d4333",x"5f412e",x"5f4230",x"634431",x"5f412f",x"593d2c",x"543b2b",x"5c4030",x"5f4434",x"5c4232",x"604535",x"684a37",x"624735",x"634634",x"644635",x"644734",x"614431",x"60432f",x"5f412f",x"5c4333",x"584030",x"544032",x"594335",x"554235",x"5d4434",x"614633",x"5e4331",x"624736",x"5e4332",x"593c2a",x"5a3c2a",x"5b3e2c",x"593a27",x"5b3d2a",x"5b3d29",x"573824",x"5a3c26",x"5d3f2b",x"553622",x"583823",x"583925",x"4f321f",x"4b301d",x"4b301d",x"4c301e",x"4a2f1d",x"4e301d",x"452d1d",x"4c2f1f",x"523727",x"553118",x"150e07",x"150e07",x"150e07",x"150e07",x"492a14",x"150e07",x"20150c",x"20150b",x"21160c",x"22170d",x"24180d",x"25190e",x"21160c",x"23180d",x"281b10",x"24190e",x"24190e",x"271b10",x"271b10",x"2a1d11",x"2d2013",x"271a0f",x"2d2013",x"2d2013",x"2c1f13",x"2b1e12",x"2d1f13",x"2d1f13",x"2e2013",x"2f2114",x"2c1e12",x"2a1d11",x"2c1e12",x"2a1d11",x"2c1e12",x"2d1f13",x"2c1e11",x"2f2013",x"281b0f",x"271b0f",x"271a0f",x"2a1c11",x"281b0f",x"271b0f",x"2b1d11",x"2b1e12",x"2f2114",x"291c11",x"2b1e12",x"2d1f13",x"2d1f13",x"2c1f12",x"2f2114",x"2b1d11",x"322316",x"2f2114",x"2c1f13",x"2b1e12",x"2d1f13",x"2b1d12",x"2b1d11",x"2b1e11",x"302114",x"2c1e12",x"2a1d11",x"312215",x"281b10",x"2d1f13",x"2d1f12",x"22170c",x"22170d",x"26190f",x"24180d",x"22170d",x"21160c",x"26190e",x"23180d",x"261a0f",x"21160c",x"261a0f",x"261a0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1a0b",x"2d1a0b",x"2f1b0c",x"301b0c",x"2a170a",x"160e07",x"170f07",x"170f07",x"1c1107",x"28180a",x"26170a",x"2d1b0b",x"331e0c",x"2e1a0b",x"321d0c",x"301c0b",x"2a170a",x"28160a",x"2a170a",x"2a180b",x"2b180b",x"2d1a0c",x"2d1a0c",x"2d1a0b",x"2a180b",x"311c0c",x"321c0d",x"2f1b0c",x"2d1a0c",x"301b0c",x"2b180b",x"2a170a",x"2d190b",x"2d190b",x"2f1a0c",x"311c0c",x"321d0d",x"301c0d",x"311c0d",x"2f1a0c",x"2e1a0b",x"2f1a0b",x"301b0c",x"331d0d",x"301b0c",x"301c0d",x"311c0d",x"341f0e",x"321d0d",x"311c0c",x"341d0d",x"2d190b",x"27160a",x"2f1a0c",x"2f1b0c",x"2f1a0c",x"2f1b0c",x"2b180b",x"2c190b",x"2a180b",x"2b180b",x"2a180b",x"29180a",x"2e1a0c",x"2c1a0c",x"321d0d",x"2e1b0c",x"311c0d",x"321c0d",x"2c190b",x"2d190b",x"331d0d",x"28180b",x"321c0d",x"29170a",x"2b180b",x"301b0c",x"301b0c",x"2d1a0b",x"2e1a0b",x"29170a",x"271609",x"28160a",x"231409",x"29170a",x"211309",x"28170a",x"261509",x"261509",x"261509",x"261609",x"29170a",x"2d190b",x"2d1a0b",x"28170a",x"2d190b",x"2a170a",x"2a180b",x"29170a",x"29170a",x"29170a",x"2c190b",x"2d1a0b",x"301b0c",x"27170a",x"2d190b",x"2b180b",x"29160a",x"29170a",x"2b180b",x"29170a",x"2d190b",x"2d190b",x"2d1a0b",x"2e1a0c",x"2d190b",x"321d0c",x"341f0c",x"37200d",x"301b0b",x"2d1a0a",x"2f1b0b",x"351f0c",x"37210d",x"2f1c0a",x"2b1b0a",x"2e1c0a",x"2f1c0b",x"341e0d",x"2e1c0a",x"2f1c0c",x"28180a",x"26160a",x"28160a",x"27160a",x"2b180b",x"29170a",x"2f1b0c",x"301c0c",x"341e0d",x"1f1408",x"1d1308",x"1a1107",x"170f07",x"180f07",x"180f07",x"1b1008",x"25150a",x"2c190b",x"2d1a0c",x"2b1a0b",x"2b180b",x"2b180b",x"2d190b",x"301a0c",x"29170a",x"2d1a0b",x"331e0d",x"3d240e",x"43280f",x"462b10",x"3e260d",x"3c250c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"2e1b0c",x"150e07",x"1e1208",x"2e1a0b",x"2e190b",x"2e190b",x"371e0d",x"311b0c",x"2d1a0b",x"2e1a0b",x"2a160a",x"2b170a",x"2c190b",x"2c190b",x"2d1a0b",x"2f1b0c",x"2d190b",x"2d1a0b",x"2e1a0c",x"2e1a0c",x"2d1a0c",x"27170a",x"29180b",x"2b180b",x"2d1a0b",x"2c190b",x"2c190b",x"2d1a0c",x"2d1a0b",x"2f1c0c",x"321d0d",x"351e0e",x"321d0e",x"341e0e",x"2d1a0b",x"311c0c",x"331d0d",x"311c0d",x"321c0d",x"2d190b",x"311b0c",x"321c0d",x"341e0e",x"2d190b",x"331d0d",x"341e0e",x"2f1b0c",x"321d0d",x"321d0d",x"301b0c",x"2f1b0c",x"301b0c",x"341e0e",x"331d0d",x"311c0d",x"2f1b0c",x"321c0d",x"361f0e",x"361f0e",x"331d0d",x"3d220f",x"180f08",x"27170a",x"341d0d",x"371f0e",x"361f0e",x"2b180b",x"3e220e",x"2e190a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492b16",x"492b16",x"4a382b",x"4f382a",x"5f412e",x"64422c",x"624028",x"6a472f",x"6b442c",x"654733",x"593d2a",x"5c402e",x"5b402f",x"523c2c",x"543928",x"583e2e",x"573c2c",x"5c3c29",x"563621",x"5d3d2a",x"5d3d27",x"5d3f2b",x"553825",x"543725",x"583a26",x"593a28",x"583926",x"5b3e2c",x"543827",x"553b2c",x"5a3c29",x"563a29",x"593d2c",x"5c3f2d",x"5c3f2e",x"5e3e2c",x"63432e",x"61432f",x"5d402f",x"624532",x"604331",x"5e412f",x"5f4330",x"60422f",x"5c4130",x"62442f",x"604331",x"5d4230",x"624632",x"644532",x"614432",x"644632",x"5a4333",x"5a4232",x"644835",x"644735",x"624736",x"584233",x"583f2f",x"5e4333",x"5f4331",x"644735",x"614534",x"654835",x"644632",x"654734",x"6a4a36",x"604433",x"624533",x"644735",x"644735",x"614735",x"664935",x"664835",x"62412d",x"654732",x"654733",x"634634",x"624939",x"5e4434",x"594335",x"574133",x"594233",x"5a4233",x"5d412f",x"5e4534",x"5c4231",x"5a3f2e",x"5a3f2e",x"553a29",x"543a29",x"593c2b",x"593b29",x"5c3d2b",x"593d2a",x"593a28",x"573a27",x"5a3b28",x"5e3c28",x"503624",x"503422",x"4c3220",x"472e1f",x"4a2d1a",x"4d301f",x"4f2f1c",x"553622",x"4d3526",x"512e15",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2c15",x"150e07",x"23180e",x"261a0f",x"251a0f",x"2a1d11",x"261a0f",x"24190e",x"2b1e12",x"25190f",x"291c11",x"24190f",x"251a0f",x"2b1e12",x"261a0f",x"291c11",x"2a1d11",x"261a0f",x"201409",x"2a1c11",x"2f2114",x"2b1e11",x"281c10",x"2c1f13",x"2e2013",x"2f2014",x"302215",x"2b1e12",x"302215",x"2c1f13",x"2e2014",x"2e2012",x"291c10",x"2a1d12",x"2b1e12",x"342516",x"2f2014",x"2e2014",x"2f2114",x"332416",x"2f2114",x"312215",x"322316",x"312215",x"322316",x"362719",x"322316",x"2b1e11",x"2a1d11",x"291d11",x"211509",x"2a1d11",x"291c11",x"2d1f12",x"2b1d11",x"302215",x"2c1f12",x"2d1f13",x"302215",x"2d1f13",x"2e2014",x"302215",x"2b1e12",x"2a1d11",x"281b0f",x"25190f",x"2b1e12",x"2d2013",x"291c11",x"2e2014",x"2b1e12",x"261a10",x"261a0f",x"281c10",x"2b1e12",x"271b10",x"271b10",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0c",x"311c0c",x"311d0c",x"321d0e",x"341e0e",x"160e07",x"170f07",x"180f08",x"1d1208",x"2c1b0a",x"2b190b",x"29180a",x"311c0c",x"351f0d",x"321d0c",x"2e1a0c",x"321d0d",x"331e0e",x"331d0e",x"2f1b0c",x"2f1b0c",x"2e1a0b",x"301b0c",x"341d0e",x"301c0d",x"311c0d",x"331d0d",x"2b190b",x"331d0d",x"321c0d",x"311c0c",x"321c0d",x"321c0c",x"311c0c",x"311c0d",x"301b0c",x"321c0d",x"311c0c",x"311c0c",x"2e1a0b",x"301b0c",x"2c180b",x"2c180b",x"2d190b",x"2d190b",x"2f1a0c",x"2f1b0c",x"311c0d",x"2f1a0c",x"2e1a0b",x"2d190b",x"2e1a0c",x"2f1a0c",x"331d0d",x"2c190b",x"271509",x"26160a",x"27160a",x"2d190b",x"301c0d",x"2d1a0c",x"2c190b",x"301c0d",x"311c0d",x"2e1b0c",x"2c190b",x"2b190b",x"2b190b",x"2a180b",x"27160a",x"2a180b",x"2e1a0b",x"2f1a0c",x"29170a",x"29180b",x"25150a",x"2a170a",x"2a180b",x"2a170a",x"2a180b",x"2c190b",x"2b180b",x"28160a",x"211309",x"241409",x"201309",x"241509",x"27160a",x"321c0c",x"2c190b",x"2a180b",x"2d190b",x"2f1c0d",x"301b0c",x"301b0c",x"311c0d",x"311c0d",x"321c0d",x"321c0d",x"2a180b",x"301c0d",x"2f1b0c",x"2c190b",x"2c1a0c",x"2e1b0c",x"2c1a0c",x"311c0d",x"311c0d",x"2f1a0c",x"321d0d",x"2b190b",x"2f1b0c",x"2d1a0c",x"28170a",x"2c190b",x"301c0d",x"2e1c0b",x"2c1a0b",x"2f1c0c",x"341f0d",x"38220e",x"301c0c",x"301d0c",x"331e0c",x"2e1b0a",x"311d0b",x"2f1c0b",x"2f1c0b",x"281909",x"2b1a0b",x"2b190b",x"27170a",x"2b190b",x"2f1b0b",x"26160a",x"29180b",x"2a180b",x"2c190b",x"2c190b",x"331d0c",x"201408",x"1e1308",x"180f07",x"180f07",x"170f07",x"1e1208",x"1c1108",x"1d1208",x"241509",x"28170a",x"29180b",x"29170b",x"2e1a0b",x"2b180b",x"2a180b",x"2c1a0b",x"2d1a0b",x"2e1a0b",x"341e0c",x"40270d",x"43290f",x"37220c",x"38220b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"191008",x"351e0e",x"150e07",x"201309",x"331d0d",x"392110",x"382010",x"1d1108",x"3e220f",x"402410",x"452712",x"472813",x"472913",x"462913",x"462812",x"452712",x"412310",x"412310",x"432611",x"442611",x"442612",x"472813",x"402511",x"442712",x"412411",x"402410",x"412410",x"422511",x"3f2310",x"422511",x"412410",x"422510",x"452712",x"442612",x"452812",x"452712",x"462812",x"412410",x"402310",x"422511",x"432611",x"412410",x"402410",x"432611",x"432611",x"432612",x"452712",x"402310",x"442711",x"452712",x"432611",x"452711",x"432611",x"492913",x"442612",x"482913",x"442712",x"472812",x"452711",x"452712",x"432611",x"462711",x"150e07",x"2b180b",x"371f0e",x"38200e",x"351e0d",x"2f1b0c",x"371e0c",x"341d0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2c17",x"4a2c17",x"543d2d",x"503421",x"553927",x"61412d",x"5e3b22",x"67412a",x"613f28",x"66442f",x"5d3e2a",x"634532",x"5e422f",x"5e4535",x"5e3f2b",x"5a4233",x"583b29",x"5c3c26",x"5b3b28",x"5e3c26",x"613d27",x"664029",x"69442d",x"67432d",x"613d27",x"573b29",x"573927",x"5a3e2d",x"60412d",x"60412d",x"614431",x"5c3f2d",x"614330",x"5a3d2c",x"5b3f2d",x"5e412f",x"614331",x"60412e",x"5f422e",x"604331",x"5d4230",x"5d402d",x"5b3f2e",x"573b2a",x"5a3d2a",x"573c2b",x"5d3f2c",x"583b29",x"5b3c28",x"553827",x"553927",x"543926",x"5b402f",x"563e2e",x"5a402f",x"543c2c",x"594131",x"584031",x"563f2f",x"5b4131",x"5e4330",x"604533",x"634633",x"644734",x"5d4232",x"604534",x"684935",x"634533",x"614532",x"5f4130",x"664835",x"5c4231",x"634632",x"654835",x"614633",x"664735",x"644734",x"624634",x"5c4232",x"5a4030",x"594334",x"573f2f",x"543d2f",x"574133",x"574132",x"5e4535",x"5e4435",x"523929",x"563b29",x"5e402e",x"5e412d",x"60422e",x"60422e",x"60412d",x"5a3d29",x"5b3e2b",x"5e3f2a",x"5b3d2a",x"5d3d27",x"5a3b29",x"593924",x"573823",x"533725",x"4f2f1b",x"573824",x"553722",x"533726",x"533c2c",x"59351a",x"150e07",x"150e07",x"150e07",x"150e07",x"4b2b15",x"150e07",x"271b0f",x"271b10",x"21160c",x"23180e",x"261a0f",x"23180e",x"22170d",x"2b1e12",x"291c10",x"25190e",x"24190e",x"281c10",x"2b1d11",x"281c10",x"2a1d11",x"2c1e12",x"2a1d11",x"2d1f13",x"2b1e12",x"2a1d11",x"2d1f13",x"2d2013",x"2d1f12",x"2b1e12",x"2e2114",x"312316",x"2e2014",x"332417",x"2f2114",x"281b0f",x"322316",x"2e2013",x"2a1d11",x"302114",x"2e2013",x"2a1d11",x"2c1e12",x"2e2013",x"302114",x"2f2114",x"322214",x"312214",x"342517",x"2c1e12",x"2e2013",x"322316",x"2d1f13",x"2c1f12",x"302114",x"2d1f13",x"302114",x"2c1e12",x"302114",x"2d2013",x"302114",x"2d1f13",x"312315",x"312316",x"2e2014",x"2e2014",x"302114",x"291d10",x"2b1e12",x"2c1e12",x"291c10",x"291d11",x"261a0f",x"271a0f",x"261a0f",x"281c10",x"281b10",x"2d2013",x"21170c",x"261a0e",x"261a0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341d0d",x"341d0d",x"331d0d",x"351d0d",x"341e0d",x"160e07",x"1d1208",x"1d1208",x"2a1a09",x"2e1c0b",x"321d0c",x"2e1b0b",x"311c0c",x"2f1b0b",x"2f1b0c",x"311c0d",x"2e1a0c",x"2f1a0b",x"311c0c",x"321d0d",x"301b0c",x"2f1b0c",x"2f1b0c",x"311c0d",x"321c0d",x"331d0d",x"311d0d",x"2e1a0c",x"311c0c",x"321c0c",x"2d1a0b",x"2e190b",x"301a0b",x"331c0d",x"311b0c",x"311c0d",x"301b0c",x"2f1b0c",x"301b0c",x"2d190b",x"2f1a0b",x"2e1a0b",x"2d1a0b",x"2f1b0c",x"341e0d",x"321d0d",x"321d0d",x"2f1b0d",x"321d0d",x"2f1b0c",x"2d190b",x"2d1a0b",x"2d1a0b",x"2a180b",x"2d1a0b",x"2e1a0c",x"2b180b",x"2a180b",x"2c1a0b",x"27160a",x"26160a",x"27170a",x"28170b",x"2b190b",x"29180b",x"2b180b",x"2a180b",x"2d1a0c",x"2e1a0c",x"2b180b",x"2a180b",x"2c190b",x"2b180b",x"29170a",x"2d190b",x"27160a",x"2f1b0c",x"2f1b0d",x"2f1c0d",x"2f1b0d",x"2c190b",x"2a180b",x"25150a",x"28170a",x"25160a",x"24150a",x"29180b",x"29170b",x"2a180b",x"29170a",x"2a180b",x"29170b",x"2c190b",x"2d1a0b",x"2b180b",x"301c0c",x"2f1b0c",x"2e1a0b",x"2c180b",x"2c190b",x"2d190b",x"2b180b",x"27160a",x"27160a",x"2c190b",x"311c0c",x"2c190b",x"2e1a0c",x"311c0d",x"2f1a0c",x"2c190b",x"2a180b",x"2d190b",x"2b180b",x"2e1a0b",x"2c190b",x"2c190b",x"2f1c0b",x"2d1a0b",x"2d1a0b",x"2e1a0b",x"35200d",x"341f0c",x"311e0b",x"331f0c",x"2c1b0a",x"24160a",x"261709",x"221509",x"2e1b0c",x"2c1a0b",x"311d0b",x"2b190b",x"2c190b",x"241509",x"231409",x"2d1a0b",x"2d1a0b",x"2e1a0c",x"1b1107",x"1c1108",x"1b1108",x"1b1107",x"190f08",x"1b1108",x"211409",x"221409",x"26160a",x"26160a",x"27170a",x"28170b",x"2e1b0c",x"2a180b",x"29180b",x"28170a",x"28170a",x"2e1b0c",x"301c0c",x"3a220d",x"3d240e",x"452910",x"36210b",x"36210b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"311c0c",x"150e07",x"150e07",x"321d0d",x"341d0d",x"321c0d",x"311d0d",x"3c2311",x"402511",x"3f2410",x"3e2310",x"3f2411",x"402512",x"412612",x"402512",x"412612",x"412612",x"402612",x"402612",x"39200e",x"38200f",x"402612",x"3e2512",x"3d2411",x"3b2310",x"3a2110",x"3a2110",x"38200f",x"3b2311",x"3b2311",x"3e2411",x"402512",x"3c2311",x"3c2310",x"3c220f",x"3c220f",x"3c2310",x"38200e",x"38200e",x"38200e",x"382210",x"3b2310",x"3c2310",x"3b2210",x"3a220f",x"38200e",x"3c230f",x"3a210f",x"3a2110",x"3d2411",x"3a2110",x"351e0e",x"3d2310",x"38200e",x"3a200e",x"391f0d",x"311a0b",x"30190a",x"321a0b",x"361e0d",x"3d2310",x"4a2b15",x"25160a",x"38200f",x"38200f",x"38200f",x"341e0e",x"40230f",x"2e190a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2e18",x"4d2e18",x"503e32",x"563e2e",x"533a29",x"5f3f2c",x"64432c",x"66452f",x"62412c",x"623f28",x"61412c",x"674833",x"594232",x"5b402e",x"614737",x"5c3d29",x"553724",x"553927",x"553622",x"5b3b27",x"5c3e2c",x"5c3c27",x"64422c",x"60412c",x"64432d",x"63422d",x"5f3f2a",x"62432f",x"5c3d29",x"61432f",x"583d2c",x"603f2a",x"664630",x"654632",x"6a4a34",x"6b482f",x"6b4a35",x"664530",x"5c3f2d",x"5c422f",x"674a35",x"614430",x"5d412f",x"5e4230",x"644734",x"644734",x"644633",x"654531",x"664935",x"644733",x"58402f",x"614736",x"5f4736",x"5e4432",x"564030",x"5f4533",x"594334",x"594233",x"5e4432",x"634633",x"604433",x"5d422f",x"634531",x"634431",x"604432",x"654734",x"674a38",x"694b36",x"6b4b37",x"634330",x"60422f",x"5f4533",x"614331",x"614432",x"533b2c",x"583c2d",x"553c2e",x"573b2b",x"624533",x"684935",x"614634",x"5d4330",x"5c4333",x"604735",x"5b4232",x"624736",x"5c4331",x"5c4332",x"614632",x"5e4332",x"654733",x"624430",x"604331",x"63432d",x"5e3f2c",x"5e3f2c",x"5f3e29",x"5b3c2a",x"5a3d2b",x"5e402e",x"553827",x"5c3a24",x"4b3121",x"50311b",x"533624",x"5d3a24",x"513826",x"563b29",x"512e16",x"150e07",x"150e07",x"150e07",x"150e07",x"4a2b15",x"150e07",x"2a1e12",x"261a0f",x"261a0f",x"281c10",x"251a0f",x"261a10",x"21170d",x"23180d",x"23180d",x"271b0f",x"2d2013",x"291c10",x"291d11",x"2c1f12",x"2d1f13",x"2b1d11",x"2a1d12",x"2b1e12",x"2c1f13",x"2d1f12",x"322316",x"2e2013",x"302215",x"2b2014",x"35281a",x"2f2215",x"372719",x"322316",x"322316",x"322417",x"2e2014",x"2c2014",x"2f2114",x"302114",x"2f2114",x"2e2013",x"2f2114",x"302215",x"2e2014",x"312215",x"291c10",x"2f2013",x"352618",x"332416",x"2f2114",x"342516",x"352517",x"332416",x"352618",x"322316",x"302215",x"2c1f12",x"2e2013",x"312215",x"39291a",x"342719",x"302417",x"312416",x"322416",x"302215",x"2f2114",x"352618",x"2e2014",x"2c2014",x"2e2114",x"302114",x"2f2114",x"2a1d11",x"2d1f13",x"302215",x"2a1d11",x"2e2013",x"26190e",x"291c0f",x"291c0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38210f",x"38210f",x"39200f",x"351e0e",x"38200f",x"160e07",x"201408",x"221509",x"271909",x"2c1b0a",x"301c0c",x"301c0c",x"311d0d",x"321d0d",x"321c0d",x"341e0e",x"311c0d",x"341e0d",x"321c0d",x"37200f",x"36200f",x"351f0e",x"331d0d",x"321d0d",x"311c0c",x"301b0c",x"2d190b",x"2a170a",x"291609",x"281609",x"2c180b",x"321c0d",x"331d0d",x"351f0e",x"311c0d",x"311d0d",x"351f0f",x"331d0e",x"341f0e",x"341f0e",x"331e0e",x"36200f",x"331e0e",x"311c0d",x"321d0e",x"311d0d",x"301c0d",x"301c0c",x"2e1a0b",x"2f1a0c",x"2d190b",x"311c0d",x"2e1a0b",x"2d190b",x"2d1a0b",x"2c190b",x"2d190b",x"2f1b0c",x"2f1b0c",x"2c190c",x"29180b",x"2b190c",x"2e1b0d",x"2d1a0c",x"2a180b",x"26160a",x"2a190b",x"2e1a0c",x"2b190b",x"2c190b",x"2c1a0c",x"29180b",x"2f1b0c",x"29170a",x"27160a",x"27160a",x"2d190b",x"2c190b",x"2b190b",x"2e1a0c",x"2d1a0c",x"2f1c0d",x"2d1a0c",x"2a180b",x"29180b",x"2d1a0c",x"2a180b",x"2c1a0c",x"2e1b0d",x"331e0e",x"321e0e",x"341f0f",x"2e1b0d",x"2b180b",x"311d0d",x"321e0e",x"331f0e",x"321d0e",x"2f1b0d",x"2d1a0c",x"301c0d",x"301c0d",x"2d1a0c",x"301c0d",x"311c0d",x"311c0d",x"311c0d",x"301b0c",x"2b190b",x"311c0d",x"2e1a0c",x"2c190b",x"29170a",x"2d1a0c",x"301d0d",x"311c0c",x"2f1c0c",x"311c0d",x"321d0c",x"2e1b0b",x"321d0d",x"351f0d",x"311d0d",x"331f0c",x"321e0c",x"301d0b",x"25160a",x"211408",x"211409",x"2b190a",x"271609",x"281709",x"271609",x"2d190b",x"2a190b",x"2c1a0c",x"36200f",x"2d1b0c",x"39210f",x"201409",x"1f1309",x"251709",x"201409",x"1d1209",x"1b1108",x"211409",x"24150a",x"24150a",x"27170b",x"2f1b0c",x"25160a",x"231409",x"28170a",x"27160a",x"2b190b",x"2e1a0b",x"2d1a0b",x"2c1a0b",x"321d0c",x"38220d",x"3f270e",x"3b250c",x"3b250c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1b1008",x"311c0d",x"150e07",x"180f08",x"24150a",x"301b0c",x"28170a",x"2f1a0b",x"381f0d",x"3a200e",x"391f0e",x"3d220f",x"412511",x"412611",x"402511",x"3e2310",x"462913",x"452813",x"452914",x"452914",x"432813",x"422612",x"3f2612",x"442913",x"422712",x"3c2411",x"472a14",x"432813",x"3f2512",x"422713",x"402612",x"452913",x"472b15",x"452914",x"432713",x"3f2411",x"3f2411",x"3c210f",x"3b210f",x"3d220f",x"391f0d",x"381f0d",x"3b210f",x"391f0e",x"3c220f",x"3b210f",x"3c220f",x"381f0d",x"3a210f",x"3b210f",x"3d2310",x"3d2310",x"3b210f",x"3d220f",x"3d2310",x"442813",x"3f2310",x"432612",x"432712",x"412612",x"432611",x"422511",x"482913",x"150e07",x"321d0d",x"301c0d",x"321d0d",x"2a180b",x"3f220e",x"361e0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492c18",x"492c18",x"564234",x"5f4736",x"5c3f2d",x"624430",x"62422e",x"684831",x"68442b",x"664731",x"64432d",x"624531",x"664b36",x"674833",x"61432e",x"5a3c28",x"583a28",x"583926",x"5c3b25",x"5e3d28",x"613e27",x"5f3d25",x"5f3d27",x"5d3d29",x"583825",x"593a27",x"583a27",x"5b3e2c",x"553c2c",x"553d2c",x"5d412d",x"634330",x"644533",x"644734",x"604533",x"624532",x"664734",x"654834",x"61432f",x"5a4231",x"624530",x"60422e",x"624735",x"573d2c",x"644632",x"614431",x"604432",x"654734",x"624532",x"694a36",x"674b37",x"614734",x"5e422f",x"624634",x"59402f",x"5a4131",x"594133",x"543c2e",x"553f31",x"5b412f",x"5e4231",x"5f4535",x"604332",x"5d412f",x"5a3f2f",x"5b3f2e",x"5c402e",x"654632",x"63442f",x"5c412f",x"604330",x"583d2a",x"664632",x"5f412d",x"63432e",x"62432e",x"674a35",x"634430",x"614432",x"5b3f2d",x"593e2c",x"5d3f2c",x"593e2d",x"553b2a",x"593f2e",x"594132",x"5b4231",x"594030",x"584030",x"5b4232",x"5e4231",x"634734",x"60432f",x"62432e",x"64432f",x"63432e",x"634532",x"624430",x"61422c",x"5f402c",x"64412b",x"5c3c27",x"5f3f2a",x"573924",x"60402c",x"623f27",x"5a3d29",x"523c2d",x"513017",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2c15",x"150e07",x"271b10",x"24190e",x"24190f",x"2d2013",x"271b10",x"261a0f",x"24190e",x"23180e",x"2b1e12",x"261a0f",x"281b10",x"2a1d11",x"25190e",x"2d1f13",x"291c11",x"2d1f13",x"2d1f13",x"2c1f13",x"312214",x"2b1e12",x"2d2013",x"302214",x"2f2114",x"2f2114",x"332416",x"352517",x"2f2114",x"312215",x"302215",x"302416",x"2c1f13",x"302215",x"2e2114",x"302214",x"302215",x"342517",x"302316",x"322316",x"302215",x"2f2114",x"2d2013",x"302214",x"2d1f13",x"312215",x"322315",x"2f2014",x"2d1f13",x"332416",x"332416",x"352617",x"312214",x"322316",x"322316",x"332416",x"322316",x"362617",x"2f2014",x"372719",x"2d2013",x"2d1f13",x"2a1d11",x"2e2215",x"2e2114",x"322416",x"2c1f13",x"2e2013",x"2c1f13",x"2f2115",x"2c2013",x"2d2013",x"2c1f13",x"291d11",x"291d11",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452813",x"452813",x"3c2411",x"37200f",x"341f0f",x"1a1107",x"1c1207",x"1c1107",x"261709",x"2d1b0b",x"301c0b",x"2a180a",x"2c190b",x"2a180b",x"311b0c",x"2f1b0c",x"2e1a0c",x"2b180b",x"2f1b0c",x"311c0c",x"321c0d",x"2e1b0c",x"301b0c",x"2f1a0c",x"2e1a0c",x"321d0d",x"331d0d",x"301c0d",x"331d0d",x"301c0d",x"321c0d",x"321c0d",x"28170b",x"2f1b0c",x"311c0d",x"2e1a0c",x"301c0d",x"2d1a0c",x"311c0d",x"2d1a0c",x"2f1b0d",x"301c0d",x"2c190b",x"28170b",x"311d0d",x"341e0e",x"311d0d",x"2d1a0b",x"2e1b0c",x"2d1a0c",x"2e1b0c",x"2f1c0d",x"2e1a0c",x"2d1a0c",x"2f1b0c",x"2f1c0d",x"301c0d",x"2f1c0d",x"2f1c0d",x"2b190c",x"2b190c",x"2a180b",x"2d1b0d",x"2c1a0c",x"2d1b0c",x"2d1b0c",x"2c190c",x"2c1a0c",x"2d1b0d",x"2d1b0d",x"2b190c",x"2a180b",x"2a180b",x"2b190b",x"28170b",x"2c1a0c",x"2c190b",x"2a180b",x"29170a",x"28160a",x"28170a",x"261509",x"27160a",x"29170a",x"26160a",x"2b190b",x"2f1b0d",x"2b190b",x"2a190b",x"28170b",x"2d1a0c",x"301c0d",x"2d1b0d",x"2d1b0c",x"2d1b0c",x"2e1b0d",x"2f1c0d",x"301d0d",x"2f1c0d",x"2e1b0d",x"2c1a0c",x"2d1b0c",x"2d1b0c",x"2b190c",x"2d1b0d",x"2f1c0d",x"301c0d",x"2f1c0d",x"2f1c0c",x"2c190c",x"29170a",x"2d190b",x"26160a",x"29170a",x"26150a",x"29170b",x"28160a",x"2f1a0b",x"2f1c0c",x"2a190b",x"29170a",x"29180b",x"2b180b",x"341f0d",x"321d0b",x"2d1b0b",x"1d1108",x"26170a",x"241709",x"2c190b",x"2d1a0c",x"2b190b",x"28170b",x"2b190b",x"29180b",x"29180b",x"2c190b",x"2f1b0c",x"321c0d",x"1f1309",x"221509",x"221509",x"1c1108",x"1d1208",x"1c1108",x"211309",x"24160a",x"27170b",x"1f1309",x"28170b",x"26160a",x"25160a",x"2a180b",x"27170a",x"27160a",x"29180b",x"331f0c",x"331d0d",x"37210d",x"42280f",x"4a2d13",x"38230b",x"38230b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231409",x"331d0d",x"150e07",x"321b0b",x"2e190b",x"301a0b",x"311b0c",x"2d190b",x"341c0c",x"391f0e",x"381f0e",x"3a210f",x"3f2310",x"3e2310",x"3f2410",x"3c220f",x"402410",x"412511",x"412611",x"3f2511",x"3f2411",x"412512",x"351d0d",x"361e0d",x"3d2411",x"361f0e",x"3e2310",x"422612",x"3f2511",x"3f2411",x"3f2411",x"3e2411",x"432713",x"412612",x"402512",x"3f2511",x"3f2512",x"3b2210",x"361e0e",x"351d0d",x"381f0e",x"341d0d",x"39210f",x"3e2410",x"3b220f",x"3f2410",x"402511",x"3b2310",x"3f2411",x"412612",x"3e2411",x"3e2410",x"3f2310",x"402511",x"3c220f",x"3c220f",x"3d2310",x"422612",x"432712",x"3d220f",x"402511",x"412611",x"4b2a14",x"341e0e",x"3b210f",x"402410",x"1d1108",x"150e07",x"391f0c",x"381f0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492c17",x"492c17",x"5d493a",x"5a402d",x"5b402d",x"5c3f2b",x"61412d",x"644531",x"65442f",x"64432c",x"62432e",x"6a4e3c",x"654835",x"694d39",x"604330",x"573a28",x"573826",x"563927",x"573723",x"4d3120",x"503524",x"533727",x"563724",x"543827",x"583b28",x"5d3f2c",x"563d2c",x"583f2e",x"664836",x"5f4331",x"614534",x"5e4534",x"614431",x"5b402f",x"624735",x"5c4434",x"594132",x"5c4434",x"614430",x"594132",x"5d4536",x"5b4333",x"5d4433",x"5e4534",x"593e2d",x"614634",x"5b4333",x"5a3f2e",x"5e4433",x"624734",x"593f2e",x"624736",x"614532",x"614432",x"614532",x"624632",x"584132",x"553f30",x"583f30",x"5b4334",x"644836",x"5e4433",x"5f4433",x"654836",x"654935",x"5d422f",x"694a36",x"644632",x"5f422f",x"5c402d",x"5d4231",x"5b402d",x"5d402d",x"5f412d",x"634531",x"63442f",x"64442f",x"5c3d2a",x"5b3d2a",x"5c3e2b",x"60402c",x"583c29",x"5b402f",x"563d2d",x"594233",x"543f31",x"5b4130",x"60422f",x"583f2f",x"664632",x"5a412f",x"5c412f",x"5d412f",x"60412e",x"604431",x"61432f",x"62432f",x"614531",x"5b402e",x"563b29",x"62412b",x"62412b",x"5f402b",x"5d3e29",x"5c3d28",x"624129",x"5d412e",x"523c2d",x"56331a",x"150e07",x"150e07",x"150e07",x"150e07",x"482a14",x"150e07",x"2a1d11",x"261a10",x"21170d",x"291c10",x"261a0f",x"291c11",x"2a1d11",x"271b10",x"261a0f",x"251a0f",x"2c1f13",x"2b1e12",x"291c10",x"281b10",x"2d2013",x"2b1e12",x"2e2014",x"2c1f13",x"312316",x"312215",x"2f2114",x"312316",x"312316",x"302215",x"312215",x"322316",x"2f2114",x"312316",x"2c1f13",x"322316",x"332416",x"2f2114",x"332416",x"2e2014",x"352618",x"2f2013",x"322315",x"322315",x"332416",x"332417",x"352517",x"2e2013",x"2c1f13",x"352517",x"312215",x"302114",x"342416",x"342416",x"332416",x"362718",x"362719",x"342516",x"342416",x"342517",x"3a291b",x"302215",x"2d1f13",x"2f2114",x"2f2114",x"2b1e12",x"2c1f13",x"2e2013",x"2e2014",x"372719",x"2e2014",x"302214",x"2a1d12",x"23180d",x"2b1d11",x"2f2114",x"2a1d11",x"2c1f13",x"2c1f12",x"2b1d12",x"2b1d12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a210f",x"3a210f",x"351e0e",x"341e0e",x"321d0d",x"160f07",x"191007",x"211509",x"271909",x"251608",x"2b190a",x"29180a",x"26160a",x"2e1c0c",x"2b190b",x"2f1b0c",x"311d0c",x"361f0e",x"2f1c0c",x"331d0e",x"2f1b0d",x"2e1a0c",x"2c190b",x"2a180b",x"29180b",x"27170a",x"2b190b",x"27170b",x"301c0d",x"2f1b0c",x"24150a",x"28170b",x"2d1a0c",x"2a180b",x"2b190b",x"25160a",x"2e1b0c",x"25160a",x"27170b",x"2a190b",x"28180b",x"2b190b",x"2c1a0c",x"26160a",x"2a190b",x"2d1a0c",x"2c1a0c",x"2b190b",x"28170a",x"2b190b",x"2d1a0b",x"27170a",x"2c1a0c",x"2a190b",x"2c1a0c",x"2c1a0c",x"2c1a0c",x"2c1a0c",x"2b190c",x"2b190c",x"28180b",x"28170b",x"28170b",x"2a190b",x"28180b",x"28180b",x"29180b",x"27170b",x"2b190c",x"2c1a0c",x"251509",x"25150a",x"28160a",x"27160a",x"241409",x"231409",x"231409",x"241409",x"251509",x"251509",x"241509",x"231409",x"241509",x"27160a",x"2a180b",x"28170b",x"25160a",x"25160a",x"24150a",x"28180b",x"27170a",x"29180b",x"28170b",x"2c1a0c",x"26160a",x"26160a",x"25150a",x"2d1a0c",x"27170a",x"2a180b",x"2c1a0c",x"28170b",x"28170b",x"29180b",x"2a190b",x"2c1a0c",x"2c1a0c",x"29180b",x"29180b",x"2a190b",x"27170a",x"26150a",x"26160a",x"2a180b",x"2b190b",x"28170a",x"2c1a0b",x"2f1c0b",x"331e0c",x"2b190b",x"24160a",x"1d1208",x"26170a",x"281909",x"27180a",x"221509",x"1f1308",x"221608",x"241708",x"1e1209",x"23150a",x"27170a",x"1e1208",x"1e1209",x"211409",x"23150a",x"25160a",x"2b190b",x"311d0d",x"1d1208",x"261709",x"1d1108",x"1d1208",x"1e1209",x"1e1309",x"1d1208",x"1e1209",x"1f1309",x"1d1208",x"1d1208",x"180f07",x"1e1208",x"221409",x"201309",x"211409",x"28180b",x"2c1a0c",x"301c0d",x"2c1b0b",x"3c250e",x"452b10",x"36210b",x"2e1d0a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"37200f",x"150e07",x"191008",x"341d0d",x"3a200f",x"3b2210",x"3f2410",x"3e220f",x"3d220f",x"3f220f",x"3f230f",x"442611",x"442611",x"462712",x"412410",x"3f230f",x"412410",x"422511",x"452813",x"432611",x"472812",x"412510",x"402410",x"3f2310",x"3d220f",x"422511",x"3e230f",x"3c210e",x"3d220f",x"3c210f",x"391e0d",x"291307",x"3a200e",x"371f0e",x"3a1f0d",x"3b210e",x"3f2410",x"402410",x"3c210f",x"361e0e",x"3f2310",x"3e2310",x"3d220f",x"3f2410",x"3c210f",x"3a200e",x"3d220f",x"402310",x"412410",x"442612",x"422511",x"442713",x"462813",x"482a14",x"492a15",x"482914",x"472914",x"442612",x"422510",x"452712",x"492a14",x"482a14",x"361f0e",x"3c210f",x"150e07",x"341d0d",x"150e07",x"341c0b",x"371e0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2e18",x"4b2e18",x"5d4534",x"5a402f",x"60412e",x"583b28",x"60402a",x"644632",x"61422c",x"64412b",x"6d4e38",x"73523c",x"6f513d",x"694731",x"69452d",x"593a26",x"5b3923",x"5c3c29",x"583f2e",x"5d3d28",x"553623",x"583927",x"613e26",x"624029",x"644532",x"654936",x"5f4331",x"593d2c",x"5d4130",x"5e3f2c",x"5c3f2d",x"5c3d27",x"5d4130",x"593f2e",x"543c2d",x"553e2f",x"573f30",x"533e30",x"573f2f",x"573f2e",x"584030",x"5a3f2f",x"553d2e",x"543b2b",x"4b372a",x"503829",x"51392a",x"51392a",x"513829",x"45342a",x"513a2c",x"523b2d",x"554032",x"543d2e",x"5a4030",x"553f32",x"574032",x"503a2c",x"583f30",x"5a4233",x"553c2d",x"5b3f2e",x"5a3f2e",x"583f2f",x"5d4231",x"583e2d",x"5d4332",x"5e412e",x"5e412e",x"644430",x"5c3f2d",x"5c3f2d",x"5b3f2b",x"5c412f",x"63412c",x"64422c",x"61402c",x"5b3f2c",x"64422c",x"61412c",x"5d3f2b",x"5d3f2c",x"533a2a",x"4e3727",x"533b2c",x"523b2c",x"5a3c2a",x"4e3a2c",x"4e392a",x"503829",x"594130",x"523d2e",x"523c2d",x"593d2c",x"553c2d",x"543a29",x"573c29",x"5c3c2a",x"543a28",x"5e3f2c",x"62412c",x"5a3d2a",x"62432d",x"5e3f28",x"583c27",x"5f402a",x"5e422f",x"5d402c",x"54331b",x"150e07",x"150e07",x"150e07",x"150e07",x"4a2b14",x"150e07",x"24190f",x"24190e",x"24190f",x"2b1e12",x"25190e",x"251a0f",x"291c11",x"25190f",x"25190e",x"281b10",x"281b10",x"281b10",x"2a1d11",x"261a0f",x"2b1e12",x"2c1f12",x"2c1f12",x"2a1d11",x"342416",x"2b1e12",x"2d1f13",x"2e2114",x"2e2114",x"332416",x"302214",x"2f2114",x"2c1f13",x"312316",x"2b1e12",x"2f2115",x"322316",x"302215",x"332417",x"302215",x"332517",x"322316",x"312214",x"2f2114",x"312315",x"322316",x"302114",x"322315",x"302114",x"291c11",x"2a1c10",x"2f2113",x"312215",x"312215",x"342516",x"322315",x"2e2013",x"342416",x"322316",x"2e2014",x"352618",x"302215",x"302214",x"362618",x"2e2014",x"342517",x"2d2013",x"312316",x"352518",x"332417",x"312215",x"2e2014",x"2a1d12",x"2f2114",x"281c10",x"2b1e12",x"291c11",x"2e2013",x"2a1d11",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281509",x"281509",x"211106",x"2b190a",x"2c190b",x"160e07",x"181007",x"1b1107",x"1e1209",x"1e1208",x"251609",x"271709",x"2c1a0b",x"2b1a0b",x"2e1b0b",x"311c0c",x"2f1b0b",x"2d1a0b",x"311c0c",x"311c0b",x"2d1a0b",x"2b190b",x"27170b",x"2d1a0c",x"2d1a0c",x"2b190b",x"2f1c0d",x"29180b",x"241509",x"28170a",x"2b190b",x"25160a",x"2c1a0c",x"2b190b",x"26160a",x"29180a",x"27160a",x"28170a",x"26160a",x"27160a",x"28170a",x"28160a",x"26160a",x"29180b",x"28170b",x"2a180b",x"2a180b",x"28170a",x"27160a",x"241509",x"26160a",x"26160a",x"29180b",x"2a180b",x"2a190c",x"2d1b0d",x"2c1a0d",x"2e1c0d",x"2c1a0c",x"2a190c",x"28180b",x"2e1b0d",x"26170b",x"2a190c",x"2a190c",x"2c1a0c",x"2c1a0c",x"2d1b0c",x"2d1b0c",x"2b190c",x"26150a",x"27160a",x"27160a",x"2c190b",x"29180b",x"231409",x"241509",x"28170a",x"2a180b",x"27170a",x"27160a",x"221409",x"28170a",x"25150a",x"25160a",x"26160a",x"241509",x"221409",x"26160a",x"241509",x"251509",x"29180b",x"25150a",x"28170a",x"29180b",x"25150a",x"24150a",x"28170a",x"27160a",x"27160a",x"231409",x"26160a",x"231409",x"251509",x"1d1007",x"1f1108",x"25150a",x"201308",x"261509",x"25150a",x"211409",x"26160a",x"241509",x"251509",x"241509",x"231409",x"261609",x"261609",x"28170a",x"251609",x"231409",x"1c1108",x"261609",x"1f1308",x"231609",x"26180a",x"261709",x"251709",x"1f1308",x"221409",x"1f1209",x"26160a",x"1f1209",x"25160a",x"23150a",x"25160a",x"2a180b",x"251509",x"25160a",x"2a180a",x"1e1308",x"1d1208",x"1c1108",x"1d1108",x"1d1108",x"1d1208",x"1d1208",x"1e1209",x"1f1209",x"1c1108",x"1a1008",x"1d1108",x"1c1108",x"1d1108",x"211409",x"23150a",x"22150a",x"22150a",x"311d0d",x"35210d",x"3f270f",x"311d0a",x"36210c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"37200f",x"150e07",x"1f1309",x"321c0c",x"361d0d",x"351c0c",x"371e0d",x"3a200d",x"3a200d",x"3b200d",x"3b200e",x"3b200e",x"3b200d",x"381e0c",x"3a1f0d",x"381e0d",x"361d0c",x"391e0c",x"3a1f0d",x"3e220f",x"422410",x"3f230f",x"3f230f",x"3d210f",x"361e0d",x"3a200e",x"422611",x"442712",x"452813",x"452812",x"432611",x"452712",x"432712",x"402410",x"402410",x"432611",x"422611",x"3e230f",x"3c210e",x"3c210f",x"402411",x"482a14",x"462914",x"432712",x"482914",x"442713",x"442712",x"482a14",x"492a14",x"482a14",x"472913",x"442712",x"432611",x"452812",x"432611",x"422511",x"3f230f",x"3e220f",x"422510",x"472912",x"472913",x"442612",x"462812",x"38200e",x"2d190b",x"3d220f",x"150e07",x"351d0b",x"351d0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f311b",x"4f311b",x"5d4331",x"583e2d",x"60422d",x"60402a",x"5c3f2b",x"593c29",x"523827",x"5e412d",x"61432f",x"654734",x"68462f",x"5f3c26",x"5c3c2a",x"5f412f",x"513421",x"533623",x"593e2d",x"533625",x"563a28",x"5b3a25",x"543725",x"533a2a",x"593f2f",x"5c402e",x"593e2c",x"5f4434",x"573c2c",x"5a4131",x"5c4333",x"503a2c",x"543f31",x"543f30",x"4b3a2e",x"4c382b",x"4d382b",x"533b2d",x"583f30",x"593d2b",x"553e2f",x"553a2a",x"533c2d",x"543c2d",x"513c2e",x"573f30",x"573e2d",x"563f2f",x"583e2d",x"573f2e",x"5a4231",x"593e2c",x"523e31",x"5a4232",x"5a412f",x"553e2f",x"553f31",x"4e3a2d",x"573e2f",x"5a402f",x"573f2e",x"5a402f",x"60422f",x"5e412d",x"634632",x"563d2c",x"5f412d",x"5c4333",x"5c402e",x"5b3f2b",x"5d412e",x"5d422f",x"573b28",x"5a3d2b",x"523a2a",x"593e2d",x"5c3d29",x"573b28",x"62432e",x"5f402d",x"573927",x"5d3d29",x"583b28",x"4e3626",x"523828",x"593d2c",x"583f2d",x"573e2d",x"4e3829",x"50392a",x"583e2c",x"563e2e",x"4f3828",x"513a2a",x"614331",x"5e412e",x"5c3f2d",x"65452f",x"5e422e",x"62422c",x"60412c",x"573925",x"563926",x"553723",x"553b29",x"60412c",x"593e2b",x"5c3f2e",x"51311b",x"150e07",x"150e07",x"150e07",x"150e07",x"462913",x"150e07",x"291c11",x"22170d",x"23180e",x"24190e",x"2a1d11",x"24190e",x"23180e",x"25190e",x"281b10",x"251a0f",x"2c1f12",x"291c10",x"2f2115",x"2d1f13",x"281c10",x"322316",x"2e2114",x"2f2114",x"2f2114",x"2c1e12",x"2d1f13",x"312215",x"2f2114",x"2e2013",x"2d1f12",x"2c1e12",x"281b10",x"2e1f13",x"2e2013",x"2f2114",x"342517",x"2e2014",x"312215",x"312215",x"322416",x"302114",x"302215",x"322416",x"342416",x"312214",x"302114",x"2f2114",x"322316",x"352516",x"362719",x"332416",x"312214",x"2d2013",x"362719",x"2f2114",x"352517",x"322315",x"312215",x"2e2013",x"312315",x"342416",x"352517",x"2e1f12",x"2a1d11",x"322315",x"312215",x"342416",x"362618",x"2c1f13",x"2e2014",x"2f2114",x"2a1d12",x"2a1d11",x"2c1f13",x"302214",x"2d2013",x"2c1e12",x"281b10",x"2b1d11",x"2b1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1a0c",x"2d1a0c",x"2a190b",x"28180a",x"2a180a",x"160e07",x"170f07",x"180f07",x"190f08",x"1c1208",x"1a1008",x"1f1209",x"28180b",x"2c1b0b",x"29190b",x"2a190b",x"2b1a0b",x"2b190b",x"2c1a0b",x"2e1b0c",x"2b190b",x"29180b",x"27170a",x"27170a",x"1e1208",x"25160a",x"211409",x"211409",x"241509",x"27160a",x"2a180b",x"26160a",x"25150a",x"29180b",x"27170a",x"25160a",x"241509",x"25150a",x"231509",x"27160a",x"211409",x"28170a",x"25160a",x"24150a",x"26160a",x"26160a",x"27170a",x"29180b",x"28180b",x"27170b",x"27170b",x"28180b",x"28180b",x"2a190c",x"28180b",x"29180b",x"27160a",x"26160a",x"27170a",x"27170b",x"2a190b",x"27170b",x"25160a",x"24150a",x"27170b",x"26160a",x"26160a",x"26160a",x"28180b",x"241509",x"28170a",x"251509",x"251509",x"26160a",x"25150a",x"26160a",x"241509",x"25150a",x"211309",x"201308",x"221309",x"231409",x"211309",x"221409",x"211309",x"211309",x"211309",x"201208",x"221409",x"1f1208",x"201208",x"1f1208",x"1f1208",x"221409",x"241509",x"211309",x"1f1208",x"241509",x"201309",x"231409",x"1f1309",x"23150a",x"1f1309",x"25160a",x"1d1208",x"1f1309",x"1d1208",x"1b1108",x"1f1309",x"211409",x"241509",x"211309",x"221309",x"24150a",x"28170b",x"22150a",x"25160a",x"221409",x"28180b",x"25160a",x"1d1108",x"23150a",x"221409",x"24160a",x"1c1108",x"201409",x"211509",x"1c1107",x"170f07",x"170f07",x"1f1208",x"1f1208",x"191008",x"1e1208",x"24150a",x"1a1008",x"211409",x"201309",x"201309",x"1c1108",x"1b1108",x"1c1108",x"1d1208",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1d1208",x"180f08",x"1f1309",x"201309",x"201309",x"22150a",x"24160a",x"24150a",x"27180a",x"2a190a",x"37210d",x"36210c",x"311e0b",x"36210c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1f1309",x"321d0d",x"150e07",x"27170a",x"2e1a0b",x"28170a",x"29170a",x"2a180a",x"28170a",x"241409",x"261509",x"251409",x"241409",x"271509",x"2b170a",x"28160a",x"251509",x"27160a",x"26160a",x"2a180a",x"28160a",x"29170a",x"2d190b",x"2a180a",x"27160a",x"29170a",x"2a180b",x"2d1b0c",x"2d1b0c",x"321d0e",x"301c0d",x"331e0e",x"2f1b0d",x"301c0d",x"2f1c0d",x"2d1b0c",x"331e0e",x"311d0d",x"2f1c0d",x"2f1a0b",x"29170a",x"2c1a0c",x"301c0d",x"321d0e",x"2f1c0d",x"321d0d",x"301c0d",x"311c0d",x"2f1b0c",x"301c0d",x"301c0d",x"2d1a0b",x"321d0d",x"2f1b0c",x"2c1a0c",x"311c0d",x"301c0d",x"311c0d",x"311c0d",x"301c0d",x"39210f",x"341e0e",x"311c0d",x"301c0d",x"301c0d",x"321d0d",x"3b210f",x"150e07",x"361e0c",x"361e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2f1b",x"4c2f1b",x"5b3f2d",x"61412d",x"5d3f29",x"61412d",x"5a3e2a",x"5b412e",x"5a3b27",x"644734",x"634531",x"62442f",x"60402b",x"664732",x"593a26",x"5b3d28",x"593c2a",x"5a3b27",x"4d321f",x"543724",x"563a27",x"543b2b",x"593f2f",x"563b29",x"554031",x"594231",x"4e3a2e",x"564438",x"584134",x"584132",x"564134",x"553e31",x"513f33",x"594233",x"564032",x"584030",x"5c4232",x"543e2f",x"574032",x"5c4232",x"5c4332",x"5a4132",x"5e4332",x"5f4232",x"604534",x"5c4332",x"5f4534",x"604432",x"5b4232",x"614634",x"614531",x"634532",x"5f4331",x"543b2b",x"5f412c",x"5f422f",x"523d2f",x"563d2e",x"624736",x"5b412f",x"574030",x"614634",x"644632",x"604431",x"634633",x"5d4130",x"5a4130",x"5f4330",x"573c2a",x"573c2a",x"573e2f",x"5d3e28",x"583c28",x"5e402c",x"5d3e2a",x"573b28",x"60422d",x"573926",x"61412a",x"61412c",x"5c3d29",x"64422c",x"543826",x"553927",x"5b3e2c",x"664531",x"5b3e2c",x"5d3e2c",x"4f392a",x"563d2c",x"59402f",x"5b4130",x"5c4130",x"593f2e",x"5a3f2e",x"5c3e2a",x"5d3f2b",x"5b3e2b",x"503627",x"5e402e",x"5b3d2b",x"533826",x"583b29",x"60412c",x"5d3f2a",x"593b27",x"5b3e2a",x"4f392a",x"55341d",x"150e07",x"150e07",x"150e07",x"150e07",x"4a2b14",x"150e07",x"23180e",x"2a1e12",x"2b1e12",x"2a1d12",x"25190f",x"291c11",x"291c11",x"2a1d12",x"2c1e12",x"2b1e12",x"2d2014",x"2e2114",x"2f2014",x"2d1f13",x"291d11",x"2f2014",x"2e2114",x"291d11",x"322316",x"322316",x"2e2013",x"322416",x"2e2013",x"2c1e12",x"2b1d11",x"302214",x"342416",x"302114",x"342416",x"352617",x"312315",x"322316",x"312215",x"352618",x"362719",x"302215",x"322316",x"332416",x"352517",x"332417",x"342517",x"312316",x"362719",x"332417",x"332416",x"312316",x"342517",x"312215",x"2d1f13",x"322416",x"2f2114",x"312215",x"342416",x"322416",x"362618",x"2d1f12",x"322214",x"302214",x"312215",x"302114",x"2e2013",x"332416",x"352517",x"342517",x"2e2014",x"2f2115",x"2f2215",x"2e2014",x"312215",x"291c11",x"2f2114",x"2e2014",x"261a10",x"2d1f14",x"2d1f14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1008",x"1a1008",x"1c1108",x"160f07",x"160e07",x"160f07",x"170f07",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1e1208",x"23160a",x"24160a",x"26170a",x"25160a",x"231609",x"25170a",x"231509",x"221509",x"241509",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1309",x"201309",x"201309",x"1f1209",x"201309",x"201309",x"1f1309",x"1f1208",x"1f1209",x"211409",x"211409",x"211409",x"201309",x"211409",x"211409",x"211409",x"221409",x"211409",x"221409",x"211409",x"221409",x"211409",x"221409",x"221409",x"221409",x"221409",x"231509",x"26160a",x"27170b",x"27170b",x"27170b",x"27170b",x"26170a",x"26160a",x"27170b",x"27170b",x"27170b",x"27170b",x"25160a",x"25160a",x"26160a",x"26160a",x"25160a",x"25160a",x"25150a",x"241509",x"25150a",x"241509",x"241509",x"241509",x"211309",x"221409",x"201208",x"201208",x"201208",x"1f1108",x"1f1108",x"1f1208",x"1f1208",x"201308",x"201309",x"201308",x"201308",x"1f1208",x"1e1208",x"1d1208",x"1e1208",x"1d1108",x"1d1108",x"1c1108",x"1e1209",x"1e1309",x"1e1209",x"1d1209",x"1c1208",x"1d1208",x"1d1208",x"1c1108",x"1e1209",x"1c1108",x"1c1108",x"1c1208",x"1b1108",x"1b1108",x"1d1108",x"1e1309",x"1f1309",x"201309",x"201309",x"1f1309",x"201309",x"1e1209",x"1d1208",x"1e1209",x"201409",x"1e1308",x"201309",x"1b1108",x"1e1209",x"180f08",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160f07",x"170f07",x"191008",x"1c1108",x"1b1008",x"1c1108",x"1d1208",x"1e1208",x"1e1208",x"1f1209",x"1f1309",x"1f1309",x"1f1309",x"1e1208",x"1d1208",x"1b1108",x"191008",x"170f07",x"160e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"25160a",x"251709",x"2f1d0b",x"3b240d",x"38230c",x"33200b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"36200f",x"150e07",x"3e230f",x"40230f",x"3d210e",x"3f220f",x"3e220e",x"40230f",x"412410",x"422410",x"442611",x"422510",x"40230f",x"422410",x"40230f",x"40240f",x"422410",x"432510",x"442611",x"432510",x"402410",x"3e220e",x"3d220e",x"3e220e",x"3d220e",x"3e220f",x"3e220f",x"432611",x"482a13",x"482913",x"462712",x"472813",x"4b2b15",x"472813",x"3d210f",x"462812",x"492b14",x"4b2c15",x"4f2e17",x"4d2e16",x"4e2f16",x"4c2d16",x"4e2e16",x"4d2d15",x"4d2d16",x"4b2b15",x"4d2d16",x"4e2e17",x"4a2b15",x"4e2d16",x"502f17",x"4a2b15",x"4e2e17",x"4e2e16",x"482913",x"452611",x"482913",x"4a2a14",x"4a2a14",x"482913",x"422410",x"4a2b14",x"4d2d16",x"482a14",x"4c2d16",x"4a2a15",x"150e07",x"3e220e",x"361e0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d301c",x"4d301c",x"5b3f2e",x"63442f",x"5d3e29",x"5b3c28",x"583d2a",x"593b28",x"583b28",x"5b3f2b",x"5f412b",x"654531",x"61402a",x"5c3f2a",x"5d3d28",x"573b28",x"533420",x"533725",x"4c3424",x"4a3121",x"573e2e",x"50392a",x"563f31",x"594131",x"5a4638",x"564336",x"564235",x"564438",x"5d4738",x"5a4333",x"5b4537",x"5f4535",x"5c4332",x"5a4130",x"5e4332",x"5e4333",x"624533",x"5e4231",x"5f4331",x"5d4332",x"573f31",x"573f2f",x"533e2f",x"593f2f",x"5b4131",x"594132",x"5b402e",x"5a4130",x"5f4432",x"5b4230",x"664733",x"61432f",x"5f4331",x"5a4232",x"604432",x"5b402e",x"574030",x"644734",x"674731",x"614430",x"61432d",x"5c412e",x"5e422f",x"61432f",x"624431",x"654632",x"654835",x"664632",x"63442f",x"5e412e",x"61432e",x"5d412e",x"60422d",x"533c2c",x"573c2a",x"543b2a",x"5c3e2b",x"593c29",x"553a28",x"5a3c2a",x"5a3d28",x"5f3e2a",x"623f29",x"5c3d28",x"65452d",x"61422e",x"614029",x"5f402d",x"5a3e2d",x"543927",x"573d2b",x"59402e",x"553b28",x"583e2b",x"573e2d",x"563d2d",x"5e402c",x"614431",x"5c412e",x"5b412f",x"62432d",x"553b28",x"5a3e2b",x"593d2b",x"4b3526",x"483223",x"533b2b",x"503928",x"52331d",x"150e07",x"150e07",x"150e07",x"150e07",x"462813",x"150e07",x"261b10",x"291c11",x"2b1e12",x"2b1e12",x"2b1e12",x"2a1d12",x"2e2014",x"271c11",x"2c1f13",x"2f2115",x"322316",x"302216",x"322416",x"2d2014",x"2d2014",x"2e2115",x"2d1f13",x"312215",x"302114",x"302114",x"2e2013",x"332416",x"352517",x"2e2013",x"342516",x"352618",x"332416",x"2f2114",x"2d1e12",x"352517",x"332417",x"352618",x"352518",x"352517",x"342517",x"342517",x"372819",x"352517",x"372719",x"38281a",x"322416",x"342517",x"372719",x"322417",x"372819",x"3a2a1b",x"372719",x"362719",x"322315",x"2c1f12",x"302114",x"302114",x"312215",x"362718",x"362618",x"352517",x"322316",x"2d1f13",x"2d1f13",x"312215",x"291c10",x"2f2114",x"352618",x"2e2114",x"332417",x"2d1f13",x"2d2014",x"2f2115",x"2d2013",x"2c1f13",x"322416",x"2f2215",x"322416",x"2e2114",x"2e2114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"160e07",x"160f07",x"170e07",x"160e07",x"170f07",x"1d1208",x"1e1208",x"1b1108",x"1d1208",x"201509",x"211409",x"211509",x"221609",x"231509",x"231409",x"24160a",x"29190b",x"26170a",x"23150a",x"23150a",x"23150a",x"24160a",x"23150a",x"211409",x"1f1209",x"201309",x"211409",x"211409",x"201309",x"1e1208",x"201309",x"211409",x"211409",x"221409",x"211409",x"221409",x"211409",x"211409",x"211409",x"221409",x"211409",x"22150a",x"23150a",x"23150a",x"23150a",x"23150a",x"24150a",x"23150a",x"24160a",x"24160a",x"25160a",x"26170b",x"27170b",x"27170b",x"27170b",x"25150a",x"26160a",x"28170b",x"28170b",x"28180b",x"26160a",x"26160a",x"27170a",x"26160a",x"26160a",x"26160a",x"26160a",x"28170b",x"27170a",x"27170a",x"26160a",x"25150a",x"241509",x"241509",x"241509",x"231409",x"231409",x"221409",x"231409",x"231409",x"241509",x"241509",x"241509",x"231409",x"221409",x"231409",x"211309",x"211309",x"211309",x"211409",x"201309",x"201309",x"1f1208",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1c1108",x"1c1108",x"1d1208",x"1e1209",x"1f1309",x"201309",x"201409",x"201409",x"211409",x"211409",x"211409",x"22140a",x"201309",x"1f1309",x"1e1209",x"231609",x"1e1208",x"1e1308",x"201409",x"1c1107",x"170f07",x"170f07",x"170f07",x"160f07",x"170e07",x"170e07",x"170f07",x"170f07",x"191008",x"1a1008",x"1c1108",x"1d1208",x"1d1208",x"1e1208",x"1f1309",x"1f1309",x"201309",x"211409",x"201409",x"201309",x"1e1209",x"1d1208",x"1b1108",x"191008",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"191107",x"241708",x"2a1b09",x"38230c",x"36220b",x"38230c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1b1108",x"351f0e",x"150e07",x"3c210e",x"381c0c",x"3b200d",x"3d210e",x"41240f",x"422510",x"462712",x"452712",x"432611",x"422510",x"40220f",x"40220f",x"452812",x"4a2b14",x"482913",x"432510",x"3e210e",x"3c210e",x"3d210e",x"402410",x"462712",x"462812",x"452712",x"462812",x"452712",x"462712",x"4a2a13",x"4d2d16",x"4b2c15",x"492a14",x"4b2b15",x"4c2d16",x"492a14",x"482a14",x"482a14",x"4c2d16",x"4d2d16",x"482a15",x"4a2b15",x"4b2c15",x"4a2c15",x"502f17",x"4d2d15",x"472913",x"472812",x"462813",x"482913",x"4a2a13",x"472812",x"492a14",x"4d2d16",x"482913",x"523118",x"58361b",x"503018",x"492a13",x"472813",x"452813",x"482a13",x"482a14",x"4c2c15",x"492a14",x"462913",x"452712",x"150e07",x"351d0b",x"2f190a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50321e",x"50321e",x"67452e",x"69472e",x"64432e",x"61402a",x"67432c",x"65432b",x"654129",x"634028",x"603f2b",x"593d2b",x"5a3d2b",x"563825",x"543928",x"593b28",x"513827",x"523d2f",x"563e2f",x"503829",x"503a2b",x"554133",x"564031",x"523d2f",x"584132",x"584335",x"5e493b",x"594233",x"594436",x"5b4333",x"5d4535",x"5a4131",x"604534",x"664935",x"664936",x"604534",x"5c4131",x"5a4233",x"5f4535",x"5f4535",x"604432",x"664937",x"624836",x"614634",x"624633",x"614634",x"5b412f",x"604535",x"644936",x"654632",x"654735",x"614431",x"654734",x"624533",x"674734",x"604734",x"624532",x"5f4533",x"664834",x"664936",x"674b38",x"664834",x"624531",x"614735",x"614433",x"5d412f",x"5e4231",x"654733",x"634432",x"5f412d",x"664631",x"5e412f",x"634430",x"63422c",x"583d2b",x"5a3d2b",x"583b27",x"5e3f2b",x"5e3e29",x"5a3c29",x"5e3f2a",x"5e3f2a",x"603f2c",x"60402b",x"5f3e29",x"5e3f2c",x"65442f",x"644731",x"664834",x"60432d",x"59402e",x"5a4130",x"553d2d",x"593f2c",x"5f422e",x"5d412f",x"5d4230",x"583f2d",x"5b3f2c",x"5f422e",x"61432e",x"513827",x"4c3729",x"583c29",x"483324",x"563b2a",x"513b2a",x"473325",x"56351e",x"150e07",x"150e07",x"150e07",x"150e07",x"472913",x"1a1108",x"25190f",x"2b1e12",x"2a1d11",x"23180e",x"251a0f",x"2a1d11",x"281c10",x"291c11",x"2a1d11",x"2a1d12",x"2a1d11",x"2b1e12",x"2b1e12",x"302214",x"2a1d11",x"2f2114",x"2d1f12",x"281c10",x"2d2013",x"332416",x"312215",x"312215",x"312316",x"2e2013",x"2e2013",x"2e2013",x"302114",x"2f2114",x"2c1e12",x"2d1f12",x"312215",x"342416",x"312215",x"312316",x"302214",x"2d2013",x"332416",x"322315",x"322316",x"2d1f12",x"332416",x"322416",x"322315",x"312215",x"312316",x"322416",x"312214",x"2f2114",x"312215",x"2e2013",x"352617",x"332416",x"322316",x"322416",x"332416",x"312215",x"312215",x"312214",x"2c1e12",x"312215",x"2e2013",x"291c11",x"2c1f12",x"2e1f13",x"312215",x"2d1f13",x"2c1f12",x"2b1e12",x"2e2013",x"2e2013",x"2c1f12",x"2b1e11",x"2c1e12",x"2a1d12",x"2a1d12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"180f07",x"170f07",x"170f07",x"170f07",x"1b1008",x"1e1308",x"221509",x"1d1208",x"1e1209",x"1f1309",x"211409",x"221409",x"211409",x"211409",x"241609",x"241609",x"241609",x"221409",x"221409",x"24150a",x"25160a",x"231409",x"25160a",x"26170b",x"25160a",x"221409",x"221409",x"221509",x"221409",x"221409",x"22140a",x"221509",x"211409",x"211409",x"201309",x"201309",x"211409",x"23150a",x"24150a",x"24160a",x"23150a",x"23150a",x"24160a",x"24160a",x"24160a",x"24160a",x"24160a",x"25160a",x"25160a",x"25160a",x"26170b",x"27170b",x"28170b",x"28170b",x"29180b",x"29190b",x"2b190c",x"2a190b",x"29180b",x"27170a",x"27170a",x"27170a",x"27160a",x"26160a",x"27170a",x"26160a",x"26160a",x"27170a",x"251509",x"251509",x"251509",x"241509",x"231409",x"231409",x"221309",x"221409",x"231409",x"241509",x"251509",x"25160a",x"25160a",x"241509",x"231409",x"221309",x"231409",x"25160a",x"24150a",x"231409",x"201308",x"1f1208",x"1e1208",x"1f1208",x"1f1308",x"1f1209",x"1f1309",x"1e1209",x"1d1208",x"1d1108",x"1d1108",x"1d1208",x"1d1209",x"1d1208",x"1d1208",x"1d1208",x"1c1208",x"1c1108",x"1c1108",x"1d1208",x"1d1209",x"1e1309",x"1e1309",x"201309",x"211409",x"211409",x"221409",x"221409",x"211409",x"211409",x"201309",x"1f1309",x"1d1208",x"211408",x"1f1308",x"1d1208",x"1c1108",x"211509",x"1a1108",x"170f07",x"180f07",x"160f07",x"170e07",x"170f07",x"170f07",x"170f07",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1f1209",x"201409",x"211409",x"211409",x"211409",x"211409",x"211409",x"1f1309",x"1e1209",x"1b1108",x"1a1008",x"180f08",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231608",x"2b1b09",x"2b1b09",x"32200a",x"321f0b",x"2f1c0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211309",x"38200f",x"150e07",x"28160a",x"2c180a",x"29170a",x"29170a",x"2a170a",x"2d190b",x"301c0c",x"311c0c",x"321c0d",x"301c0c",x"301b0c",x"301b0c",x"2f1b0b",x"341d0d",x"321d0c",x"2f1a0b",x"2d190b",x"301c0d",x"2b190b",x"351f0f",x"351e0e",x"361e0e",x"3a2110",x"341e0e",x"301b0c",x"2f1a0b",x"361f0f",x"341e0e",x"311d0d",x"2f1c0c",x"311b0c",x"331d0d",x"2c190b",x"311b0c",x"321c0d",x"2f1b0c",x"311d0d",x"2b190b",x"321d0e",x"2d1a0c",x"331d0e",x"351e0e",x"331d0d",x"25160a",x"28170a",x"2f1b0c",x"27160a",x"321d0d",x"2f1b0d",x"37200f",x"361f0f",x"311c0d",x"37200f",x"38210f",x"341f0e",x"331d0e",x"301c0d",x"38200f",x"36200f",x"2f1b0c",x"2f1b0c",x"331e0e",x"38210f",x"3f2511",x"150e07",x"3a200d",x"361e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50321e",x"50321e",x"61422f",x"5b3f2a",x"5e3d27",x"583a28",x"5f412c",x"61422e",x"5e3d28",x"573722",x"593a27",x"5e402d",x"5f3f2a",x"573a29",x"60412d",x"523826",x"493223",x"523524",x"4d3729",x"4c3628",x"563f31",x"564335",x"533c2c",x"574538",x"4f3e33",x"523f31",x"574538",x"5c483a",x"584435",x"574131",x"584132",x"614533",x"604332",x"5b4130",x"634532",x"5b3f2e",x"593e2d",x"61432f",x"60422f",x"63432d",x"5f412e",x"5a3e2b",x"61422e",x"5e422f",x"5e412d",x"5b4030",x"5b4130",x"5b4130",x"5c4230",x"5a3f2e",x"583d2b",x"573f2f",x"583d2c",x"573d2d",x"5b3e2c",x"593f2f",x"593b28",x"573d2c",x"5b3e2a",x"61412c",x"66432e",x"593f2e",x"5e422f",x"5d402d",x"664733",x"5e4333",x"634632",x"684935",x"614431",x"604533",x"644733",x"5d402e",x"614430",x"624530",x"63442f",x"62432d",x"5c3e2b",x"664530",x"66442d",x"5f3f2b",x"5e3e29",x"603f2a",x"66432c",x"66432b",x"6a472f",x"62422a",x"61402a",x"603f2a",x"5a3f2e",x"5f4230",x"634531",x"5e4331",x"594233",x"573f30",x"5c4332",x"543c2d",x"594132",x"5a3f2e",x"5c412f",x"553c2c",x"573d2b",x"4c3729",x"4d3728",x"4a3425",x"4f3626",x"4a3527",x"463428",x"403429",x"53341f",x"150e07",x"150e07",x"150e07",x"150e07",x"452711",x"1c1208",x"23180e",x"291c11",x"2b1d12",x"2b1e12",x"251a0f",x"291c11",x"291c11",x"291d11",x"2d1f13",x"2a1d11",x"2e2014",x"2a1d11",x"2c1f13",x"2e2014",x"302215",x"2d1f13",x"2e2014",x"291d11",x"2a1d12",x"2b1d12",x"2a1d11",x"312215",x"302215",x"312316",x"2e2014",x"352517",x"342417",x"352618",x"322316",x"342417",x"2d1f13",x"342517",x"2f2114",x"342517",x"312215",x"352517",x"312316",x"342517",x"2a1d11",x"312215",x"2e2014",x"2c1e12",x"342517",x"2d1f13",x"312215",x"352517",x"332416",x"2d1f13",x"2e2014",x"2d1f13",x"322416",x"332315",x"322315",x"372718",x"362719",x"352619",x"342517",x"352517",x"322316",x"332416",x"312215",x"2f2114",x"302114",x"322416",x"2f2114",x"2d1f13",x"2d1f13",x"2d1f13",x"2b1e12",x"2d1f13",x"2a1d11",x"2b1e12",x"2e2114",x"291c11",x"291c11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"191007",x"180f08",x"221509",x"211409",x"1e1308",x"1d1208",x"1f1309",x"201309",x"201309",x"211409",x"241609",x"241509",x"241509",x"231509",x"23150a",x"24150a",x"24160a",x"25160a",x"24150a",x"26160b",x"25160a",x"25160a",x"24150a",x"23150a",x"23150a",x"24150a",x"231409",x"211409",x"23150a",x"23150a",x"23150a",x"23150a",x"23150a",x"211309",x"211409",x"211409",x"221409",x"23150a",x"23150a",x"231509",x"24150a",x"24160a",x"24150a",x"24150a",x"24160a",x"25160a",x"241509",x"26160a",x"26170a",x"27170a",x"27170b",x"27170b",x"27170a",x"27170b",x"26160a",x"27170a",x"26160a",x"241509",x"26160a",x"241509",x"26160a",x"27160a",x"241509",x"27170a",x"26160a",x"251509",x"241509",x"241509",x"261609",x"251509",x"241509",x"231409",x"221308",x"221309",x"231409",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"25150a",x"241509",x"241509",x"25160a",x"221409",x"211309",x"221409",x"221409",x"211409",x"221409",x"1f1309",x"1f1309",x"201309",x"1e1208",x"1d1108",x"1d1108",x"1e1209",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1b1108",x"1c1108",x"1d1108",x"1d1208",x"1e1209",x"201309",x"201309",x"201309",x"211409",x"211409",x"23150a",x"201309",x"201309",x"201309",x"1f1309",x"1f1309",x"21150a",x"1e1308",x"201409",x"231609",x"1d1208",x"191007",x"170f07",x"170f07",x"171007",x"180f07",x"181007",x"170f07",x"191008",x"1a1108",x"1c1108",x"1d1208",x"1d1108",x"1d1108",x"1e1208",x"1f1209",x"201309",x"211409",x"201309",x"201309",x"201309",x"1e1209",x"1c1108",x"1a1108",x"191008",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"2b1b09",x"2f1e0a",x"2b1b09",x"2e1c0b",x"2c1c0a",x"2c1b0a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"341e0e",x"150e07",x"231409",x"311b0b",x"3d210e",x"40230f",x"3f240f",x"402310",x"3e220f",x"442611",x"412410",x"412410",x"40220f",x"40240f",x"452712",x"432611",x"422511",x"412410",x"412410",x"3e230f",x"412410",x"3f2410",x"402410",x"452611",x"3e230f",x"432711",x"402411",x"432611",x"432611",x"432611",x"462813",x"452813",x"452813",x"492a14",x"3f2410",x"3e220f",x"3a1f0e",x"3f2410",x"3a210f",x"3b220f",x"3e2310",x"3f2410",x"432813",x"462812",x"452712",x"432711",x"462813",x"472913",x"472a14",x"422611",x"4c2d16",x"4d2e16",x"482a14",x"402410",x"412410",x"482914",x"3f2410",x"432510",x"432611",x"492b14",x"492b14",x"442813",x"492a14",x"3d2310",x"2b190b",x"39200e",x"150e07",x"361e0c",x"2e190a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"51341f",x"51341f",x"573d2c",x"593f2d",x"5f3e27",x"64442f",x"5e3d28",x"62422c",x"63432e",x"62422e",x"624029",x"563825",x"5e3e28",x"67452f",x"5d3e28",x"543826",x"4e3423",x"4f3525",x"4f3625",x"553c2d",x"573e2d",x"594232",x"5a4334",x"513e31",x"594336",x"554134",x"594336",x"5c4738",x"594436",x"5c4536",x"5c4535",x"5e4637",x"644937",x"614838",x"634837",x"634835",x"574234",x"5e4433",x"604637",x"5d4231",x"604634",x"634736",x"614634",x"614432",x"614735",x"5d4231",x"5c4333",x"5b4332",x"574233",x"5f4533",x"5c4535",x"5e4230",x"644835",x"584031",x"594233",x"5b4434",x"5b4536",x"5b4435",x"5d4333",x"5f4331",x"694b37",x"644936",x"60432f",x"5c412f",x"5b4333",x"604330",x"694b36",x"654835",x"5c3f2d",x"644733",x"62432f",x"5e422f",x"573f2e",x"5d4230",x"593e2d",x"523829",x"593d2c",x"62432c",x"62432e",x"64432d",x"5f3f2a",x"5b3e2a",x"5f3f28",x"5e3e2a",x"563926",x"573b2a",x"5b3c28",x"62412b",x"573c2b",x"51392a",x"583d2d",x"563f31",x"5d412f",x"5d4230",x"573f2f",x"584234",x"4e3c2f",x"553e2f",x"553e2f",x"543d2e",x"4c382a",x"4d392b",x"4f392b",x"3e3227",x"3c2f25",x"5a3c2a",x"503b2d",x"4c3b2e",x"563620",x"150e07",x"150e07",x"150e07",x"150e07",x"482913",x"1c1208",x"251a0f",x"23180e",x"261b10",x"24190e",x"2a1d11",x"312216",x"2c1f12",x"2f2115",x"2e2114",x"2c1f13",x"322416",x"2e2115",x"322316",x"362719",x"302215",x"2f2115",x"342518",x"342517",x"322316",x"312215",x"312215",x"322316",x"342517",x"322416",x"332417",x"2f2114",x"352618",x"332416",x"332416",x"2e2014",x"2e2013",x"322316",x"312215",x"322316",x"332417",x"352517",x"342517",x"332417",x"332416",x"352618",x"352518",x"332417",x"302214",x"3a2a1b",x"352518",x"332417",x"2f2215",x"312216",x"2f2115",x"2e2013",x"342416",x"342416",x"312215",x"322316",x"362618",x"302215",x"362719",x"322316",x"362719",x"302215",x"332416",x"2d1f13",x"322316",x"322316",x"2e2014",x"2f2114",x"2e2014",x"2c1f12",x"2c1f12",x"312216",x"2c1f12",x"2d1f13",x"2e2014",x"2c1f13",x"2c1f13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"1b1107",x"170f07",x"1a1108",x"271909",x"201408",x"1d1208",x"1e1208",x"211409",x"201309",x"221509",x"26170a",x"231509",x"28180a",x"25160a",x"24150a",x"24150a",x"26170b",x"25160a",x"231509",x"221409",x"24160a",x"231409",x"211309",x"231409",x"24150a",x"24160a",x"24150a",x"23150a",x"23150a",x"231509",x"211309",x"1f1208",x"201208",x"211309",x"211409",x"1f1208",x"1e1208",x"1f1208",x"201308",x"221409",x"23150a",x"221409",x"221409",x"221409",x"221409",x"231509",x"231509",x"24150a",x"25150a",x"25150a",x"25150a",x"26160a",x"26160a",x"28180b",x"29180b",x"28170b",x"27170a",x"27170a",x"29180b",x"28170b",x"28170a",x"27170a",x"28170b",x"29180b",x"27170a",x"27160a",x"27160a",x"26160a",x"26160a",x"26150a",x"241409",x"231409",x"241509",x"26160a",x"25150a",x"25150a",x"26160a",x"26160a",x"26160a",x"231409",x"231409",x"251509",x"25150a",x"24150a",x"241509",x"221409",x"221409",x"201309",x"201309",x"201309",x"1f1208",x"1e1208",x"1e1208",x"1f1309",x"1d1208",x"1d1108",x"1d1208",x"1d1208",x"1d1208",x"1d1208",x"1d1208",x"1c1108",x"1b1008",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1e1208",x"1e1209",x"201409",x"211409",x"201309",x"221409",x"221409",x"211409",x"221509",x"221409",x"1f1309",x"201409",x"23150a",x"211409",x"1d1208",x"1b1108",x"1c1208",x"1b1107",x"181007",x"160f07",x"170f07",x"180f07",x"160f07",x"170f07",x"180f08",x"191008",x"1a1008",x"1a1008",x"1c1108",x"1d1208",x"1d1108",x"1c1108",x"1d1108",x"1d1108",x"1f1208",x"201309",x"1f1209",x"1d1108",x"1c1108",x"1a1008",x"191008",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1308",x"2b1b09",x"261809",x"261809",x"2c1b0a",x"241608",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"3a2210",x"150e07",x"1c1108",x"3a1f0d",x"321b0c",x"381e0d",x"371e0c",x"371e0c",x"3a200e",x"3b200e",x"3c200d",x"3f230f",x"442611",x"412410",x"412410",x"3f2410",x"412411",x"422511",x"452712",x"422611",x"412410",x"3f230f",x"412511",x"452812",x"412410",x"3f2410",x"3e2310",x"412410",x"391e0d",x"361c0c",x"321a0b",x"381d0c",x"381e0d",x"3f2410",x"3d2310",x"412511",x"3f2310",x"351d0d",x"351d0d",x"321b0c",x"371e0d",x"391f0d",x"3b200e",x"391f0d",x"3d220f",x"3c210e",x"3d210f",x"3f220f",x"39200e",x"402511",x"482a14",x"472a14",x"432713",x"452914",x"4a2d15",x"432712",x"432712",x"452712",x"3f2410",x"422712",x"3b210f",x"462812",x"331d0d",x"3c210f",x"150e07",x"2e1a0b",x"150e07",x"3c210e",x"311b0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533520",x"533520",x"523928",x"543927",x"533a2a",x"60402c",x"5c3d29",x"62412c",x"60422e",x"583b28",x"563a28",x"593c28",x"533828",x"4a3223",x"553725",x"553c2c",x"513727",x"573a28",x"543a29",x"5b402f",x"5b4333",x"5d4333",x"543f32",x"533f32",x"533f32",x"544236",x"574234",x"584335",x"5c4537",x"5c4434",x"5f4433",x"5e4737",x"5d4535",x"5a4334",x"604736",x"5d4433",x"5a4334",x"634633",x"644836",x"5b4132",x"634532",x"6b4c37",x"644735",x"5f4231",x"5d4332",x"5e4333",x"5a4334",x"554033",x"543f33",x"533d30",x"563e30",x"543b2d",x"5f4432",x"5e4230",x"5b4130",x"583f30",x"563c2b",x"553e2f",x"543d2e",x"563d2d",x"563d2e",x"563c2c",x"573c2b",x"513829",x"563d2d",x"543b2b",x"5d4332",x"5c4334",x"604534",x"654733",x"634836",x"694934",x"60432f",x"5b402e",x"583c28",x"593f2d",x"5b3e2b",x"603f29",x"5d3e28",x"5e3f2a",x"543927",x"503624",x"523624",x"523624",x"5a3a25",x"5e3d27",x"573824",x"5a3d29",x"543726",x"513727",x"543a2a",x"553a29",x"61422e",x"5c402d",x"503c2e",x"45352a",x"4c392b",x"4f392b",x"533a2a",x"433226",x"4d382b",x"453225",x"413127",x"533a2a",x"392f26",x"4b372a",x"4b3729",x"4b3a2f",x"593a23",x"150e07",x"150e07",x"150e07",x"150e07",x"452711",x"1a1107",x"281c10",x"281c11",x"2a1d11",x"281c10",x"251a0f",x"2c1e12",x"2b1e12",x"2d1f13",x"2b1e13",x"2e2114",x"2f2115",x"2d1f13",x"302215",x"2d1f12",x"322315",x"2f2014",x"312214",x"2b1d11",x"2d1e12",x"2e1f12",x"312114",x"2e2013",x"302013",x"302114",x"392819",x"352517",x"342416",x"2d2013",x"312316",x"342517",x"322316",x"352618",x"362618",x"38281a",x"342517",x"322316",x"2e2013",x"2e1f13",x"342416",x"372719",x"342518",x"322417",x"342517",x"332517",x"332417",x"312215",x"2d1f12",x"2f2014",x"2e2013",x"2a1d11",x"2a1d11",x"2e1f12",x"2c1e11",x"312214",x"2d1e12",x"302114",x"352517",x"342416",x"312215",x"322316",x"342517",x"382819",x"382719",x"2d1f13",x"2d2013",x"302215",x"2e2013",x"2c1e12",x"312215",x"312214",x"2d2013",x"2a1e12",x"2b1e13",x"2f2115",x"2f2115",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"180f07",x"191007",x"1d1208",x"1d1108",x"1a1108",x"221509",x"1e1308",x"1c1108",x"1d1108",x"1e1108",x"231508",x"201308",x"231508",x"26160a",x"211309",x"231409",x"24150a",x"26160a",x"25160a",x"26160a",x"26170b",x"24150a",x"24150a",x"24150a",x"231509",x"25160a",x"221409",x"23150a",x"221409",x"221409",x"211309",x"201208",x"221409",x"221409",x"221409",x"211409",x"201308",x"211309",x"211309",x"201309",x"221409",x"221409",x"221409",x"231409",x"221409",x"231409",x"231509",x"231409",x"231409",x"241509",x"25160a",x"27170a",x"27170a",x"27160a",x"26160a",x"26160a",x"27160a",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"241509",x"251509",x"26160a",x"26160a",x"27170a",x"27170a",x"26160a",x"26160a",x"251509",x"241509",x"231409",x"231409",x"231409",x"231409",x"241509",x"231409",x"241409",x"26160a",x"26160a",x"25150a",x"25150a",x"25160a",x"241509",x"231409",x"24150a",x"231509",x"201309",x"211409",x"201409",x"1f1309",x"1d1108",x"1e1208",x"1d1208",x"1c1108",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"1f1309",x"1f1309",x"201309",x"1e1309",x"201408",x"1f1308",x"211409",x"191008",x"1b1107",x"191007",x"170f07",x"160f07",x"180f07",x"160e07",x"160f07",x"170f07",x"180f07",x"1a1008",x"1c1108",x"1d1108",x"1d1208",x"1d1108",x"1d1208",x"1e1208",x"1e1208",x"1f1309",x"1f1309",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"191008",x"180f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1e1308",x"241608",x"251809",x"241609",x"221509",x"1f1409",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"38210f",x"150e07",x"271609",x"2a170a",x"2a170a",x"231409",x"2d190b",x"3b210e",x"381f0d",x"311a0b",x"341c0c",x"351d0d",x"381f0e",x"331c0c",x"331c0c",x"361e0d",x"351d0d",x"3e220f",x"381f0e",x"3b210f",x"3b210f",x"341c0d",x"38200e",x"3a200f",x"3b210f",x"331c0c",x"3c2310",x"3b200e",x"402511",x"3d2411",x"38200f",x"3c2310",x"3c2210",x"37200f",x"3b2311",x"3d2311",x"412612",x"422712",x"3a2210",x"3a200f",x"39200e",x"3a210f",x"3d2310",x"3a210f",x"3b200e",x"3a210f",x"3a200e",x"39200e",x"39200f",x"3e2411",x"3d2411",x"3e2310",x"3d2310",x"361e0d",x"341c0c",x"361d0d",x"361e0d",x"361e0d",x"331c0c",x"351d0d",x"321c0c",x"3c210e",x"231409",x"311b0c",x"371f0e",x"150e07",x"1c1108",x"402410",x"3b2210",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482f1d",x"482f1d",x"593f2d",x"553a29",x"5d412f",x"593c28",x"563c2a",x"5f412e",x"543927",x"563b2a",x"523827",x"523726",x"543826",x"4f3626",x"52392a",x"583c2b",x"5f3e29",x"5a3e2a",x"583c2b",x"563e2f",x"513728",x"553c2d",x"543928",x"543827",x"4f3526",x"543826",x"583e2d",x"50392c",x"584132",x"5a4131",x"604737",x"5c4637",x"5a4335",x"5d4231",x"5a4233",x"604433",x"63442f",x"60432f",x"5e402d",x"5b4030",x"5d402d",x"60422d",x"61412d",x"5e402d",x"60432f",x"523b2c",x"5f4330",x"5e412d",x"5d412f",x"5d4230",x"5f422e",x"5e4330",x"654733",x"614532",x"654733",x"65452e",x"5b4231",x"5a4030",x"593f2d",x"604432",x"634632",x"644735",x"5b4231",x"5a402f",x"553c2d",x"5f4535",x"5e4636",x"614432",x"5f4432",x"644a37",x"614533",x"624330",x"553b2b",x"583e2d",x"563d2d",x"583b2a",x"563b2a",x"523827",x"523828",x"4d3424",x"513726",x"4f3424",x"503523",x"563925",x"593c29",x"60412b",x"553824",x"5b3e2c",x"533928",x"573b2a",x"543927",x"5f3f2a",x"604330",x"5a4131",x"543f31",x"513e31",x"563f30",x"4c3a2c",x"4e392b",x"4b382b",x"4d3a2e",x"513b2d",x"513a2a",x"3d3229",x"4b382a",x"3d332b",x"4b3729",x"4b3a2d",x"4f3320",x"150e07",x"150e07",x"150e07",x"150e07",x"432611",x"191007",x"281b10",x"2c1f13",x"2b1e13",x"2f2114",x"2c1f13",x"2b1e12",x"302215",x"2e2114",x"312316",x"302215",x"322416",x"2f2114",x"372719",x"302114",x"322316",x"322316",x"2e2013",x"2d1f12",x"2e2012",x"322315",x"342416",x"342416",x"362617",x"392819",x"342517",x"372719",x"302114",x"302215",x"342517",x"322316",x"372719",x"39291b",x"362719",x"39291b",x"322316",x"332417",x"372719",x"342517",x"372719",x"39291a",x"342517",x"322416",x"372719",x"352618",x"302215",x"2c1e12",x"322316",x"312215",x"2f2113",x"332214",x"2f2113",x"342416",x"2e2013",x"342416",x"2f2114",x"352517",x"372719",x"372719",x"332316",x"2e2014",x"362719",x"352518",x"332517",x"352718",x"3a2a1b",x"302216",x"322316",x"2f2114",x"2e2014",x"2f2115",x"302215",x"302215",x"2d2014",x"312315",x"312315",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"160e07",x"150e07",x"160f07",x"160e07",x"170f07",x"211509",x"1e1208",x"1f1308",x"201308",x"1f1308",x"211408",x"201309",x"221409",x"241509",x"241609",x"241509",x"231609",x"241609",x"24150a",x"25160a",x"24150a",x"24150a",x"221409",x"211309",x"211309",x"211309",x"211309",x"211309",x"221409",x"201309",x"201309",x"201309",x"201309",x"221409",x"24150a",x"25160a",x"24160a",x"24150a",x"23150a",x"221409",x"221409",x"221409",x"231509",x"231509",x"24150a",x"24150a",x"23150a",x"231509",x"24150a",x"24150a",x"241509",x"24150a",x"26160a",x"26160a",x"25160a",x"26160a",x"27170a",x"27170a",x"28170a",x"28170b",x"27160a",x"26160a",x"251509",x"251509",x"241509",x"241409",x"241509",x"241509",x"26160a",x"27170a",x"27160a",x"26160a",x"251509",x"241509",x"221409",x"231409",x"241509",x"241509",x"251509",x"241509",x"211208",x"231409",x"241509",x"241509",x"241509",x"221309",x"221409",x"221409",x"221409",x"24150a",x"221409",x"221409",x"201309",x"1f1208",x"201309",x"201309",x"1e1208",x"1f1309",x"1e1209",x"1e1209",x"1e1209",x"1e1209",x"1d1208",x"1d1208",x"1d1208",x"1d1208",x"1d1209",x"1d1208",x"1e1209",x"1e1209",x"1d1208",x"1d1208",x"1e1208",x"1f1309",x"1f1309",x"1f1309",x"201309",x"201309",x"1f1209",x"201309",x"201409",x"211409",x"1f1309",x"1d1208",x"1f1308",x"241609",x"1e1209",x"180f07",x"170f07",x"180f07",x"160f07",x"160e07",x"170f07",x"170f07",x"160e07",x"170f07",x"191008",x"1b1108",x"1c1108",x"1d1209",x"1f1209",x"1e1208",x"1e1208",x"1f1208",x"1f1309",x"201309",x"201309",x"1f1309",x"1e1208",x"1d1208",x"1c1108",x"1a1008",x"180f08",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"211508",x"231608",x"1f1408",x"211508",x"231509",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"3b2311",x"150e07",x"1c1108",x"311c0d",x"301c0c",x"2e1b0c",x"301c0c",x"3b210e",x"361d0c",x"341c0c",x"39200e",x"3b210f",x"3f2410",x"412410",x"3f2410",x"3b210f",x"3f2411",x"3e2310",x"3f2310",x"3e2310",x"3b220f",x"3b210f",x"3e2310",x"3d2310",x"3a200e",x"3e2310",x"39200e",x"371e0d",x"371e0d",x"39200e",x"3b210f",x"351d0d",x"38200e",x"3d2310",x"442813",x"3c210f",x"3f2411",x"432712",x"3a200f",x"341c0c",x"3b210f",x"3f2411",x"402511",x"371e0d",x"3c220f",x"3d220f",x"3f2310",x"3b2310",x"402512",x"402512",x"432713",x"3f2511",x"402411",x"402511",x"3f2410",x"3f2410",x"3f2410",x"3d2310",x"3e2310",x"3d2310",x"3c210f",x"432712",x"150e07",x"2e1a0b",x"301b0c",x"341e0d",x"2d1a0b",x"412511",x"371f0e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e321f",x"4e321f",x"4b3a2e",x"5d412f",x"5e402b",x"64442f",x"543b2b",x"523727",x"4e3526",x"4a3426",x"513828",x"4f3424",x"543724",x"503523",x"563928",x"5b3d2b",x"5d3e2b",x"553c2b",x"5f4332",x"5a402f",x"574031",x"5f4332",x"5c4231",x"5b4131",x"604330",x"624736",x"614332",x"5d402f",x"5e4331",x"5a4131",x"634837",x"654a39",x"614837",x"5b4333",x"634b3a",x"664b39",x"664a37",x"684b38",x"5f4534",x"654b3a",x"684c3a",x"644a39",x"624837",x"604738",x"5a4334",x"544133",x"564132",x"5e4433",x"604534",x"5c4433",x"5d4535",x"634733",x"5e4535",x"634632",x"5f4432",x"5c4230",x"624734",x"543d2f",x"594132",x"624531",x"654633",x"5c3f2d",x"5e4332",x"614532",x"5b402f",x"5c412f",x"664835",x"644734",x"614533",x"624532",x"654835",x"5c4231",x"5f422f",x"58402f",x"5f4330",x"593b28",x"533826",x"583b27",x"553926",x"593c28",x"543724",x"4a3223",x"573826",x"573a28",x"523726",x"523625",x"583a26",x"563926",x"5a3c28",x"553b29",x"533928",x"5b3e2b",x"5a3e2b",x"4e3b2e",x"513b2b",x"5a4131",x"563f2f",x"503d30",x"49382c",x"523d2e",x"463326",x"563b29",x"48372a",x"3d3229",x"49382d",x"423429",x"533a2a",x"392e26",x"563722",x"150e07",x"150e07",x"150e07",x"150e07",x"422611",x"191007",x"2d2012",x"23170d",x"2d1f13",x"2a1d12",x"291c11",x"2c1f13",x"2c1f13",x"2c1e12",x"302215",x"2e2014",x"352517",x"332416",x"2f2114",x"312114",x"2f2013",x"322315",x"302114",x"2e2013",x"2f2113",x"332315",x"2d1f12",x"322315",x"382819",x"362517",x"362617",x"332416",x"332416",x"382819",x"3b2a1b",x"332417",x"322316",x"352617",x"342517",x"302114",x"342517",x"2e2013",x"312315",x"39291a",x"332416",x"312214",x"332416",x"352517",x"332416",x"332416",x"322315",x"322315",x"312214",x"2d1f12",x"2c1e12",x"302114",x"2b1d11",x"2f2113",x"332316",x"322315",x"342417",x"342416",x"382719",x"352618",x"362718",x"362619",x"38281a",x"352517",x"362617",x"2b1e12",x"342517",x"322315",x"2b1e12",x"2c1f12",x"2d1f13",x"2e2114",x"302215",x"312214",x"2a1d11",x"302114",x"302114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"180f07",x"1c1208",x"211409",x"1f1309",x"261709",x"231509",x"201309",x"201308",x"211409",x"241609",x"241609",x"251509",x"26160a",x"24160a",x"25160a",x"24160a",x"23150a",x"231509",x"24150a",x"23150a",x"231509",x"231509",x"231509",x"24150a",x"231409",x"24150a",x"221409",x"211309",x"221409",x"231509",x"231509",x"221409",x"221409",x"221409",x"231509",x"24150a",x"24150a",x"23150a",x"24150a",x"24150a",x"24150a",x"24150a",x"24160a",x"24150a",x"26160a",x"24150a",x"231409",x"24150a",x"26160a",x"26160a",x"25160a",x"27170a",x"27170a",x"27170a",x"25150a",x"241509",x"231409",x"231409",x"241509",x"241509",x"241409",x"241509",x"231409",x"27160a",x"26160a",x"25150a",x"25150a",x"25150a",x"251509",x"26160a",x"27170a",x"28170a",x"27170a",x"27160a",x"26160a",x"251509",x"25150a",x"241409",x"26160a",x"27170a",x"27160a",x"26160a",x"25150a",x"26160a",x"241509",x"231509",x"221409",x"201309",x"201309",x"211409",x"1f1309",x"1e1208",x"1e1209",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1c1108",x"1c1108",x"1d1208",x"1c1108",x"1c1108",x"1e1208",x"1f1309",x"1e1208",x"1e1208",x"1f1309",x"201309",x"201309",x"211409",x"201409",x"221409",x"201409",x"1e1308",x"1c1108",x"1e1308",x"201409",x"1e1309",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"180f07",x"191008",x"1a1008",x"1c1108",x"1d1108",x"1e1208",x"1f1309",x"1f1309",x"201309",x"201309",x"201309",x"1f1309",x"1e1209",x"1d1208",x"1c1108",x"1b1108",x"191008",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"221608",x"231608",x"221508",x"241608",x"251709",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"392210",x"150e07",x"25160a",x"371f0e",x"3a210f",x"361f0e",x"341e0d",x"351f0e",x"381f0e",x"351d0d",x"321c0d",x"321d0d",x"381f0d",x"331c0b",x"301a0a",x"321c0b",x"301a0a",x"321c0b",x"391f0d",x"3e2310",x"3b220f",x"3e2410",x"361e0d",x"3a210f",x"371f0e",x"3a210f",x"3b210f",x"3e2310",x"402411",x"3b210f",x"3a210f",x"38200e",x"3b220f",x"3d2310",x"3d2310",x"402511",x"422612",x"3e2410",x"3e2310",x"371f0e",x"39200f",x"3a210f",x"381f0e",x"402511",x"3d2310",x"3d230f",x"422712",x"432713",x"452914",x"3e2411",x"3a2210",x"3d2411",x"3c210f",x"3c2210",x"402511",x"402512",x"432712",x"3c220f",x"3a220f",x"3c2310",x"3c2210",x"472914",x"1e1209",x"3d2311",x"3c2311",x"392110",x"2d190b",x"361e0e",x"3a2110",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c311f",x"4c311f",x"513c2f",x"5d4331",x"5e412f",x"5d402c",x"5b3e2a",x"563a28",x"5a3f2d",x"5c402d",x"5b3f2d",x"593c2a",x"5c3d27",x"61412a",x"5f3f2a",x"61412c",x"5a402f",x"5d3f2c",x"62412c",x"664732",x"634431",x"614532",x"5e4332",x"684833",x"634532",x"5e422f",x"654633",x"664836",x"5f4533",x"6c4d39",x"624634",x"5d4535",x"544134",x"574235",x"523f31",x"584233",x"654937",x"614838",x"614735",x"644937",x"5c4435",x"614736",x"5d4435",x"604634",x"5c4434",x"604636",x"644835",x"654836",x"664936",x"634836",x"614534",x"5d4534",x"644733",x"634735",x"684a36",x"644937",x"634836",x"644734",x"664835",x"674934",x"624534",x"644836",x"674a37",x"5f4432",x"5a4231",x"5e4331",x"6a4c37",x"614532",x"5f4432",x"634532",x"5a402e",x"5a4131",x"5a4130",x"553d2d",x"5a402d",x"553b2a",x"4e3626",x"5f3e27",x"5b3c27",x"533827",x"4b3323",x"513625",x"553a26",x"583b27",x"4a3120",x"513625",x"5b3c27",x"65422b",x"5c3c27",x"61402a",x"513828",x"4c3525",x"4f392a",x"5b402f",x"563d2b",x"5a3f2e",x"503b2d",x"543e2f",x"513b2c",x"594030",x"543e2e",x"5a3f2d",x"423125",x"47352a",x"362e26",x"3e3228",x"453529",x"563c2b",x"523520",x"150e07",x"150e07",x"150e07",x"150e07",x"4a2a14",x"191007",x"302113",x"291c10",x"2a1d11",x"2a1e12",x"261a0f",x"2d2014",x"2b1e12",x"2e2014",x"312216",x"302114",x"2f2114",x"2d2013",x"322316",x"2f2114",x"312315",x"342416",x"362718",x"342516",x"342517",x"362719",x"322214",x"332314",x"342416",x"392819",x"332416",x"342416",x"3a291a",x"382719",x"382819",x"362619",x"362619",x"39291b",x"332416",x"332416",x"322316",x"2f2114",x"382819",x"322316",x"362719",x"302215",x"372719",x"3a281a",x"382719",x"2f2114",x"342416",x"382719",x"332416",x"322315",x"392819",x"342516",x"332416",x"362718",x"322315",x"2f2013",x"312214",x"362718",x"39281a",x"342416",x"342517",x"342417",x"362719",x"362619",x"342517",x"37281a",x"302214",x"312215",x"2c1e12",x"2a1e12",x"261a0f",x"302215",x"2d2014",x"302215",x"342517",x"2e2014",x"2e2014",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"160e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"191008",x"1d1208",x"201409",x"211408",x"221409",x"211408",x"25170a",x"241609",x"251609",x"251609",x"26160a",x"25170b",x"24150a",x"23150a",x"24150a",x"221409",x"221409",x"23150a",x"24150a",x"24160a",x"23150a",x"231409",x"25160a",x"24160a",x"25160a",x"25160a",x"26160a",x"26170b",x"26160b",x"221409",x"25160a",x"27170b",x"24160a",x"24150a",x"24150a",x"24150a",x"25160a",x"24150a",x"24160a",x"25160a",x"25160a",x"25160a",x"26170b",x"26170b",x"26170b",x"26170b",x"27170b",x"27170b",x"25160a",x"241509",x"28180b",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"25160a",x"26160a",x"27170a",x"25160a",x"28170b",x"27160a",x"26160a",x"26160a",x"27170a",x"28170b",x"28170b",x"28180b",x"28180b",x"28170b",x"27160a",x"26160a",x"26150a",x"241509",x"29190b",x"27170a",x"251509",x"211308",x"201308",x"201308",x"201208",x"221409",x"231409",x"231409",x"221409",x"221409",x"211409",x"1f1208",x"1f1309",x"1f1209",x"1e1208",x"1e1209",x"1e1208",x"1d1208",x"1d1208",x"1d1208",x"1c1108",x"1d1108",x"1d1108",x"1d1208",x"1d1208",x"1d1108",x"1d1108",x"1d1208",x"1e1208",x"1d1108",x"1e1208",x"1f1309",x"1f1309",x"1f1309",x"201409",x"21140a",x"201309",x"211509",x"201408",x"211408",x"1b1108",x"1b1108",x"1c1208",x"1d1208",x"1e1209",x"181007",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"1a1008",x"1d1209",x"1e1209",x"1f1209",x"1f1209",x"1f1309",x"201309",x"201409",x"1f1309",x"1f1309",x"1f1309",x"1d1208",x"1c1108",x"1b1108",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"261809",x"291a09",x"251708",x"251709",x"271909",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"37200f",x"150e07",x"231409",x"381f0e",x"361f0e",x"38200f",x"221409",x"3c220f",x"452712",x"3f2310",x"3a200d",x"371e0c",x"432510",x"44250f",x"3c210d",x"3c210d",x"42240f",x"43250f",x"3f220e",x"3b200d",x"432712",x"452712",x"402310",x"452813",x"432611",x"482a14",x"482914",x"462712",x"462711",x"442712",x"412511",x"472812",x"462812",x"472812",x"472812",x"462711",x"492913",x"472913",x"502f18",x"482b14",x"442813",x"462812",x"442711",x"452712",x"4a2b14",x"462913",x"4a2b15",x"503017",x"513017",x"4b2c15",x"482a13",x"432611",x"442611",x"3d220f",x"432611",x"482913",x"452712",x"452712",x"472913",x"4a2a14",x"4d2c14",x"150e07",x"26160a",x"351e0d",x"38200f",x"3c2210",x"37200f",x"3b210f",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c321e",x"4c321e",x"513b2d",x"563e2e",x"5e4230",x"593e2d",x"614330",x"5e3f2b",x"5d412f",x"5d3f2c",x"583b2a",x"583825",x"5d3e2b",x"5d3c29",x"563927",x"5f3f2c",x"644530",x"684833",x"664531",x"654531",x"604433",x"5a4131",x"614331",x"684834",x"644733",x"6b4a35",x"664631",x"624634",x"594132",x"563f31",x"644533",x"5e4535",x"5b4637",x"594335",x"5e4637",x"614635",x"644939",x"5b4436",x"684b3a",x"614838",x"664a37",x"654c3b",x"634938",x"624735",x"684d3b",x"614838",x"634837",x"694d3b",x"6b4d3a",x"6b4d39",x"674a38",x"624635",x"654734",x"614534",x"614533",x"634634",x"6a4933",x"6c4a34",x"694833",x"664531",x"664530",x"614331",x"61422e",x"604431",x"584031",x"5d412e",x"5f4635",x"5f4535",x"63442f",x"5f4534",x"5a4333",x"553e2e",x"4e392b",x"4c3526",x"503828",x"4e3828",x"593c29",x"553826",x"563a27",x"563b28",x"4f3524",x"4d3424",x"473122",x"4f3524",x"513623",x"523724",x"4f3422",x"593823",x"5a3a23",x"5c3c26",x"4e3321",x"4b3121",x"5d3d2a",x"60412e",x"573d2c",x"583d2b",x"543d2f",x"533d2e",x"503827",x"4c3729",x"49372b",x"5b412e",x"52392a",x"47362a",x"453428",x"47382d",x"3d332a",x"453529",x"4a301e",x"150e07",x"150e07",x"150e07",x"150e07",x"472914",x"181007",x"2f2011",x"2a1d11",x"302214",x"261a0f",x"2a1d11",x"291d11",x"2e2013",x"2c1e12",x"2e1f13",x"2c1e12",x"2d1f12",x"302114",x"322215",x"2e2013",x"312315",x"322316",x"342516",x"342517",x"312215",x"342415",x"342415",x"2e2012",x"322214",x"312215",x"2f2013",x"2e1f12",x"2f2013",x"312215",x"332416",x"382819",x"352517",x"352617",x"342416",x"352517",x"352517",x"39281a",x"322315",x"382718",x"362618",x"322316",x"362517",x"322315",x"2d1f12",x"372618",x"322315",x"362618",x"332416",x"382719",x"312215",x"2e2013",x"2e2013",x"342415",x"362516",x"2d1f12",x"2e1f12",x"2f2114",x"2f2013",x"2c1e12",x"2b1d11",x"2d1f12",x"332416",x"322416",x"342416",x"352517",x"2c1e12",x"322416",x"332416",x"2b1e12",x"281c10",x"2d2013",x"2a1d11",x"2a1d11",x"2a1d11",x"2b1e12",x"2b1e12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"201409",x"231509",x"211508",x"24150a",x"221509",x"231509",x"261709",x"25160a",x"24150a",x"24160a",x"23150a",x"231509",x"221409",x"211409",x"211409",x"211409",x"221409",x"221409",x"221409",x"231509",x"25160a",x"241509",x"25160a",x"24150a",x"241509",x"26170a",x"25160a",x"27170b",x"28180b",x"24150a",x"24150a",x"25160a",x"25160a",x"25160a",x"24160a",x"25160a",x"25160a",x"24150a",x"24150a",x"231509",x"221409",x"24150a",x"25160a",x"25150a",x"24150a",x"24150a",x"25150a",x"25160a",x"25150a",x"25160a",x"25160a",x"26160a",x"26160a",x"26160a",x"25160a",x"25150a",x"25150a",x"26160a",x"25150a",x"241509",x"241509",x"27170a",x"28180b",x"27170a",x"27170a",x"27160a",x"26160a",x"27160a",x"28180b",x"28170b",x"28170a",x"28170a",x"29180b",x"241509",x"231409",x"251509",x"261609",x"241509",x"221409",x"221409",x"241409",x"241409",x"1f1208",x"221409",x"211309",x"201309",x"201309",x"201409",x"1f1209",x"201309",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1e1309",x"1d1209",x"1d1208",x"1d1208",x"1d1208",x"1d1208",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"201309",x"201408",x"1e1208",x"221509",x"1d1108",x"1a1008",x"1b1008",x"1b1108",x"1b1107",x"1a1007",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"191008",x"1b1108",x"1d1108",x"1d1108",x"1e1209",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1d1208",x"1c1108",x"1a1008",x"191008",x"180f08",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1f1408",x"1d1308",x"211508",x"231608",x"251708",x"271909",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1e1208",x"361f0f",x"150e07",x"1e1208",x"311b0c",x"371f0e",x"3b2311",x"482a14",x"28170a",x"2b180b",x"2b180a",x"2f1a0b",x"281609",x"251509",x"2b180a",x"2a180a",x"28170a",x"2a170a",x"241409",x"27160a",x"271609",x"29170a",x"2a190b",x"27170a",x"2b190c",x"2a180b",x"2b180b",x"28170a",x"2a180b",x"28170a",x"2c190b",x"28170a",x"27170a",x"2f1c0d",x"2e1b0c",x"2e1a0c",x"29170a",x"2c190b",x"2b180b",x"2b180b",x"251509",x"28170a",x"2c190b",x"2f1b0c",x"2d1a0b",x"2e1a0b",x"2a180b",x"29180b",x"29180b",x"2b190b",x"29180a",x"29170a",x"26160a",x"251509",x"27160a",x"241409",x"271509",x"28160a",x"2b180a",x"28160a",x"311c0c",x"341d0d",x"2b180b",x"1c1108",x"2d190b",x"2f1a0b",x"301b0c",x"331d0d",x"3c210f",x"301b0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482e1c",x"482e1c",x"58402e",x"59402f",x"644632",x"654733",x"61432e",x"5c3e29",x"60402b",x"593c2b",x"573928",x"553825",x"5c3a26",x"5b3b27",x"573a29",x"543825",x"5e402c",x"5e412f",x"5c3e2d",x"5a3e2c",x"5a3e2d",x"533a2b",x"603f2b",x"66452f",x"6c4b34",x"684934",x"5c4232",x"5f4230",x"5d4231",x"5c4231",x"543e30",x"563f30",x"5b4334",x"594233",x"5e4331",x"594030",x"5a402e",x"624532",x"543d2e",x"644734",x"614533",x"654936",x"604533",x"5c4231",x"644532",x"5d4230",x"5d3f2d",x"61412d",x"6a4731",x"624431",x"614431",x"654834",x"664735",x"644735",x"644837",x"634837",x"5d4434",x"5f4535",x"604637",x"624737",x"684b38",x"5f4534",x"5c4434",x"584334",x"5d4636",x"5e4636",x"5d4638",x"533e30",x"553f30",x"543e2f",x"4d3a2d",x"503d2f",x"4d392b",x"443227",x"4e382b",x"473327",x"493427",x"4d3423",x"422e21",x"453023",x"513524",x"4d3121",x"442f20",x"422f22",x"4f3524",x"4e3423",x"4e3626",x"5f4029",x"5c3c25",x"583b27",x"503323",x"523625",x"493121",x"533a2b",x"513929",x"593c2a",x"543c2d",x"513b2d",x"48372a",x"49382c",x"392d24",x"573c2c",x"4a3527",x"47372c",x"4a392d",x"4c3a2c",x"45372d",x"423327",x"452c1c",x"150e07",x"150e07",x"150e07",x"150e07",x"4b2c15",x"150e07",x"25190e",x"271b10",x"271b10",x"2c1e12",x"2a1d11",x"2e2014",x"291d11",x"2d1f13",x"302114",x"2f2114",x"2a1d11",x"2d1f12",x"2c1e12",x"332416",x"322315",x"2e2013",x"2e2013",x"312215",x"322315",x"2e1f12",x"2a1c10",x"2f2013",x"322314",x"302214",x"332314",x"2e2013",x"312215",x"322315",x"312215",x"3b2a1a",x"342416",x"322315",x"352517",x"352517",x"312215",x"322315",x"362517",x"372718",x"2d1f13",x"352517",x"362618",x"322316",x"2b1e12",x"2f2013",x"332415",x"362517",x"362517",x"312214",x"342415",x"312215",x"302114",x"2e1f12",x"2f2013",x"312214",x"362617",x"342416",x"2f2013",x"302114",x"312215",x"322315",x"322316",x"2f2114",x"2a1d11",x"2c1f12",x"2d1f13",x"291c11",x"312215",x"2e2013",x"2e1f13",x"2e2114",x"271b10",x"2b1e12",x"271b10",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"1f1308",x"221509",x"211408",x"231509",x"201309",x"221509",x"25160a",x"201309",x"211409",x"201309",x"201309",x"201208",x"201208",x"1f1208",x"1e1208",x"1c1108",x"1e1208",x"1f1208",x"201309",x"211309",x"221409",x"221409",x"231409",x"231409",x"241509",x"241509",x"25160a",x"27170b",x"27170b",x"27170b",x"27170b",x"24150a",x"211309",x"211309",x"221409",x"24150a",x"24160a",x"25160a",x"24150a",x"25160a",x"24150a",x"231509",x"231509",x"241509",x"231509",x"231509",x"25160a",x"25160a",x"25160a",x"25160a",x"26160a",x"25160a",x"241509",x"231409",x"211309",x"221309",x"241509",x"25150a",x"25150a",x"231409",x"231409",x"241409",x"251509",x"241509",x"241509",x"241509",x"26160a",x"28170b",x"2a190b",x"28170b",x"241509",x"261609",x"221308",x"261609",x"211308",x"231409",x"251509",x"251509",x"241509",x"211309",x"201208",x"231409",x"1e1208",x"211309",x"211409",x"221409",x"211409",x"1f1209",x"1e1209",x"1e1208",x"1d1108",x"1d1108",x"1d1208",x"1d1208",x"1d1108",x"1d1208",x"1c1108",x"1b1108",x"1b1008",x"1a1008",x"1b1108",x"1b1108",x"1b1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1e1208",x"1d1208",x"201409",x"1e1208",x"1f1309",x"201409",x"1c1108",x"180f07",x"170f07",x"1a1107",x"1a1107",x"171007",x"170e07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"180f07",x"1a1108",x"1c1108",x"1d1208",x"1e1209",x"1e1209",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1d1209",x"1c1108",x"1b1108",x"1a1008",x"180f08",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1308",x"191007",x"251809",x"2d1c09",x"231608",x"241709",x"241708",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1e1208",x"392110",x"150e07",x"201309",x"311c0d",x"321c0d",x"301b0c",x"2d1a0b",x"341d0d",x"351e0c",x"391f0d",x"311b0b",x"361d0c",x"3b210e",x"371f0d",x"391f0d",x"391f0d",x"3c210e",x"3c210e",x"311a0a",x"391f0d",x"321c0b",x"402511",x"432712",x"3a2110",x"3f2410",x"3f2410",x"38200e",x"3c220f",x"3b210f",x"3a200e",x"3e2310",x"402511",x"3f2410",x"422611",x"422511",x"402511",x"3f2511",x"442813",x"3e2310",x"3e2310",x"422511",x"432713",x"402511",x"3e2411",x"422612",x"3e2411",x"3e2411",x"402511",x"3a200f",x"3c210f",x"351d0c",x"361d0d",x"351d0d",x"3b200e",x"351d0c",x"3b210e",x"412511",x"39210f",x"3e2310",x"3d2310",x"3c220f",x"3c210e",x"150e07",x"2d190b",x"2a170a",x"2e1a0b",x"27160a",x"3d220f",x"311c0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d311e",x"4d311e",x"5f4737",x"583f2d",x"573c2c",x"614533",x"5c3f2d",x"634532",x"62422b",x"5e3e2a",x"61422d",x"60402a",x"593d2b",x"593c2a",x"523725",x"593b29",x"65432d",x"674734",x"61432f",x"5d4230",x"5d4230",x"5b4130",x"583e2d",x"5f4330",x"60432f",x"5a4130",x"5b402e",x"5b402e",x"5d4332",x"543f31",x"624432",x"614635",x"564032",x"574335",x"5b4535",x"5f4536",x"5a4537",x"684c3a",x"60493a",x"624837",x"654c3b",x"674b38",x"684c3a",x"6a4e3c",x"674b39",x"6b503e",x"634a3a",x"644938",x"654a38",x"684d3b",x"654a38",x"614737",x"664b39",x"654b3a",x"644938",x"644936",x"614634",x"654b39",x"674936",x"674936",x"634736",x"614634",x"614735",x"5c4332",x"5b4233",x"533f30",x"584131",x"5a4436",x"534033",x"503f33",x"4f3e32",x"4f3d31",x"4a3528",x"4f3a2d",x"5c3f2d",x"523827",x"4f3625",x"503727",x"433225",x"423022",x"422e22",x"453023",x"402e22",x"3c2b20",x"402c1f",x"462f20",x"382a1f",x"4d3222",x"4f3323",x"493121",x"613e25",x"583924",x"452f21",x"5c3d27",x"5f3f2a",x"5c3e2c",x"483123",x"47372c",x"3d2e23",x"413025",x"47382d",x"45362c",x"453327",x"302720",x"473427",x"463326",x"433328",x"4b3b30",x"4e321e",x"150e07",x"150e07",x"150e07",x"150e07",x"40240f",x"150e07",x"22170d",x"261a0f",x"281c10",x"261a0f",x"2b1e12",x"2c1e12",x"271a0f",x"291d11",x"291d11",x"332416",x"312316",x"2c1e12",x"312215",x"322315",x"372718",x"352517",x"302114",x"362517",x"302114",x"372719",x"362517",x"342517",x"362617",x"322316",x"322316",x"362617",x"392819",x"342516",x"342416",x"352517",x"342417",x"312214",x"2f2013",x"2e2013",x"312214",x"332415",x"312214",x"352517",x"302114",x"352516",x"352517",x"332416",x"372719",x"342416",x"362618",x"372718",x"3b2a1a",x"352517",x"342415",x"322315",x"352516",x"372719",x"392818",x"352517",x"342416",x"312215",x"322316",x"312214",x"392819",x"312215",x"2c1e12",x"322315",x"312215",x"291d11",x"291c10",x"2e2013",x"2a1d11",x"281c10",x"261a0f",x"2e2013",x"281c10",x"2d1f13",x"2b1e12",x"2c1e12",x"2c1e12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1b1108",x"201408",x"231509",x"26170a",x"211409",x"241609",x"27170a",x"201309",x"1f1309",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1d1108",x"1f1209",x"201309",x"201309",x"211409",x"221409",x"211309",x"201208",x"221409",x"211309",x"231509",x"221409",x"211308",x"221409",x"231409",x"231509",x"231409",x"23150a",x"231509",x"23150a",x"24150a",x"24150a",x"231509",x"211309",x"211309",x"221409",x"221409",x"211409",x"221409",x"221409",x"231409",x"231509",x"221409",x"211409",x"231509",x"221409",x"231509",x"24150a",x"23150a",x"231509",x"24150a",x"221409",x"231509",x"231409",x"231409",x"24150a",x"26160a",x"25160a",x"25160a",x"27170b",x"26160a",x"25160a",x"27170a",x"26160a",x"231409",x"26160a",x"211308",x"261509",x"211308",x"261609",x"251509",x"231409",x"231409",x"241409",x"241509",x"211308",x"211308",x"201308",x"211309",x"211409",x"22140a",x"201309",x"1f1209",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1b1108",x"1b1108",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1108",x"1a1008",x"1b1008",x"1d1208",x"1c1108",x"221508",x"1b1107",x"211508",x"1d1208",x"181007",x"170f07",x"181007",x"181007",x"191007",x"171007",x"170e07",x"160f07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"190f07",x"1a1008",x"1b1108",x"1c1108",x"1d1208",x"1d1208",x"1d1208",x"1d1209",x"1c1108",x"1b1108",x"191008",x"180f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1408",x"221508",x"2b1b09",x"281909",x"241709",x"261809",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1f1309",x"37210f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"321d0d",x"381f0d",x"331c0b",x"311b0b",x"361e0c",x"341d0c",x"311b0b",x"301a0a",x"2e190a",x"331c0b",x"341d0c",x"321c0b",x"2f190a",x"371e0d",x"321b0b",x"341d0d",x"361e0d",x"331d0d",x"321b0c",x"321b0c",x"29170a",x"2f1a0b",x"311b0c",x"311b0c",x"301b0b",x"381f0d",x"381f0e",x"3b210f",x"391f0d",x"3c220f",x"3c220f",x"3a200f",x"3a210f",x"3c2210",x"3b2210",x"3d2310",x"381f0e",x"341d0d",x"321c0c",x"39210f",x"3d2310",x"39200f",x"3a200f",x"371f0e",x"3e220f",x"3b200e",x"381f0e",x"39200f",x"39200e",x"351e0e",x"3f2411",x"361e0d",x"3a220f",x"402512",x"3f2410",x"482913",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"381f0d",x"321c0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50331f",x"50331f",x"563f31",x"5a4131",x"5c4130",x"614532",x"614532",x"644633",x"624532",x"5e402c",x"5b3c2a",x"5c3d28",x"583c29",x"573b28",x"563a28",x"5e3f2b",x"62422c",x"5a3c29",x"5e402e",x"563c2c",x"543c2c",x"563e2e",x"594030",x"5c412f",x"593e2d",x"593f2e",x"553e2f",x"593f2f",x"523e30",x"5a4130",x"553f30",x"4f3b2c",x"4f3c30",x"533c2e",x"583e2e",x"604532",x"5c4536",x"624736",x"604839",x"654a3a",x"62493a",x"614939",x"604533",x"5b4132",x"5c4333",x"604737",x"5d4331",x"5c4333",x"604534",x"5c4333",x"5b4333",x"624735",x"5c4536",x"5e4839",x"644a38",x"644a3a",x"614939",x"664b39",x"694d3b",x"664b3a",x"5e4636",x"5c4536",x"5f4737",x"5f4535",x"584435",x"584131",x"594233",x"523e2f",x"513d2f",x"5a4131",x"553d2d",x"523b2c",x"563d2e",x"553b2a",x"5f412d",x"51392a",x"4c372a",x"543b2a",x"4e3727",x"483121",x"4f3423",x"483325",x"473021",x"473022",x"432d1f",x"4d3120",x"472f21",x"4b301e",x"503422",x"503522",x"5e3c26",x"5f3e27",x"493222",x"503421",x"503524",x"4d3524",x"543928",x"463427",x"483223",x"3d2d22",x"46352a",x"46362a",x"4a3629",x"453529",x"463223",x"48362a",x"4e3b2d",x"483628",x"4c311e",x"150e07",x"150e07",x"150e07",x"150e07",x"3e220e",x"150e07",x"291d11",x"261a10",x"2a1d11",x"2c1f12",x"2a1d11",x"342517",x"2d1f13",x"2c1e12",x"312214",x"302114",x"2e2013",x"322316",x"332416",x"332416",x"352517",x"312215",x"322315",x"372719",x"3a281a",x"312215",x"302114",x"2f2114",x"322214",x"342415",x"382718",x"312214",x"342416",x"392819",x"322316",x"362618",x"3a2b1c",x"38291a",x"362618",x"352517",x"352517",x"342416",x"382819",x"382819",x"352517",x"332416",x"322315",x"352517",x"332416",x"362618",x"342516",x"352517",x"312315",x"342416",x"342416",x"372719",x"362617",x"322416",x"332315",x"352516",x"2f2013",x"2d1e12",x"2d1f13",x"342416",x"332315",x"362618",x"2e2013",x"332416",x"302316",x"342618",x"2b1f13",x"332416",x"2e2014",x"281c10",x"2a1d11",x"2b1e12",x"312315",x"2c1e12",x"2c1e12",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"180f07",x"191008",x"1b1108",x"1d1108",x"1f1208",x"201308",x"211408",x"241609",x"231509",x"1f1309",x"1f1208",x"1f1209",x"1e1208",x"1e1208",x"1d1208",x"1e1208",x"1d1208",x"1d1208",x"1f1209",x"1e1208",x"1f1309",x"221409",x"221409",x"231509",x"24150a",x"24150a",x"231509",x"231409",x"241509",x"241509",x"221409",x"231409",x"25160a",x"25150a",x"24150a",x"24150a",x"24150a",x"24150a",x"231509",x"221409",x"221409",x"221409",x"211409",x"221409",x"221409",x"221409",x"211409",x"221409",x"221409",x"211409",x"221409",x"221409",x"231509",x"231509",x"221409",x"221409",x"211309",x"231509",x"24150a",x"231509",x"211309",x"231509",x"24150a",x"231509",x"221409",x"231409",x"231409",x"25150a",x"25150a",x"25160a",x"26160a",x"27160a",x"231409",x"261609",x"211308",x"261509",x"251509",x"221408",x"201308",x"201208",x"221309",x"241509",x"221409",x"201308",x"201308",x"211309",x"1f1309",x"1f1208",x"1e1208",x"1c1108",x"1b1108",x"1b1008",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1b1008",x"1b1108",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1108",x"1a1008",x"1b1008",x"1d1208",x"1c1208",x"1d1208",x"201409",x"1d1208",x"1f1308",x"1c1107",x"1a1007",x"180f07",x"170f07",x"180f07",x"181007",x"180f07",x"180f07",x"160e07",x"150e07",x"170f07",x"160e07",x"170f07",x"180f07",x"191008",x"1b1108",x"1d1208",x"1d1108",x"1d1209",x"1e1209",x"1d1208",x"1c1108",x"1b1108",x"1a1108",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1308",x"1a1107",x"261809",x"291a09",x"201408",x"211508",x"211508",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1d1208",x"36200f",x"150e07",x"150e07",x"3e220f",x"3a200e",x"3a200e",x"3b210f",x"3a200d",x"3e220e",x"351c0b",x"391f0d",x"3a200d",x"351d0b",x"331c0b",x"341c0b",x"3b200d",x"40230f",x"3d210e",x"3b200d",x"3d210e",x"3c210e",x"371e0d",x"301b0b",x"2e1a0b",x"331c0c",x"301b0b",x"361e0d",x"341d0c",x"391f0d",x"39200e",x"361d0c",x"351c0b",x"351c0c",x"381e0c",x"371c0c",x"391f0d",x"361d0c",x"391e0d",x"381f0d",x"3d220f",x"3d220f",x"3e230f",x"3f2410",x"3d220f",x"412411",x"402411",x"412411",x"422611",x"432611",x"3f230f",x"3d210f",x"422611",x"3f2310",x"3e230f",x"3d220f",x"3e230f",x"3c210f",x"381f0e",x"3b210e",x"3a200e",x"391f0d",x"381e0c",x"361d0c",x"3c210e",x"2a180a",x"1e1208",x"150e07",x"331c0c",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c301d",x"4c301d",x"5d4333",x"563c2b",x"614634",x"5b4232",x"5b4131",x"5e4333",x"573c2c",x"5b3f2d",x"583f2f",x"503524",x"533b2a",x"583e2c",x"573e2e",x"523729",x"523a29",x"573b29",x"5b3f2e",x"563d2e",x"573d2d",x"533b2b",x"543c2d",x"573e2d",x"593e2d",x"5d3f2d",x"543a2a",x"563c2b",x"5b3e2b",x"583d2b",x"523b2c",x"503a2c",x"533d2e",x"564031",x"634735",x"5f4635",x"5c4434",x"674936",x"5b4536",x"644b3b",x"654b3b",x"6b4f3e",x"664d3c",x"664b3a",x"664b3a",x"624a39",x"634c3d",x"664c3c",x"5e4433",x"5d4537",x"574234",x"594538",x"5c473a",x"594436",x"574335",x"5b473a",x"5f493b",x"664a39",x"614939",x"644937",x"644a39",x"624939",x"61493a",x"634937",x"634837",x"5e4637",x"624a3a",x"5a4334",x"594234",x"5c4535",x"594335",x"583f2f",x"543e2f",x"573f31",x"594030",x"533929",x"523a2a",x"4e3626",x"463226",x"433024",x"443024",x"3b2b20",x"463022",x"3f2c1e",x"36271d",x"3e2c1f",x"402c1f",x"402c1f",x"492f1f",x"4c3323",x"553825",x"432d1f",x"452e20",x"412d20",x"3a291e",x"4a301f",x"442f22",x"4b3627",x"513828",x"3b2d23",x"48372b",x"423024",x"3a3027",x"423328",x"45352a",x"453429",x"45352a",x"46372b",x"51331f",x"150e07",x"150e07",x"150e07",x"150e07",x"361d0b",x"150e07",x"2a1d11",x"2e2013",x"2a1d11",x"2b1d12",x"2c1e12",x"342416",x"2d1f12",x"2c1f12",x"2d1f13",x"322315",x"2e1f13",x"2e2013",x"2f2114",x"312215",x"342416",x"352517",x"312215",x"342516",x"342516",x"322315",x"352516",x"332416",x"342416",x"322215",x"372617",x"3a291a",x"3c2a1b",x"3a2a1b",x"3d2b1c",x"3b2a1b",x"392819",x"372719",x"392819",x"3a2819",x"322315",x"342516",x"322215",x"382718",x"3a2919",x"322316",x"352517",x"362517",x"302114",x"382718",x"3a291a",x"332416",x"342416",x"382719",x"2f2114",x"362617",x"3a291a",x"3a2818",x"372718",x"332416",x"322315",x"322215",x"342416",x"322316",x"332416",x"342517",x"312215",x"322416",x"352517",x"332517",x"332416",x"2e2013",x"281c10",x"2b1d11",x"2a1d11",x"2e2013",x"2b1d11",x"2a1d11",x"2c1e12",x"2c1e12",x"2c1e12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"201409",x"231509",x"201408",x"201408",x"251609",x"24150a",x"201409",x"1f1309",x"1e1208",x"1d1108",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1108",x"1e1208",x"1f1208",x"211309",x"221409",x"221409",x"221409",x"221409",x"221409",x"211309",x"241509",x"231509",x"221409",x"201309",x"201308",x"1f1208",x"201208",x"201309",x"1f1208",x"201309",x"1f1308",x"201308",x"1f1208",x"201208",x"211409",x"1f1208",x"211309",x"201309",x"221409",x"211409",x"201309",x"211309",x"201309",x"211309",x"211409",x"221409",x"211409",x"221409",x"221409",x"1f1208",x"201309",x"211309",x"231409",x"231409",x"241509",x"231409",x"231409",x"241509",x"251509",x"241509",x"211308",x"261509",x"221308",x"261609",x"241509",x"211308",x"201308",x"201308",x"231409",x"241509",x"201308",x"231409",x"1e1208",x"201309",x"201309",x"201309",x"1e1208",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"190f07",x"190f07",x"191008",x"190f07",x"190f07",x"190f07",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1a0f08",x"1e1309",x"201409",x"201408",x"1c1107",x"191007",x"1a1007",x"181007",x"170f07",x"180f07",x"170f07",x"180f07",x"150e07",x"170f07",x"160f07",x"160e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"190f08",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"201408",x"1d1208",x"2a1a09",x"2c1c09",x"211508",x"221608",x"231609"),
(x"150e07",x"150e07",x"150e07",x"1b1008",x"341e0e",x"150e07",x"1e1108",x"2c180a",x"150e07",x"3f230f",x"331b0c",x"3b200d",x"3d210e",x"371e0c",x"3a200d",x"3b200e",x"3b200d",x"371e0c",x"381f0d",x"3e220e",x"3d220e",x"301a0a",x"3b210e",x"341c0b",x"391f0e",x"3c220f",x"361d0d",x"381f0d",x"2f1a0b",x"30190b",x"2c170a",x"361d0c",x"371e0d",x"3a200e",x"3b210e",x"371e0d",x"39200e",x"3c210f",x"3e220f",x"3e230f",x"412410",x"3c210f",x"3c210f",x"3b200f",x"391f0e",x"3a200e",x"3a200e",x"391f0d",x"361e0d",x"381e0d",x"361e0d",x"391f0d",x"331c0c",x"381f0d",x"391f0d",x"381e0d",x"391f0d",x"321b0b",x"311a0b",x"3d220f",x"3d2310",x"402410",x"3f2410",x"3c210f",x"3d210e",x"381f0d",x"2c180b",x"331c0c",x"150e07",x"2f1a0b",x"150e07",x"371e0d",x"341e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452c1a",x"452c1a",x"553f31",x"5d4435",x"554133",x"573f2f",x"5c4435",x"5a4335",x"563f31",x"543b2c",x"4e3728",x"4f3728",x"513a2b",x"523b2c",x"4a3223",x"4c3527",x"4b3427",x"513829",x"513a2b",x"513c2e",x"4b382d",x"4e3a2d",x"4c382c",x"503829",x"553c2c",x"583c2a",x"543a2a",x"593e2d",x"523827",x"5b402f",x"563c2c",x"5b4130",x"563f30",x"614635",x"654735",x"5e4332",x"654837",x"5d4434",x"684935",x"5f4535",x"5c4334",x"614736",x"614939",x"594133",x"5d473a",x"5e4638",x"604737",x"5e4432",x"5f4534",x"624838",x"654a39",x"5b4233",x"614736",x"614736",x"604737",x"644a39",x"5f4636",x"61493a",x"604736",x"5e4535",x"614837",x"614a3b",x"614737",x"624a3b",x"624a3b",x"5a4131",x"5c4537",x"5b4333",x"5b4434",x"5c4538",x"5a4436",x"574235",x"503c2f",x"564134",x"594031",x"60432f",x"5a3e2c",x"563b29",x"4d3526",x"4b3425",x"462f21",x"422d20",x"422c1f",x"412d21",x"422f23",x"36291f",x"422f22",x"412d20",x"452e1f",x"513524",x"462e1d",x"442d1f",x"49301f",x"3a281d",x"513523",x"442e21",x"3e2d21",x"473326",x"473225",x"46362b",x"423328",x"3f3227",x"4a382b",x"3c2e24",x"443429",x"413329",x"3f3127",x"433429",x"50321f",x"150e07",x"150e07",x"150e07",x"150e07",x"40230f",x"150e07",x"24190e",x"2c1f13",x"2b1e12",x"2d2013",x"2e2014",x"2d2013",x"302114",x"2e2013",x"322316",x"322315",x"2d1f13",x"342416",x"322315",x"2e2013",x"302114",x"322315",x"342516",x"352516",x"312215",x"332416",x"342416",x"352617",x"342516",x"312215",x"322315",x"2c1c10",x"352516",x"312214",x"382718",x"39291a",x"3d2c1c",x"382819",x"322214",x"392919",x"322315",x"3a2819",x"362718",x"3c2b1b",x"3b2a1a",x"382718",x"362618",x"3b291a",x"352517",x"342416",x"322315",x"322315",x"372718",x"322315",x"382818",x"352516",x"392819",x"332416",x"322315",x"342416",x"322316",x"2f2114",x"322315",x"281a0e",x"302214",x"2e2013",x"342416",x"352618",x"312216",x"302214",x"2d1f12",x"302215",x"2f2114",x"2f2114",x"2c1f13",x"2b1e12",x"2c1e12",x"281c10",x"2a1d11",x"2d1f13",x"2d1f13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"191008",x"1f1408",x"1f1308",x"251709",x"211409",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1008",x"1b1008",x"1c1108",x"1e1208",x"1e1208",x"1f1309",x"201309",x"201208",x"201309",x"211309",x"201309",x"201308",x"211309",x"231409",x"231409",x"231509",x"231409",x"231409",x"231409",x"211309",x"211309",x"211309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1e1108",x"1d1108",x"1e1108",x"1e1208",x"1e1208",x"1f1208",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"211309",x"221409",x"221409",x"1f1208",x"1f1208",x"1f1208",x"201208",x"201208",x"201208",x"201208",x"211309",x"251509",x"231409",x"231409",x"211308",x"261609",x"211308",x"261509",x"261509",x"241509",x"231409",x"241509",x"251509",x"221409",x"211308",x"221409",x"221409",x"221409",x"1d1108",x"1e1208",x"1d1108",x"1c1108",x"1b1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1008",x"1b1108",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"190f08",x"1a1008",x"191008",x"191008",x"191008",x"191008",x"190f07",x"190f07",x"180f07",x"180f07",x"1c1107",x"1c1107",x"1b1107",x"211508",x"1b1107",x"1c1107",x"191007",x"170f07",x"191007",x"180f07",x"160e07",x"191007",x"160e07",x"160e07",x"160f07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1008",x"1a1008",x"190f07",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"1c1208",x"301e0a",x"1f1408",x"211508",x"251809",x"1d1308"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"38210f",x"150e07",x"150e07",x"191008",x"150e07",x"150e07",x"1a1008",x"150e07",x"1b1008",x"1c1108",x"1a1008",x"180f07",x"1c1108",x"150e07",x"150e07",x"191007",x"170f07",x"150e07",x"150e07",x"1b1108",x"180f07",x"1a1008",x"170f07",x"150e07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"1e1208",x"150e07",x"221409",x"1a1008",x"150e07",x"1f1309",x"1a1008",x"1c1108",x"1c1108",x"180f08",x"190f08",x"150e07",x"180f07",x"180f07",x"170f07",x"170f07",x"150e07",x"1a1008",x"1a1008",x"170f07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"1b1008",x"180f07",x"150e07",x"190f07",x"1f1208",x"231409",x"150e07",x"351c0c",x"341d0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f311d",x"4f311d",x"594537",x"584234",x"604737",x"584030",x"5f4737",x"604534",x"5a402f",x"523a2a",x"442f22",x"453225",x"4e372a",x"4d3728",x"50392a",x"543929",x"4b372b",x"513a2b",x"4f3a2c",x"533e31",x"4f3a2d",x"4e392b",x"533e30",x"543d2f",x"593e2d",x"543b2a",x"533b2d",x"5c3f2d",x"543b2c",x"523d2f",x"553b2a",x"5a3e2c",x"584031",x"573f2d",x"533c2d",x"674835",x"5b4332",x"604737",x"604737",x"5f4636",x"664a38",x"5f4738",x"5e493c",x"5c483b",x"584639",x"5a483b",x"584232",x"5e4637",x"5f4737",x"654b3a",x"674b3a",x"644c3c",x"654b3a",x"634c3d",x"5b4536",x"5e4637",x"634a39",x"5a4334",x"5f4637",x"644937",x"604534",x"5e4332",x"604432",x"634735",x"5b4232",x"5f4331",x"5f4534",x"644a38",x"614635",x"5f4432",x"5e4535",x"5f4635",x"5b4435",x"574132",x"503d30",x"563d2c",x"50392b",x"4b3629",x"50382a",x"513829",x"493224",x"4a3326",x"3f2c21",x"3a2b21",x"31251d",x"39291f",x"372a20",x"4a3120",x"402c1f",x"48301f",x"563826",x"513626",x"442f21",x"3e2d22",x"483224",x"4a3324",x"493021",x"442f23",x"473124",x"48382d",x"413328",x"443227",x"513b2c",x"433022",x"4c382a",x"4b382c",x"473529",x"46362b",x"4f321e",x"150e07",x"150e07",x"150e07",x"150e07",x"3e220e",x"150e07",x"281b10",x"2a1d11",x"261a0f",x"291c11",x"2a1d11",x"302114",x"312315",x"312215",x"312215",x"2d1f12",x"2f2114",x"342416",x"332416",x"302114",x"2f2114",x"352618",x"2d1f13",x"3a291a",x"362719",x"3b2a1b",x"362618",x"352618",x"352517",x"3d2b1c",x"3b2a1b",x"3f2d1d",x"382719",x"382819",x"3f2d1d",x"382819",x"39281a",x"3a2819",x"332316",x"362516",x"352516",x"332315",x"3a2819",x"3b2a1b",x"3e2c1c",x"392819",x"3a2919",x"342416",x"382718",x"382718",x"372718",x"352516",x"342415",x"3c2b1c",x"39281a",x"382819",x"39291a",x"3c2b1c",x"3a291a",x"3b2a1a",x"352517",x"322316",x"38281a",x"362618",x"342416",x"382819",x"372819",x"342517",x"312315",x"312215",x"302114",x"2e2013",x"2b1d11",x"302114",x"302114",x"302114",x"2b1e12",x"291c11",x"2b1d11",x"2d1f12",x"2d1f12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1f1309",x"211409",x"211408",x"251609",x"201308",x"201308",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1d1108",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201208",x"201208",x"201208",x"201208",x"211309",x"24150a",x"24150a",x"24150a",x"231409",x"201308",x"1f1208",x"201309",x"201208",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"1f1208",x"201308",x"201309",x"211409",x"211309",x"201309",x"201208",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1108",x"1e1108",x"1f1208",x"201208",x"201309",x"1f1208",x"1f1208",x"201309",x"211309",x"211309",x"211309",x"211308",x"231409",x"231409",x"231409",x"231409",x"231409",x"251509",x"241509",x"211308",x"251509",x"251509",x"251509",x"241409",x"201208",x"231409",x"221409",x"221409",x"221409",x"201309",x"201309",x"1e1208",x"1d1108",x"1b1008",x"1b1008",x"1b1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"1a1008",x"1b1008",x"1a1008",x"1b1108",x"1f1309",x"1d1208",x"1c1107",x"1b1107",x"1a1007",x"181007",x"160f07",x"170f07",x"180f07",x"170f07",x"160e07",x"170f07",x"160e07",x"150e07",x"160e07",x"160e07",x"160e07",x"180f07",x"191008",x"1b1108",x"1b1108",x"1b1008",x"1a1008",x"1b1008",x"1a1008",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1308",x"211508",x"231608",x"1c1208",x"211508",x"211508"),
(x"150e07",x"150e07",x"150e07",x"180f07",x"281509",x"2f1b0b",x"341d0c",x"351d0d",x"341d0d",x"3c210f",x"3c220f",x"381f0e",x"3a1f0d",x"351d0b",x"3a200d",x"381f0d",x"361e0c",x"381f0d",x"3a200d",x"3a200d",x"361e0c",x"381f0d",x"2e180b",x"311b0c",x"341c0c",x"381f0d",x"361d0c",x"361e0d",x"3a200e",x"361e0d",x"361e0d",x"311b0b",x"301a0b",x"351d0d",x"341d0d",x"361e0d",x"381f0e",x"3c220f",x"3c220f",x"3f2410",x"3b220f",x"3d2310",x"3b210f",x"3d2310",x"39200f",x"371f0e",x"371f0e",x"331c0c",x"331c0d",x"38200e",x"39200e",x"38200f",x"3d2310",x"371f0e",x"31190b",x"331b0c",x"371d0c",x"331c0c",x"3b200e",x"381f0d",x"341d0c",x"371e0d",x"3a200e",x"3a200e",x"361d0c",x"391f0e",x"3a200e",x"3a200e",x"3b210f",x"371f0e",x"371f0e",x"361e0d",x"301b0b",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2e1b",x"4b2e1b",x"544235",x"5b4638",x"543e2f",x"513b2d",x"574336",x"513b2d",x"554033",x"563a2a",x"553928",x"4f382a",x"4e382a",x"51382a",x"563d2d",x"52392a",x"4d382c",x"49372c",x"48362b",x"4f3a2c",x"543c2d",x"50392b",x"563d2d",x"553d2d",x"583d2d",x"5c3f2e",x"593f2e",x"4e392b",x"573d2c",x"583d2c",x"543c2d",x"513c2e",x"513c2d",x"5a4334",x"553f30",x"543e31",x"604635",x"5c4435",x"684b3a",x"604535",x"5c4536",x"5b4435",x"5c483a",x"5b4435",x"5a473a",x"554338",x"574538",x"5b4234",x"5b4638",x"594537",x"614838",x"634a39",x"5b4232",x"644a39",x"634a39",x"604839",x"644a38",x"604736",x"654d3c",x"634938",x"614737",x"644b3b",x"624a3b",x"6a4f3d",x"604535",x"604737",x"5f4838",x"5c4434",x"5d4333",x"5a4336",x"563c2b",x"5b4335",x"574032",x"553f30",x"4f3c2e",x"543d2f",x"543d2e",x"4e3626",x"4b3629",x"533928",x"4c3526",x"493325",x"402e22",x"3f2e23",x"3c2d22",x"3c2d22",x"3f2e22",x"473022",x"452d1e",x"3e2b1e",x"442e20",x"482f20",x"4c3323",x"4f3626",x"503422",x"4b3528",x"503524",x"433126",x"413126",x"422d20",x"443225",x"433327",x"4e3729",x"47362a",x"48392e",x"4d3a2e",x"493a2f",x"4d3c30",x"50311c",x"150e07",x"150e07",x"150e07",x"150e07",x"42240f",x"150e07",x"291c11",x"2c1e12",x"271b0f",x"271b10",x"2d1f13",x"2a1d11",x"302114",x"2c1e12",x"2f2113",x"312214",x"2d1f12",x"2f2013",x"342416",x"2c1e12",x"312214",x"352517",x"312214",x"382718",x"3a281a",x"362618",x"322316",x"322416",x"352517",x"342416",x"362617",x"322316",x"332315",x"342417",x"382718",x"332316",x"3c2a1a",x"3a2819",x"372718",x"3b291a",x"372618",x"332316",x"372718",x"332415",x"352517",x"332416",x"342416",x"352516",x"362517",x"342415",x"362517",x"372617",x"322315",x"382718",x"362617",x"382718",x"3a281a",x"3d2b1c",x"362618",x"342517",x"312315",x"342416",x"312214",x"382718",x"302114",x"2f2014",x"352517",x"322215",x"342517",x"312215",x"2b1e11",x"342416",x"312215",x"2c1e12",x"2c1e12",x"2c1e12",x"2e2013",x"2a1d11",x"2b1e11",x"291c10",x"291c10",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1f1208",x"211409",x"1f1308",x"1f1308",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1f1208",x"1f1208",x"201309",x"221409",x"221409",x"221409",x"231409",x"231409",x"231409",x"231409",x"231409",x"221409",x"231409",x"221409",x"211409",x"201308",x"201309",x"201309",x"1f1308",x"1e1208",x"1e1208",x"1e1208",x"1f1208",x"201308",x"201309",x"201308",x"201308",x"1f1208",x"201308",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"201309",x"201309",x"211309",x"211309",x"201208",x"1f1208",x"1e1108",x"1e1108",x"211409",x"231409",x"221409",x"231409",x"231409",x"201208",x"26160a",x"261609",x"211308",x"251509",x"261609",x"241409",x"231409",x"231409",x"251509",x"241509",x"1f1208",x"231409",x"201308",x"221409",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"180f07",x"1b1107",x"190f07",x"1c1107",x"201408",x"1c1107",x"180f07",x"180f07",x"170f07",x"170f07",x"160e07",x"170e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1f1408",x"1c1208",x"201508",x"201508",x"201408"),
(x"150e07",x"150e07",x"150e07",x"180f07",x"211309",x"2a170a",x"311c0c",x"361e0d",x"38200e",x"371f0e",x"351c0c",x"371f0e",x"39200f",x"391f0d",x"351d0c",x"2f1a0a",x"2c180a",x"2e190a",x"2c180a",x"331c0c",x"311b0c",x"311c0c",x"301a0b",x"331c0c",x"331c0c",x"361f0d",x"351d0d",x"341c0c",x"2d190b",x"341c0c",x"311b0b",x"341c0c",x"371f0e",x"371f0e",x"3a210f",x"371f0e",x"3a210f",x"3d2310",x"39200e",x"39200e",x"361e0d",x"351d0d",x"351d0d",x"331c0c",x"351d0d",x"2f1a0b",x"321c0c",x"2e190b",x"301b0c",x"2e1a0b",x"371f0e",x"361e0d",x"2d190b",x"331d0c",x"371f0e",x"351d0d",x"361e0d",x"341d0c",x"321c0c",x"331c0c",x"341d0c",x"331c0c",x"351d0c",x"361e0d",x"361e0d",x"301b0b",x"331c0c",x"371f0e",x"351e0d",x"351e0d",x"381f0e",x"351e0d",x"301b0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482d19",x"482d19",x"563e2f",x"49372a",x"554134",x"5a4638",x"534032",x"554031",x"544033",x"533d2f",x"543d2f",x"4c3729",x"523b2c",x"4e3a2d",x"4c3629",x"4a372b",x"433127",x"463429",x"513c2f",x"543c2d",x"553f30",x"563d2e",x"543d2d",x"573e2d",x"513a2a",x"4a372b",x"563e2e",x"553f31",x"543c2d",x"4e3b2e",x"503e31",x"523d30",x"553f31",x"563f30",x"594333",x"564133",x"604736",x"5c4535",x"5c4537",x"5b4435",x"5a4333",x"523f32",x"503f32",x"4f3e32",x"524236",x"47392f",x"4b3d32",x"534336",x"554236",x"584639",x"5c493b",x"5d493b",x"574437",x"5a4536",x"5b4739",x"5d4738",x"61493a",x"5e483a",x"574436",x"5c473a",x"5c4334",x"5e4536",x"604636",x"5f4636",x"5b4334",x"5f4433",x"573f30",x"533c2e",x"5f4330",x"5a4132",x"5d4231",x"573e2f",x"50392a",x"513d30",x"4f3c2f",x"503b2e",x"523c30",x"4d3a2d",x"4c392b",x"503829",x"483427",x"473427",x"473122",x"443124",x"352920",x"3e2b1f",x"38291d",x"513523",x"483123",x"433023",x"4c3323",x"4f3424",x"503422",x"4f3322",x"483325",x"473124",x"4c3526",x"4f3728",x"503a2c",x"453429",x"4d382b",x"3e3127",x"4b382c",x"46362b",x"473427",x"4c3c30",x"4b3c31",x"4d3c30",x"4b2f1b",x"150e07",x"150e07",x"150e07",x"150e07",x"442510",x"150e07",x"281c10",x"291c11",x"2c1e12",x"2d1f13",x"2b1d11",x"2d1f12",x"2d1f12",x"291c11",x"322315",x"2f2113",x"2a1c11",x"322215",x"332315",x"2f2013",x"2f2013",x"332416",x"362517",x"362618",x"3c2a1b",x"3a291a",x"382819",x"382718",x"322316",x"352617",x"382819",x"322316",x"382718",x"342416",x"302214",x"302114",x"362617",x"352416",x"3a291a",x"3a291a",x"372718",x"3c2a1b",x"362517",x"382718",x"342415",x"312114",x"352517",x"362617",x"312214",x"2f2013",x"302214",x"302114",x"362517",x"332416",x"352517",x"392819",x"3d2b1c",x"3e2c1d",x"3a291a",x"322315",x"342516",x"342416",x"312215",x"2e2013",x"2d1f13",x"312214",x"2f2113",x"2d1f13",x"302114",x"2f2013",x"2e2013",x"312215",x"302114",x"2d1f13",x"2d1f12",x"291c11",x"281b0f",x"261a0f",x"291c11",x"2a1d11",x"2a1d11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"1c1108",x"1c1108",x"1f1308",x"241609",x"221409",x"1f1308",x"1d1208",x"1e1209",x"1e1209",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1f1208",x"201208",x"201208",x"211409",x"221408",x"221409",x"231509",x"24150a",x"241509",x"231509",x"231409",x"211409",x"201309",x"1f1208",x"201208",x"201309",x"201309",x"201309",x"211309",x"211309",x"211309",x"211309",x"211409",x"1f1308",x"211409",x"1e1208",x"211309",x"201309",x"201309",x"211309",x"1f1209",x"1f1309",x"201309",x"1e1208",x"1f1208",x"1f1208",x"201308",x"1f1208",x"1d1108",x"1a0f07",x"190f07",x"190e07",x"1d1108",x"1f1108",x"201208",x"211308",x"221409",x"231409",x"26160a",x"241509",x"251509",x"211308",x"251509",x"261509",x"251509",x"251509",x"251509",x"211308",x"42260f",x"4a2c11",x"4b2d11",x"4e2e13",x"492b11",x"452810",x"482a11",x"4b2c12",x"4d2d12",x"4a2b13",x"4b2c12",x"4d2d13",x"4f2d14",x"4c2d13",x"452811",x"412510",x"422610",x"41260e",x"3f230f",x"442610",x"3f240f",x"3f240f",x"3f240f",x"3b200d",x"3d220e",x"371e0d",x"361e0d",x"3c210f",x"3e230f",x"3d220f",x"3f230f",x"3e230f",x"402410",x"3d220f",x"3c210e",x"3c210e",x"3c210f",x"3b210e",x"391f0d",x"3c210e",x"3d210f",x"3d220f",x"3b210e",x"3a1f0d",x"3a1f0d",x"3c210e",x"39200e",x"3d220f",x"402410",x"3e2310",x"402410",x"3c220f",x"3e2310",x"422511",x"3e2310",x"3f230f",x"3d210f",x"3e230f",x"3f220f",x"3d210f",x"3f230f",x"402410",x"432611",x"4a2913",x"492913",x"472813",x"472813",x"442611",x"422511",x"402410",x"371e0d",x"170f07",x"371f0e",x"150e07",x"150e07",x"150e07",x"160f07",x"221608",x"201508",x"231609",x"211508",x"221608"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"28160a",x"331c0d",x"341e0d",x"37200f",x"3c2310",x"371f0e",x"311c0c",x"321c0c",x"2b170a",x"351e0e",x"2e1a0c",x"2b190b",x"301b0c",x"311c0c",x"29170a",x"311b0c",x"2d190b",x"2c190b",x"311b0c",x"361f0e",x"361f0e",x"321c0c",x"331c0c",x"2f190b",x"361e0d",x"301c0c",x"301b0c",x"361f0e",x"361f0e",x"361f0d",x"361f0e",x"361e0e",x"351e0e",x"311c0d",x"3b2210",x"361f0e",x"2f1b0c",x"341d0d",x"331d0d",x"351e0e",x"311b0c",x"321c0d",x"321c0d",x"2c190b",x"301b0c",x"361f0e",x"351e0d",x"321c0d",x"351d0d",x"311c0c",x"301a0b",x"311b0b",x"2e190b",x"2a170a",x"2b170a",x"281609",x"29160a",x"2d180a",x"2c180a",x"2d190b",x"301a0b",x"2d190b",x"2e1a0b",x"2f1b0b",x"2e1a0b",x"2b180b",x"2c190b",x"1f1208",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482c18",x"482c18",x"554337",x"564235",x"574437",x"574639",x"59473a",x"5a4436",x"544439",x"514338",x"533e30",x"523e31",x"564132",x"513d2f",x"513929",x"5c4434",x"543b2a",x"533e30",x"574132",x"573d2d",x"554032",x"533e2f",x"584334",x"543f30",x"624735",x"523d2f",x"563f31",x"503c2f",x"573f2f",x"4f3c2f",x"554133",x"584132",x"573f2f",x"594437",x"574131",x"5d4536",x"5f4332",x"584334",x"4e3b2e",x"534133",x"534135",x"4e3f34",x"413529",x"4f3f33",x"4c3c30",x"44392f",x"45372d",x"513d30",x"4f3c2e",x"533d2d",x"4c3b2f",x"543d2f",x"503d30",x"543e2f",x"584233",x"5a4436",x"5b4638",x"5f4738",x"574234",x"584336",x"5b4537",x"5a4538",x"584336",x"614838",x"5d4536",x"614838",x"5d4433",x"5f4839",x"5e4637",x"584233",x"5b4537",x"564235",x"56453a",x"503f32",x"4f3e33",x"503e32",x"503b2e",x"493528",x"4b382b",x"4c382c",x"4a372a",x"3f3229",x"463428",x"4d3627",x"402f24",x"4e3627",x"473326",x"4e3524",x"422f23",x"442f22",x"4c3424",x"543928",x"4d3424",x"4c3628",x"513828",x"4c3628",x"503829",x"513d2f",x"433226",x"4e392b",x"574234",x"46392e",x"4a3b31",x"483a30",x"49382c",x"493b30",x"514236",x"4e4137",x"4b2d1a",x"150e07",x"150e07",x"150e07",x"150e07",x"40230e",x"150e07",x"2d1f12",x"2b1e12",x"332416",x"302215",x"352618",x"2e2013",x"2c1e12",x"2f2114",x"2f2013",x"332315",x"322316",x"2d1f12",x"342416",x"302114",x"362517",x"352516",x"322315",x"362517",x"322316",x"342416",x"3b2a1b",x"3b291a",x"3f2d1d",x"39281a",x"3a291a",x"362517",x"372618",x"362618",x"3a2919",x"362517",x"3a2919",x"3a2919",x"3d2a1a",x"3f2d1c",x"3d2c1c",x"3c2b1c",x"3e2c1d",x"3a2919",x"382819",x"3c2a1b",x"322214",x"362617",x"362618",x"332315",x"342416",x"352517",x"382719",x"312214",x"312214",x"332315",x"342416",x"39281a",x"3b2a1b",x"342416",x"3a291a",x"332416",x"332416",x"2c1f12",x"302114",x"352517",x"332415",x"2f2114",x"372718",x"332416",x"312215",x"352517",x"302215",x"2a1d12",x"312215",x"2c1e12",x"302214",x"2f2114",x"291c10",x"2c1f12",x"2c1f12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"543116",x"462811",x"4a2b12",x"3c220e",x"432710",x"412510",x"3d230f",x"3a210e",x"381f0d",x"331c0c",x"341d0b",x"371e0b",x"351d0c",x"38200c",x"341c0c",x"30190b",x"311b0b",x"331c0b",x"351c0b",x"2d190b",x"331c0c",x"331c0c",x"371e0d",x"341d0d",x"381f0e",x"422510",x"2f1a0b",x"4c2b10",x"43280f",x"42270e",x"462910",x"43280f",x"3f250e",x"41270f",x"422710",x"402610",x"371f0d",x"351e0c",x"331b0b",x"2d180a",x"3b210e",x"3c220e",x"311b0c",x"3b210e",x"331c0b",x"331c0c",x"3e2310",x"361e0d",x"3a210f",x"3a210f",x"3a210f",x"3f2310",x"321c0d",x"361e0d",x"462711",x"42240f",x"3b200d",x"422410",x"472812",x"4a2a13",x"4c2c14",x"442610",x"432510",x"4c2b13",x"4a2a13",x"442610",x"482911",x"4c2c13",x"4e2d14",x"4a2912",x"4c2b12",x"4d2c12",x"502e13",x"553114",x"553113",x"45280c",x"543114",x"533114",x"37220c",x"3c240d",x"3f260e",x"3c240d",x"42270f",x"3e250d",x"40270f",x"3b230c",x"38210c",x"3f250e",x"3c230d",x"3d240e",x"3e250e",x"3b220e",x"3c240f",x"3c240e",x"38200d",x"3b220e",x"371f0e",x"331d0d",x"311d0c",x"311c0b",x"361f0c",x"321c0c",x"311c0c",x"2e1a0b",x"301b0c",x"2f1a0b",x"2d190b",x"2c190b",x"2f1b0c",x"301c0d",x"2b180b",x"2c190b",x"28160a",x"251509",x"29170a",x"281609",x"271509",x"271509",x"231409",x"271509",x"291609",x"28160a",x"28170a",x"2a180a",x"2b180a",x"28170a",x"29170a",x"2e1a0c",x"2d190b",x"311b0c",x"2d190b",x"28160a",x"241509",x"29170a",x"2c190b",x"2d190b",x"2d190b",x"2c190b",x"2e1a0b",x"311c0c",x"2f1b0c",x"321d0d",x"2d1a0b",x"321c0d",x"2d1a0b",x"2c190b",x"2d1a0b",x"211309",x"211309",x"180f07",x"1c1108",x"221508",x"301c0c",x"271809",x"271809",x"221608",x"201508",x"231609",x"211508",x"221608"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160f07",x"191008",x"201409",x"1c1108",x"25150a",x"150e07",x"150e07",x"160f07",x"1e1209",x"1e1209",x"201309",x"23150a",x"211409",x"201409",x"24150a",x"24160a",x"21140a",x"1b1108",x"1d1208",x"1b1108",x"1b1108",x"170e07",x"150e07",x"150e07",x"170f08",x"211309",x"241509",x"29170a",x"241509",x"251509",x"2a180b",x"2f1b0c",x"2a170a",x"261609",x"251509",x"211309",x"251509",x"27160a",x"201208",x"271509",x"241409",x"221308",x"261509",x"26160a",x"29170b",x"241509",x"2b180a",x"2f1a0b",x"3a200e",x"3c210f",x"391f0d",x"3a200e",x"311c0c",x"331d0d",x"26160a",x"21150a",x"2c190b",x"301b0c",x"2c190b",x"170f08",x"231409",x"2e1b0c",x"241509",x"473f36",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462b18",x"462b18",x"5d483a",x"5b483b",x"594436",x"4e4137",x"534133",x"594537",x"483e34",x"4e4035",x"46392f",x"463a31",x"503c2e",x"503e32",x"513f31",x"48362a",x"4f3d31",x"4f3c30",x"513b2d",x"543e2f",x"584031",x"513d2f",x"533d2f",x"513d31",x"513e32",x"493b30",x"564336",x"513f33",x"533f32",x"514034",x"5d4537",x"624836",x"543f32",x"5c4435",x"5c4537",x"5e4536",x"594537",x"5c4537",x"514236",x"614b3b",x"514337",x"4d3f35",x"4f4035",x"4e4035",x"4b3f35",x"504236",x"4e433a",x"56473b",x"4f4135",x"574437",x"524337",x"524337",x"524134",x"504237",x"503d2f",x"514236",x"504338",x"584538",x"594538",x"564437",x"584539",x"574539",x"54453a",x"524033",x"5c473a",x"5c483a",x"5e4636",x"554234",x"634837",x"564334",x"594334",x"544236",x"564437",x"564438",x"524135",x"4e4035",x"523d30",x"4c3c31",x"493a30",x"46392f",x"46382d",x"47362a",x"4e3829",x"45352a",x"413227",x"3c3128",x"433328",x"432f23",x"3d2e23",x"493324",x"483528",x"4a3527",x"513728",x"4a3324",x"5a3f2f",x"503828",x"4c3628",x"4c3b2f",x"503e32",x"574133",x"513f32",x"514034",x"4e4036",x"4f4136",x"504136",x"473d33",x"4b4137",x"453d35",x"492d19",x"150e07",x"150e07",x"150e07",x"150e07",x"44250f",x"150e07",x"2a1d11",x"2f2114",x"302215",x"312316",x"312215",x"332316",x"312214",x"2d1f13",x"2f2012",x"332315",x"342517",x"2d1f12",x"2f2013",x"322214",x"342416",x"332415",x"362618",x"352516",x"352516",x"332315",x"362516",x"28190c",x"2b1c0f",x"342316",x"342416",x"382718",x"382718",x"372718",x"3a2819",x"3c2a1b",x"392819",x"3c2b1b",x"412e1d",x"3d2b1b",x"3d2c1c",x"3a291a",x"3a291a",x"3a2819",x"382718",x"3a2819",x"332314",x"362516",x"3b291a",x"352416",x"2f2013",x"342315",x"3b291a",x"352416",x"342416",x"312214",x"332415",x"332315",x"312214",x"27180c",x"2d1d0f",x"332315",x"322315",x"362617",x"332316",x"302114",x"362617",x"382718",x"312214",x"332416",x"362618",x"3a281a",x"352517",x"2b1e12",x"2f2014",x"302114",x"24180e",x"302114",x"2d2012",x"312214",x"312214",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"40240f",x"40240f",x"39200d",x"1b1108",x"201408",x"211508",x"211508",x"1c1208",x"231608",x"1f1408",x"191007",x"170f07",x"191007",x"191007",x"1f1408",x"1d1308",x"160e07",x"170e07",x"1d1208",x"1b1207",x"1c1207",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"1a1007",x"190f07",x"4c2d11",x"301e0a",x"3f260e",x"36210b",x"3b240c",x"341f0b",x"321d0b",x"271709",x"2c1a0a",x"28170a",x"26170a",x"221509",x"231409",x"1f1308",x"201309",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"321c0c",x"1b1008",x"1b1008",x"231409",x"231509",x"211309",x"261509",x"301a0b",x"311b0b",x"39200e",x"371e0d",x"381f0d",x"3d210e",x"381f0d",x"3a200c",x"3a200d",x"452711",x"472812",x"502f16",x"4c2d13",x"523114",x"593616",x"502f13",x"4f2e15",x"513013",x"291a0a",x"321f0b",x"3a230d",x"3d250d",x"40280e",x"3f270e",x"40260e",x"3d250e",x"3f260e",x"3f250e",x"3c240e",x"3c240e",x"3b230f",x"3a230d",x"361f0d",x"39210c",x"341e0d",x"36200e",x"341f0d",x"341e0d",x"36200d",x"321d0c",x"2d1a0b",x"321d0c",x"311c0b",x"2c190b",x"2b180b",x"2c190b",x"2b180a",x"2a170a",x"2e1a0b",x"2e1a0b",x"2b190b",x"2d1a0b",x"2d190b",x"29170a",x"2d190b",x"2a180a",x"28170a",x"2d190b",x"29170a",x"261509",x"2a170a",x"2c180a",x"2a170a",x"281609",x"2a170a",x"2a170a",x"2a170a",x"2b180a",x"2a170a",x"2a170a",x"2c190b",x"2b190b",x"2a180b",x"2d190b",x"2a170a",x"2d190b",x"301b0b",x"2a180b",x"2a180b",x"2c190b",x"2c190b",x"301b0c",x"2e1a0b",x"301b0c",x"2f1b0c",x"2f1a0c",x"2a180b",x"27170a",x"241509",x"211309",x"211408",x"201509",x"221509",x"271809",x"271809",x"261709",x"291909",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"341d0d",x"3f2410",x"462912",x"452812",x"442611",x"442611",x"452711",x"432610",x"432510",x"442610",x"3d210e",x"41230f",x"402410",x"432611",x"432711",x"3d220f",x"40230f",x"3b200d",x"3f230f",x"462712",x"472811",x"452711",x"412611",x"442712",x"472812",x"462812",x"462812",x"4a2b14",x"462913",x"432712",x"472914",x"4b2b15",x"492a14",x"482913",x"472812",x"4b2b15",x"492a13",x"472812",x"482912",x"4c2c15",x"3f230f",x"381e0c",x"3d2310",x"492a13",x"4a2a13",x"472913",x"482913",x"412410",x"422510",x"472913",x"492a13",x"482913",x"452711",x"452711",x"422511",x"402410",x"452711",x"422510",x"3f230f",x"3a200e",x"402310",x"3c210e",x"412310",x"422510",x"361e0d",x"26160a",x"2b180b",x"27160a",x"150e07",x"473f36",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482f1f",x"412612",x"321e10",x"3a2212",x"362011",x"2d1b0f",x"2c1a0f",x"2b1a0e",x"402714",x"402614",x"402614",x"402615",x"3a2313",x"3a2314",x"392314",x"402817",x"352215",x"3b2515",x"392416",x"382417",x"3d2718",x"3a2618",x"3d2719",x"382416",x"362417",x"3a2518",x"392416",x"392517",x"3c2617",x"3d2516",x"3d2616",x"3f2818",x"442a18",x"3f2716",x"382314",x"442916",x"432916",x"412715",x"422917",x"422916",x"412816",x"412715",x"402616",x"412715",x"372213",x"3b2314",x"3a2313",x"3d2414",x"3b2413",x"3b2414",x"3e2615",x"3c2515",x"382112",x"3f2615",x"3d2515",x"382112",x"362012",x"382112",x"321e10",x"341f11",x"301d10",x"362011",x"341f11",x"3a2312",x"331e10",x"351f11",x"382313",x"3a2414",x"342013",x"3b2413",x"311f12",x"382213",x"3b2313",x"3a2313",x"3c2414",x"3e2615",x"382214",x"382313",x"3c2415",x"3d2515",x"3c2415",x"3c2414",x"3a2414",x"392414",x"3b2515",x"3b2414",x"3a2313",x"3c2414",x"382111",x"3b2311",x"3b2312",x"3a2111",x"3b2310",x"3e2411",x"3e2410",x"3d2410",x"3e2411",x"3e2412",x"3d2412",x"382110",x"392313",x"321e10",x"332011",x"2e1c0f",x"2f1d10",x"2f1d11",x"291a0e",x"4b3a2e",x"150e07",x"150e07",x"150e07",x"150e07",x"42240f",x"150e07",x"2d1f13",x"2e2013",x"2d2013",x"2e2013",x"322315",x"352617",x"332416",x"302114",x"352517",x"302114",x"302114",x"362517",x"382718",x"392818",x"352517",x"342416",x"372718",x"392819",x"3c2a1a",x"352516",x"302013",x"382717",x"372718",x"3a2819",x"3e2b1b",x"322315",x"372718",x"3c2a1b",x"402e1c",x"3b291a",x"3e2c1c",x"3d2b1b",x"372718",x"3a291a",x"412e1e",x"422e1d",x"412d1c",x"3c2b1b",x"3d2b1c",x"3d2b1a",x"3c2a1a",x"392819",x"372618",x"372718",x"382718",x"372718",x"352517",x"382718",x"322315",x"342416",x"332316",x"342415",x"332315",x"362617",x"372718",x"362617",x"352516",x"362517",x"342416",x"382718",x"392818",x"382718",x"342416",x"362617",x"332416",x"332416",x"2f2114",x"2d1f12",x"302114",x"2f2114",x"302214",x"291c11",x"2d1f12",x"2d1f12",x"2d1f12",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2d13",x"4e2c13",x"462911",x"3d230e",x"231608",x"201508",x"261809",x"231608",x"1f1408",x"241708",x"201408",x"191007",x"181007",x"191007",x"191007",x"1d1308",x"1c1208",x"170e07",x"170f07",x"1f1408",x"1a1107",x"1b1107",x"170f07",x"180f07",x"180f07",x"190f08",x"190f08",x"1a1108",x"191008",x"4a2d11",x"2f1e0a",x"2f1d0a",x"2c1c09",x"301e0a",x"2c1c09",x"251709",x"1b1108",x"251809",x"1a1107",x"1a1107",x"1a1107",x"150e07",x"170f07",x"1c1208",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"29170a",x"180f07",x"180f07",x"1a1008",x"170f07",x"1c1108",x"1b1108",x"24150a",x"251509",x"2f1b0c",x"361f0e",x"38200e",x"3b220f",x"3a200e",x"3c220f",x"3c210e",x"3d230e",x"3e230f",x"41240f",x"43270f",x"4a2b11",x"4d2e11",x"4d2d12",x"482910",x"492b11",x"2f1d0a",x"3a240c",x"38220c",x"40270d",x"3e260e",x"38220c",x"39220d",x"3e260e",x"42280e",x"3e250e",x"41270f",x"40260f",x"37210e",x"39220f",x"3e250f",x"351e0e",x"311d0c",x"341e0d",x"36200e",x"36200e",x"351f0c",x"301c0b",x"341e0d",x"321d0c",x"2d190a",x"2d190b",x"301c0c",x"301c0c",x"2f1c0c",x"321d0d",x"311c0c",x"2b180b",x"2d1a0b",x"2f1b0c",x"2d1a0b",x"2c190b",x"2b180b",x"2b180b",x"2b180b",x"2b190b",x"2e1a0b",x"2d190b",x"301b0c",x"29170a",x"2c190b",x"2b180a",x"2d190b",x"2f1a0c",x"301b0c",x"27160a",x"2e1a0b",x"2a180b",x"2b180b",x"29170a",x"261509",x"28170a",x"2c180b",x"2f1a0b",x"2a180b",x"2c190b",x"2f1a0c",x"28170a",x"2c190b",x"2b180a",x"2b180b",x"2c190b",x"2c190b",x"2d1a0c",x"29170a",x"26150a",x"231409",x"221409",x"1f1308",x"201409",x"241609",x"211509",x"251709",x"261709",x"281909",x"281809",x"281809",x"000000"),
(x"150e07",x"150e07",x"150e07",x"180f07",x"231409",x"2e190b",x"341d0d",x"331d0d",x"361f0e",x"351e0e",x"3b2210",x"422611",x"3e2410",x"3f2411",x"3c2310",x"37200e",x"3a210f",x"3a210f",x"39200f",x"3a200e",x"371f0d",x"321c0c",x"331c0c",x"39200e",x"3b220f",x"371f0d",x"361e0d",x"371f0e",x"381f0e",x"341d0d",x"331c0c",x"351d0d",x"361e0d",x"361d0d",x"341d0d",x"402411",x"3b220f",x"351e0e",x"341d0d",x"3b2310",x"3b2210",x"3b220f",x"422612",x"3a2310",x"321c0d",x"301c0c",x"372210",x"392310",x"3a2210",x"38210f",x"38200e",x"38200f",x"37210f",x"3a210f",x"38200f",x"3b2310",x"3a210f",x"3c2310",x"3b220f",x"351e0e",x"381f0e",x"361e0d",x"2e1a0b",x"2d190b",x"301b0b",x"311b0c",x"381f0e",x"39200e",x"38200e",x"391f0e",x"351e0d",x"2e1a0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412612",x"321e10",x"3a2212",x"362011",x"2d1b0f",x"2c1a0f",x"2b1a0e",x"402714",x"402614",x"402614",x"402615",x"3a2313",x"3a2314",x"392314",x"402817",x"352215",x"3b2515",x"392416",x"382417",x"3d2718",x"3a2618",x"3d2719",x"382416",x"362417",x"3a2518",x"392416",x"392517",x"3c2617",x"3d2516",x"3d2616",x"3f2818",x"442a18",x"3f2716",x"382314",x"442916",x"432916",x"412715",x"422917",x"422916",x"412816",x"412715",x"402616",x"412715",x"372213",x"3b2314",x"3a2313",x"3d2414",x"3b2413",x"3b2414",x"3e2615",x"3c2515",x"382112",x"3f2615",x"3d2515",x"382112",x"362012",x"382112",x"321e10",x"341f11",x"301d10",x"362011",x"341f11",x"3a2312",x"331e10",x"351f11",x"382313",x"3a2414",x"342013",x"3b2413",x"311f12",x"382213",x"3b2313",x"3a2313",x"3c2414",x"3e2615",x"382214",x"382313",x"3c2415",x"3d2515",x"3c2415",x"3c2414",x"3a2414",x"392414",x"3b2515",x"3b2414",x"3a2313",x"3c2414",x"382111",x"3b2311",x"3b2312",x"3a2111",x"3b2310",x"3e2411",x"3e2410",x"3d2410",x"3e2411",x"3e2412",x"3d2412",x"382110",x"392313",x"321e10",x"332011",x"2e1c0f",x"2f1d10",x"2f1d11",x"291a0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200d",x"150e07",x"2a1d11",x"2d1f12",x"2e1f13",x"312214",x"322315",x"302114",x"2e2013",x"342516",x"2f2014",x"342416",x"372718",x"3a2919",x"342416",x"352517",x"3b291a",x"392819",x"3d2b1b",x"3d2b1c",x"3d2b1b",x"3c2a1a",x"3e2b1b",x"3f2c1c",x"382718",x"3b2919",x"3a2919",x"3d2b1b",x"3c2a1a",x"3b2919",x"3f2c1c",x"402d1d",x"392819",x"392819",x"3a2819",x"392819",x"3a2919",x"422e1d",x"3b2919",x"3c2a1a",x"3f2d1c",x"3f2d1c",x"3f2d1c",x"3b2a1a",x"3a2919",x"332416",x"342416",x"352517",x"322416",x"362617",x"382819",x"362618",x"322316",x"332416",x"322315",x"3b291a",x"382718",x"382718",x"362517",x"352516",x"352516",x"382718",x"332416",x"362617",x"362517",x"382718",x"362617",x"352517",x"362517",x"312215",x"2e2013",x"332315",x"342416",x"2f2114",x"352517",x"322215",x"322215",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2911",x"512e15",x"512e14",x"41260f",x"39220f",x"1a1107",x"1f1408",x"231608",x"221608",x"1e1308",x"241708",x"201408",x"1a1107",x"1a1107",x"191007",x"1a1107",x"1b1108",x"1a1107",x"170f07",x"170f07",x"1f1408",x"1a1007",x"1a1107",x"180f07",x"180f07",x"190f08",x"191008",x"191008",x"191008",x"191008",x"41270f",x"32200a",x"2e1d0a",x"2c1c09",x"2c1c09",x"281a09",x"231608",x"1c1208",x"221508",x"170f07",x"191007",x"191007",x"150e07",x"160f07",x"1b1108",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"191008",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"241509",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"1b1008",x"1d1108",x"261509",x"2d1a0b",x"321c0c",x"3a210e",x"37200e",x"422711",x"3c2310",x"412711",x"432711",x"462912",x"492b13",x"4c2d13",x"4d2e11",x"462a11",x"452911",x"4b2d12",x"331f0b",x"311d0b",x"35200c",x"38210d",x"35200c",x"3a230d",x"341f0c",x"3d250e",x"3d240d",x"3e250d",x"39220c",x"38210d",x"3f250e",x"3a230c",x"3a220d",x"3b230d",x"351f0d",x"36210d",x"331e0d",x"39220e",x"37210e",x"321d0c",x"311d0d",x"351f0d",x"2d1a0c",x"2d1b0c",x"27180b",x"2d1c0d",x"2d1c0d",x"2f1b0c",x"2b190b",x"2b190b",x"2e1b0c",x"2a180b",x"2c190b",x"2c1a0c",x"2f1c0d",x"2d1a0c",x"28170b",x"2d1a0c",x"2c180b",x"2a180a",x"2e1a0b",x"2c180a",x"2c190b",x"2e1a0b",x"2b180b",x"2d190b",x"2e1a0c",x"2e1a0b",x"2e1a0b",x"29180a",x"2d190b",x"2b180a",x"29170a",x"27160a",x"2b180a",x"2d190b",x"301b0c",x"2c190b",x"301c0c",x"2c190b",x"2b180b",x"271609",x"29160a",x"29170a",x"2a170a",x"28160a",x"26160a",x"231409",x"231309",x"29170a",x"1c1108",x"211308",x"211409",x"291909",x"241509",x"241609",x"271809",x"271809",x"2a1a09",x"35200c"),
(x"150e07",x"150e07",x"150e07",x"1d1108",x"2e1a0b",x"331d0d",x"3a210f",x"381f0e",x"3a210f",x"3a210f",x"3e2410",x"39200e",x"422611",x"3b210f",x"3a200e",x"3b200e",x"381f0d",x"361e0d",x"341d0c",x"341d0c",x"341d0c",x"351c0c",x"301a0b",x"321b0b",x"311b0b",x"2f1a0b",x"361e0d",x"3b200e",x"3c220f",x"381f0e",x"39200e",x"361e0d",x"321b0b",x"381e0d",x"381e0d",x"381f0d",x"3a200e",x"341d0d",x"371f0e",x"341d0d",x"361e0d",x"361e0e",x"2f190a",x"321b0b",x"3b210f",x"422712",x"3e2411",x"3b2411",x"452914",x"3e2712",x"3a2512",x"3a2310",x"37200f",x"37200e",x"381f0e",x"3b210f",x"3c220f",x"3d2210",x"3b220f",x"38200e",x"3f2410",x"3d2410",x"3f2410",x"3c220f",x"3c220f",x"3c230f",x"3f2411",x"3c230f",x"402511",x"3b2210",x"3c230f",x"371f0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"452813",x"150e07",x"2c1e12",x"2d2013",x"312215",x"302215",x"372719",x"342517",x"372819",x"392919",x"322316",x"372719",x"3e2d1d",x"3f2d1d",x"3d2c1c",x"362618",x"39291a",x"3d2b1c",x"3f2d1c",x"382718",x"3d2b1b",x"3c2a1b",x"3a2919",x"382718",x"352516",x"362617",x"362516",x"362617",x"392818",x"352415",x"362718",x"3c2a1a",x"402e1c",x"3d2b1b",x"3e2b1b",x"402d1d",x"3d2b1c",x"453120",x"402e1e",x"3d2c1c",x"3a291a",x"392919",x"3a291a",x"3c2a1b",x"38281a",x"3c2b1c",x"3e2d1d",x"3f2c1c",x"412f1f",x"362618",x"362617",x"362517",x"382819",x"392819",x"382617",x"362517",x"2f2114",x"312215",x"2f2113",x"312214",x"312214",x"322214",x"332416",x"322315",x"332416",x"3b291a",x"362617",x"382719",x"2e2013",x"362718",x"362719",x"372719",x"362618",x"332416",x"302114",x"332416",x"332416",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462811",x"42250f",x"543115",x"482911",x"4a2911",x"38200e",x"231609",x"3c2410",x"211508",x"231608",x"211508",x"221608",x"221608",x"241708",x"211508",x"1f1408",x"1a1107",x"1a1107",x"191007",x"191007",x"191007",x"170e07",x"180f07",x"1c1208",x"1a1007",x"1a1007",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"452910",x"2c1c09",x"2f1d0a",x"2b1b09",x"281909",x"241708",x"231608",x"221508",x"1f1408",x"160e07",x"180f07",x"180f07",x"160e07",x"170f07",x"1a1107",x"170f07",x"180f08",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"190f08",x"180f08",x"231409",x"180f07",x"180f07",x"170f07",x"170f07",x"180f07",x"170f07",x"170f07",x"1a1008",x"27160a",x"2f1c0c",x"341d0d",x"311c0c",x"361e0e",x"3a200e",x"3f250f",x"3e240f",x"3d230f",x"3b210e",x"41260f",x"3d230e",x"3f250d",x"3d240d",x"44280e",x"4a2c12",x"2b1a0a",x"2f1d0a",x"321f0a",x"321e0b",x"331f0a",x"351f0b",x"35200b",x"331e0b",x"331e0b",x"341f0c",x"38210c",x"351f0c",x"38220c",x"39220c",x"3a230d",x"351f0c",x"36200c",x"321d0c",x"321c0c",x"2d1a0b",x"2d1a0b",x"261509",x"211308",x"2b180b",x"28180b",x"2d1a0c",x"2b1a0c",x"2a1a0c",x"2c1a0c",x"2f1c0d",x"2a190b",x"2a180b",x"27170a",x"28170a",x"24150a",x"27160a",x"29180b",x"25160a",x"2b190b",x"2b190b",x"2b190b",x"2f1c0c",x"2d1a0c",x"28170a",x"2d1a0c",x"311c0d",x"2d1a0c",x"2f1b0c",x"301c0d",x"2d1a0c",x"2e1b0c",x"2a180b",x"2a180b",x"2b190b",x"2c190b",x"28170a",x"2a180a",x"251509",x"28170a",x"2e1a0c",x"26160a",x"27160a",x"2a180a",x"301b0c",x"2d1a0b",x"2c190b",x"29170a",x"2b190b",x"201309",x"29180b",x"27160a",x"221409",x"241509",x"261609",x"241609",x"24150a",x"271809",x"251609",x"251609",x"261809",x"301d0a",x"35200c"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2e1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a220f",x"37200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"462813",x"150e07",x"221508",x"261a0f",x"291c10",x"2d2013",x"302214",x"2e2013",x"312215",x"332416",x"362719",x"3a291a",x"362718",x"392819",x"392819",x"3d2b1c",x"382718",x"372617",x"372617",x"372617",x"382819",x"3a2819",x"3a291a",x"3d2b1b",x"382718",x"382718",x"362617",x"3a2919",x"3c2a1a",x"362617",x"342416",x"382717",x"372617",x"342314",x"2a1a09",x"382818",x"382719",x"412e1e",x"362618",x"3a2919",x"362618",x"372718",x"3e2c1d",x"3d2b1c",x"352617",x"3b2a1a",x"3f2d1d",x"3b2a1b",x"362617",x"382718",x"312214",x"312114",x"362617",x"362618",x"3c2a1b",x"3c2a1b",x"322315",x"2f2013",x"302114",x"2a1d11",x"342417",x"302214",x"312114",x"2f2013",x"322315",x"291b0f",x"241608",x"2f2113",x"372618",x"342416",x"382819",x"312214",x"332316",x"312215",x"342517",x"2e2014",x"2e2014",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2e15",x"4b2a12",x"432610",x"42250f",x"42250f",x"543115",x"361f0b",x"26170a",x"27180a",x"39200e",x"251709",x"211508",x"1f1408",x"211508",x"221608",x"231608",x"251708",x"1d1308",x"1b1108",x"170f07",x"180f07",x"170f07",x"180f07",x"160f07",x"170f07",x"1b1007",x"190f08",x"1a1008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"3f250f",x"281909",x"281909",x"291a09",x"231608",x"1f1408",x"1b1108",x"181007",x"1c1208",x"150e07",x"160f07",x"170f07",x"160e07",x"180f07",x"191007",x"180f07",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"241509",x"2f1a0c",x"2e1b0c",x"311c0d",x"2f1b0c",x"2e190b",x"321d0d",x"2b180b",x"301a0b",x"26160a",x"211409",x"2e1a0b",x"321c0c",x"341d0c",x"3c230e",x"3a210e",x"3d240e",x"3c230f",x"452812",x"3f240f",x"3e240f",x"452810",x"452810",x"452710",x"442811",x"2a1909",x"2b1b09",x"2b1a0a",x"2d1b0a",x"2d1b0a",x"2a1809",x"2f1b0a",x"2b1a09",x"331e0b",x"311d0a",x"2f1c0b",x"2b190a",x"331e0c",x"2f1c0b",x"311c0c",x"321e0c",x"2a180b",x"331e0c",x"301b0b",x"2c190b",x"26160a",x"251509",x"231409",x"251509",x"28170a",x"27170a",x"26160a",x"24150a",x"2a180b",x"28170a",x"221409",x"28180b",x"2a190b",x"231509",x"1e1208",x"26160a",x"2c190b",x"28180b",x"2d1b0c",x"2f1b0c",x"2d1a0c",x"2d1a0c",x"2f1c0d",x"29180b",x"2d1a0c",x"2e1b0c",x"2f1b0c",x"2c190b",x"2e1a0c",x"2d1a0c",x"311c0d",x"28170a",x"2c1a0c",x"2b190b",x"2d1a0c",x"29180b",x"25150a",x"2b190b",x"2a180b",x"28170a",x"2b190b",x"29170a",x"2a180a",x"29170a",x"2b180b",x"241509",x"26160a",x"211309",x"1f1208",x"261509",x"231409",x"1f1208",x"201309",x"25150a",x"1e1208",x"1f1308",x"231509",x"231509",x"24160a",x"2f1d0b",x"311f0b",x"35200c"),
(x"150e07",x"150e07",x"150e07",x"1e1209",x"39210f",x"150e07",x"251509",x"301a0b",x"261509",x"351b0b",x"331a0b",x"331b0b",x"321b0b",x"331b0b",x"381f0d",x"381e0d",x"361e0c",x"371e0d",x"2e190b",x"2c180a",x"2d170a",x"2d170a",x"2d170a",x"281408",x"2a1609",x"391f0d",x"3d210e",x"3a200e",x"3b210e",x"3b200d",x"351d0c",x"3a1f0d",x"391f0d",x"341d0c",x"381f0d",x"3b200d",x"351d0c",x"391f0d",x"3a200e",x"3a210e",x"361e0d",x"381f0e",x"3d230f",x"371f0e",x"3b210f",x"412411",x"3f2410",x"3f2511",x"412511",x"3e2310",x"422511",x"3e2310",x"3e2310",x"3a210f",x"412511",x"3f2410",x"3f2410",x"402411",x"3b210f",x"3e2310",x"3d220f",x"412511",x"3f2411",x"3e2310",x"3b200e",x"3b200e",x"3d220f",x"27170a",x"432611",x"150e07",x"3d2210",x"36200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"432713",x"150e07",x"2d1f12",x"271b0f",x"2c1d11",x"281b0f",x"2a1c10",x"2a1c11",x"2a1d11",x"302114",x"302114",x"322315",x"362618",x"372718",x"352517",x"3e2c1c",x"382819",x"3d2b1b",x"3b291a",x"44311f",x"3d2c1c",x"3c2a1b",x"3e2c1c",x"402d1c",x"402d1d",x"372618",x"362617",x"3e2b1b",x"3b2a1a",x"3f2d1c",x"3c2a1b",x"43301f",x"3b2919",x"3e2c1a",x"3a2819",x"362517",x"382717",x"3a2818",x"322214",x"322315",x"342416",x"362617",x"362517",x"3a291a",x"332316",x"382819",x"3d2a1b",x"3d2b1b",x"3a291a",x"382718",x"382718",x"3b2a1b",x"3c2b1b",x"382719",x"3c2a1b",x"372618",x"382819",x"362618",x"352517",x"362617",x"362618",x"322316",x"352517",x"352517",x"322214",x"382717",x"2d1e12",x"2c1e12",x"2c1e11",x"2d1f12",x"2f2012",x"312214",x"291c10",x"291c11",x"2b1d11",x"2d1f13",x"2d1f13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492a13",x"553218",x"4f2e15",x"472912",x"3f230f",x"41250e",x"3c240e",x"2d1b0a",x"2e1c0b",x"241609",x"3d230f",x"211508",x"231608",x"231608",x"241608",x"231608",x"201508",x"1e1308",x"1f1408",x"1b1108",x"191007",x"160f07",x"160e07",x"160e07",x"160f07",x"170f07",x"180f08",x"180f08",x"180f07",x"191008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"3b220e",x"231608",x"261809",x"271909",x"241608",x"221508",x"160f07",x"160e07",x"160f07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"190f07",x"190f08",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"3c220f",x"2c190b",x"2c190b",x"26160a",x"2d190b",x"2c180b",x"281609",x"2d180a",x"2d190b",x"2e190b",x"321c0c",x"2b190b",x"331c0b",x"38200c",x"351e0b",x"361d0b",x"351c0b",x"381f0c",x"381f0d",x"3b220d",x"3a210c",x"3e240e",x"43270e",x"3d230d",x"42260f",x"191007",x"1d1107",x"1f1208",x"1e1107",x"1f1208",x"28170a",x"221509",x"29190a",x"251609",x"2a1909",x"28180a",x"2c190a",x"29180a",x"29180a",x"281709",x"281609",x"261609",x"26150a",x"271609",x"29180b",x"221409",x"27160a",x"27160a",x"28170a",x"29180b",x"24150a",x"27170a",x"27170b",x"2a180b",x"25150a",x"27160a",x"26160a",x"1f1309",x"25160a",x"211409",x"26160a",x"28170b",x"27170a",x"29180b",x"28170b",x"28170a",x"2d1a0c",x"29180b",x"27160a",x"27160a",x"27160a",x"29180b",x"2a180b",x"2b190b",x"2d1a0c",x"2a180b",x"27160a",x"251509",x"251509",x"27160a",x"27160a",x"27160a",x"26160a",x"261609",x"28160a",x"28160a",x"231409",x"231409",x"251509",x"241409",x"211309",x"1f1208",x"201309",x"231409",x"241509",x"1e1208",x"1d1108",x"1d1208",x"1e1208",x"1f1208",x"1e1208",x"1e1208",x"231509",x"2a1a09",x"2d1b0b",x"2f1d0b",x"35200c"),
(x"150e07",x"150e07",x"150e07",x"170f07",x"3f2411",x"191008",x"191008",x"432611",x"402410",x"472912",x"3d220f",x"361e0c",x"361d0d",x"391f0d",x"3c200e",x"3b200e",x"3b200e",x"391f0e",x"3e2310",x"402510",x"402511",x"3e230f",x"3a1f0d",x"381f0d",x"3d220f",x"39200d",x"3c200e",x"3f240f",x"432510",x"402410",x"3f2410",x"3a210f",x"3c210f",x"3a200e",x"3c220f",x"3c220f",x"3c210f",x"412511",x"452813",x"402512",x"3d2411",x"412612",x"3d2411",x"402512",x"422612",x"422611",x"432712",x"442712",x"452914",x"422712",x"3f2411",x"412511",x"412511",x"432712",x"432712",x"412511",x"402411",x"3d220f",x"371e0d",x"3e220f",x"3b210f",x"3d2310",x"422611",x"3f2410",x"472812",x"3b210f",x"3e220f",x"180f08",x"2a180b",x"150e07",x"3c220f",x"36200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"432711",x"150e07",x"2e2114",x"2f2115",x"2b1d12",x"302215",x"332416",x"362618",x"342517",x"382718",x"3b2a1b",x"392819",x"3c2b1c",x"3c2b1c",x"382719",x"362618",x"382718",x"3a2819",x"291a0b",x"382618",x"382718",x"3c2a1a",x"3d2b1b",x"402e1e",x"3e2c1c",x"3a291a",x"412f1f",x"382819",x"412f1f",x"412e1e",x"402d1d",x"3f2c1b",x"3a2918",x"3f2d1d",x"3e2c1c",x"43301f",x"3c2a1b",x"3f2d1d",x"402d1d",x"3d2b1c",x"3a291a",x"3a2819",x"3f2d1d",x"3d2c1c",x"433120",x"443120",x"3e2c1c",x"392819",x"3b291a",x"342416",x"26180a",x"342416",x"392819",x"3c2a1a",x"3b291a",x"3c2b1c",x"3a2819",x"3a291a",x"39291a",x"362617",x"352618",x"3c2a1b",x"39281a",x"322315",x"332314",x"362718",x"352617",x"342416",x"352517",x"3a2a1a",x"312215",x"322416",x"312215",x"322315",x"302114",x"312216",x"312216",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"42240f",x"41220e",x"513016",x"442812",x"2b1a0b",x"462913",x"2e1d0a",x"2f1d0b",x"311e0b",x"321e0c",x"241609",x"3c230f",x"1f1408",x"231608",x"221508",x"231608",x"201408",x"1f1408",x"1f1408",x"1a1107",x"191007",x"170f07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"482a10",x"271909",x"271809",x"281909",x"271909",x"181007",x"150e07",x"150e07",x"150e07",x"160e07",x"180f07",x"1d1208",x"1b1107",x"1c1107",x"1c1107",x"1c1208",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"3b210f",x"26160a",x"2b190b",x"2f1b0c",x"2d1a0b",x"261509",x"2b1809",x"351e0c",x"38200d",x"361f0c",x"3c230e",x"3c230f",x"351f0d",x"3e240e",x"3e240f",x"3b210d",x"381f0d",x"381f0c",x"391f0d",x"3b220d",x"3c220e",x"472911",x"43270f",x"482911",x"482912",x"1a1107",x"191107",x"1d1108",x"170f07",x"170f07",x"1b1008",x"1c1108",x"1d1108",x"221409",x"27170a",x"27180a",x"27170a",x"2d1a0a",x"241609",x"28180a",x"261609",x"29180a",x"201409",x"27170b",x"28190b",x"25160a",x"24150a",x"23150a",x"22150a",x"23150a",x"211409",x"211409",x"27170b",x"28170b",x"24150a",x"25160a",x"221409",x"221409",x"25160a",x"24150a",x"26160a",x"241509",x"251509",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"26160a",x"241509",x"26160a",x"26160a",x"251509",x"27160a",x"26160a",x"241509",x"231409",x"201309",x"25160a",x"201309",x"231409",x"241509",x"221409",x"241409",x"261509",x"231409",x"231409",x"221409",x"231409",x"231409",x"211309",x"1e1208",x"201208",x"1e1208",x"231409",x"201309",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1f1309",x"1f1208",x"231509",x"2b1b0a",x"2c1b0a",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"432713",x"150e07",x"150e07",x"150e07",x"201308",x"28170a",x"341d0d",x"3a1f0e",x"311b0b",x"2e190a",x"321b0b",x"321c0c",x"381f0d",x"381f0e",x"361e0d",x"38200e",x"351d0d",x"3a200e",x"371e0d",x"361e0d",x"341d0d",x"341d0d",x"371e0d",x"331c0c",x"371e0d",x"331c0c",x"371e0d",x"361e0d",x"381f0d",x"371f0d",x"39200e",x"3a210f",x"3d2310",x"371f0e",x"351d0d",x"341d0d",x"341d0d",x"331c0c",x"2f1a0c",x"351f0e",x"3a210f",x"3e2411",x"3d2410",x"3c2310",x"3d2310",x"39200f",x"381f0e",x"381f0d",x"351d0d",x"361e0d",x"381f0e",x"3b210f",x"3b220f",x"38200f",x"341d0d",x"3a210f",x"3a210f",x"331d0d",x"3b200e",x"351d0d",x"3d220e",x"150e07",x"180f07",x"1c1108",x"1d1108",x"201208",x"3b210f",x"392110",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"402310",x"19120b",x"322519",x"2e2216",x"312417",x"302114",x"302214",x"312215",x"322215",x"382718",x"302213",x"312214",x"3a2a1a",x"3e2b1b",x"392819",x"392819",x"372718",x"3b2919",x"362517",x"3c2a1b",x"3a2919",x"382718",x"412e1d",x"453120",x"3a291a",x"3c2a1b",x"43301f",x"42301f",x"422f1e",x"463321",x"493422",x"3b2919",x"43301f",x"412e1d",x"3f2d1c",x"392819",x"3d2b1b",x"3a2919",x"3b2a1a",x"392819",x"3c2a1b",x"39281a",x"382817",x"3e2c1b",x"412e1e",x"3b2919",x"3a291a",x"3e2c1c",x"392819",x"3b2919",x"3d2a1b",x"332416",x"342416",x"3b291a",x"3d2b1c",x"3f2d1c",x"372718",x"332416",x"3f2d1d",x"3a2a1a",x"3b2a1b",x"3d2b1c",x"362618",x"332414",x"3a281a",x"382718",x"362617",x"312215",x"312214",x"322315",x"322315",x"302114",x"332416",x"352517",x"2e2113",x"322416",x"322416",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1108",x"1d1108",x"1f1309",x"2c190a",x"2f1b0b",x"412611",x"2d1c0a",x"2c1b0a",x"2c1b0a",x"301d0b",x"291909",x"38210f",x"201508",x"1f1408",x"201508",x"211508",x"1f1408",x"1f1408",x"1e1308",x"1c1208",x"1a1107",x"170f07",x"150e07",x"160e07",x"160e07",x"170f07",x"181007",x"180f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"462910",x"2e1d0a",x"2e1d0a",x"2c1c09",x"251709",x"1c1208",x"191007",x"150e07",x"160e07",x"180f07",x"1a1107",x"181007",x"251708",x"1f1309",x"1b1108",x"1d1208",x"1d1208",x"1d1208",x"1c1108",x"1d1108",x"1d1208",x"1d1208",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"3f2410",x"2f1b0c",x"311c0c",x"2e1b0c",x"2d190b",x"2e1a0b",x"321c0b",x"341d0b",x"371f0d",x"39210e",x"38210d",x"3a210e",x"361f0d",x"351e0d",x"3b210e",x"381f0d",x"3b210d",x"371e0c",x"381f0c",x"3a200c",x"45280f",x"43270f",x"4a2b11",x"4c2d12",x"4a2a11",x"1c1108",x"160f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f08",x"191008",x"1d1208",x"201309",x"1e1208",x"201409",x"231509",x"2a1a09",x"25170a",x"241609",x"201309",x"211409",x"1e1208",x"1d1108",x"1f1209",x"1f1309",x"1f1309",x"211409",x"201309",x"211409",x"201309",x"1f1309",x"1e1208",x"1f1208",x"201309",x"1f1208",x"1f1208",x"211309",x"221409",x"201309",x"211309",x"24150a",x"231509",x"201309",x"201309",x"201208",x"1f1208",x"201208",x"201208",x"201308",x"1f1208",x"1f1208",x"211309",x"201309",x"201309",x"211309",x"201308",x"1e1208",x"1f1208",x"1f1308",x"1d1108",x"1c1008",x"1c1008",x"1d1208",x"1e1208",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"201309",x"1e1208",x"1f1208",x"1f1208",x"201408",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"26170b",x"402511",x"150e07",x"261609",x"321b0c",x"361e0d",x"38200e",x"371f0d",x"39200e",x"351e0d",x"3e230f",x"3d220f",x"3a200e",x"381f0e",x"3c220f",x"39200f",x"3b2210",x"3d2410",x"3a210f",x"3a210f",x"3a210f",x"3c220f",x"3a210f",x"3c220f",x"39200e",x"381f0e",x"351d0c",x"3b200e",x"341c0c",x"3a200e",x"3e2310",x"3c220f",x"351e0d",x"311c0c",x"38200e",x"371e0d",x"381f0e",x"38200e",x"371f0e",x"351e0e",x"3b2210",x"38200e",x"3d2310",x"3c2310",x"3c2310",x"412612",x"402512",x"3a210f",x"3b210f",x"3b2210",x"3d2310",x"3c2310",x"3d2411",x"38200e",x"3c2310",x"3a2210",x"3f2511",x"412410",x"402511",x"462813",x"422712",x"472914",x"180f08",x"392110",x"3d2411",x"3c2311",x"331e0e",x"3d220f",x"3a2210",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422511",x"251e17",x"392c20",x"3d2e22",x"36281c",x"322418",x"3b2a1b",x"3a291a",x"3b2a1b",x"392819",x"332314",x"332415",x"3d2c1c",x"3e2c1c",x"3b2a1a",x"3b2a1a",x"382818",x"3c2a1b",x"3d2c1c",x"3c2a1b",x"3f2d1d",x"3e2c1c",x"402e1d",x"3f2d1c",x"453220",x"3e2f1f",x"3e2f1f",x"493625",x"453221",x"453221",x"43301f",x"4a3724",x"453221",x"423020",x"453220",x"44311f",x"44311f",x"43301f",x"44301f",x"402e1e",x"3c2b1c",x"3b2919",x"3b2919",x"3a2818",x"453220",x"3c2b1b",x"3c2b1b",x"3f2c1c",x"3d2b1c",x"3e2c1c",x"412f1f",x"412e1e",x"3f2d1d",x"392819",x"3c2b1c",x"39291a",x"3f2e1f",x"413222",x"413221",x"423122",x"402f20",x"412f20",x"3c2c1d",x"413121",x"3f2f20",x"423121",x"38291c",x"352719",x"3a2b1c",x"3a2a1c",x"38291c",x"36271b",x"382a1c",x"322418",x"322418",x"34261a",x"34261a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"181007",x"181007",x"221509",x"301c0b",x"3a230d",x"41250f",x"2e1c0b",x"281909",x"25170a",x"28180a",x"261709",x"452913",x"2b1b09",x"201408",x"211508",x"201408",x"1e1308",x"1d1308",x"1c1208",x"191007",x"180f07",x"160e07",x"160e07",x"160e07",x"180f07",x"170f07",x"1b1107",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1208",x"1e1209",x"1e1209",x"1e1209",x"1e1209",x"4a2d12",x"311f0a",x"301f0a",x"2b1b09",x"221508",x"1e1308",x"1a1007",x"160e07",x"160f07",x"180f07",x"170f07",x"190f07",x"1e1308",x"191008",x"221509",x"201409",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1a1008",x"1b1008",x"1c1108",x"1d1208",x"1e1208",x"1c1108",x"3b210f",x"2a180b",x"27160a",x"29160a",x"28170a",x"311c0d",x"321d0c",x"311c0c",x"2d190b",x"38200d",x"311c0b",x"351e0c",x"381f0d",x"371f0d",x"3d230f",x"361f0d",x"3b220f",x"39200e",x"432710",x"3c220d",x"41260e",x"482a11",x"4b2c12",x"513014",x"4f3014",x"190f07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"190f08",x"190f07",x"191008",x"1a1008",x"1a1008",x"1d1208",x"201308",x"241609",x"241609",x"251709",x"221509",x"1f1208",x"1d1108",x"1f1309",x"1f1208",x"201309",x"201309",x"1f1208",x"201309",x"201409",x"201409",x"211409",x"201309",x"1f1209",x"1f1309",x"201309",x"201309",x"201309",x"201309",x"201309",x"211409",x"221409",x"211409",x"201309",x"231409",x"23150a",x"24150a",x"24150a",x"24150a",x"24150a",x"24160a",x"24160a",x"24160a",x"23150a",x"23150a",x"23150a",x"211409",x"211409",x"201309",x"201309",x"201309",x"1f1308",x"201309",x"211409",x"201309",x"1e1208",x"1e1108",x"1e1208",x"201309",x"201409",x"201309",x"201309",x"201309",x"1f1208",x"1d1108",x"1c1108",x"201309",x"201309",x"1d1108",x"1f1208",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"3d2310",x"150e07",x"2a180b",x"28170a",x"321c0c",x"301b0c",x"3b210e",x"351d0d",x"351d0c",x"301a0b",x"371e0d",x"361e0d",x"381f0e",x"361e0d",x"3c210f",x"402410",x"381f0e",x"3d220f",x"361e0d",x"3a210f",x"3a200e",x"341d0c",x"341d0c",x"351c0c",x"341c0c",x"351c0c",x"361d0c",x"31190b",x"291308",x"321a0b",x"371e0d",x"331c0c",x"321b0c",x"381f0d",x"371f0e",x"39200e",x"361f0d",x"38200e",x"361f0e",x"3d2310",x"3c220f",x"3d2310",x"3d220f",x"3c220f",x"402511",x"3a200f",x"3a210f",x"412511",x"3f2411",x"402511",x"3d220f",x"412612",x"3a2210",x"3f2411",x"3d230f",x"39200e",x"3b200e",x"3c210f",x"3d220f",x"3d2410",x"150e07",x"2a180b",x"351e0e",x"3d2411",x"3d2411",x"351f0e",x"39200e",x"341e0d",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"432611",x"29221c",x"3b2e22",x"392d22",x"3b2d20",x"3e2d1f",x"2f2216",x"382819",x"352618",x"3b2a1a",x"342416",x"3a281a",x"392819",x"392819",x"3a291a",x"3e2c1c",x"402d1c",x"3b2a1a",x"463220",x"412f1e",x"3e2c1b",x"3f2d1c",x"3b2a1a",x"412e1e",x"3f2d1d",x"402d1d",x"3e2c1c",x"3f2e1d",x"44311f",x"463221",x"463220",x"433322",x"3f2d1d",x"443120",x"463221",x"453220",x"433120",x"412e1e",x"423120",x"422f1e",x"453220",x"3e2c1c",x"3c2a1b",x"3e2c1c",x"3f2c1c",x"3f2c1c",x"3e2b1b",x"3a291a",x"3f2d1c",x"3e2c1c",x"3c2b1b",x"3b2b1c",x"3a291a",x"3f2e1e",x"3b2b1c",x"3d2d1d",x"3f2e1f",x"3d2c1d",x"402e1f",x"413121",x"3d2c1e",x"423121",x"3a2b1e",x"3d3021",x"3e2f20",x"3e2e1f",x"3d2d1f",x"423121",x"3b2d1f",x"3a2c1f",x"3b2c1f",x"392a1c",x"3a2c1e",x"3a2b1e",x"3f2f21",x"3a2c1f",x"3a2c1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1107",x"1a1107",x"251609",x"321c0b",x"3d240e",x"432711",x"27180a",x"2a190a",x"28180a",x"27180a",x"231509",x"472a11",x"1d1308",x"1f1408",x"201508",x"201408",x"1f1408",x"1c1208",x"1a1107",x"191007",x"150e07",x"150e07",x"160e07",x"160e07",x"181007",x"181007",x"1a1007",x"180f08",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1d1208",x"1d1209",x"1d1208",x"1e1209",x"1e1209",x"41270f",x"2c1c09",x"311f0a",x"281909",x"2c1c09",x"191007",x"1a1007",x"160e07",x"160f07",x"1b1107",x"191007",x"180f08",x"231609",x"191008",x"1f1309",x"1c1108",x"1f1308",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"3a200e",x"26160a",x"231409",x"261509",x"241509",x"2a180b",x"2e1b0b",x"2d1a0b",x"2c190b",x"311c0c",x"37200d",x"351e0d",x"321c0b",x"37200c",x"39210d",x"361e0d",x"37200d",x"361e0c",x"371f0c",x"38200d",x"3e240e",x"472a0f",x"45290f",x"4c2d12",x"492b11",x"25150a",x"28170a",x"29170a",x"26160a",x"29170a",x"28160a",x"26160a",x"28160a",x"28170a",x"2c180b",x"28160a",x"271509",x"27160a",x"29170b",x"2c190b",x"2b180b",x"2a180a",x"2a180a",x"26150a",x"211409",x"211309",x"211309",x"221409",x"24150a",x"26160a",x"26160a",x"27170b",x"27170a",x"26160a",x"27160a",x"27170a",x"251509",x"221308",x"221409",x"241509",x"27160a",x"27170b",x"27160a",x"25160a",x"25160a",x"25160a",x"221409",x"221409",x"241509",x"25160a",x"25160a",x"26170a",x"24150a",x"24150a",x"23150a",x"221409",x"211309",x"201309",x"201309",x"211309",x"26160a",x"27160a",x"28160a",x"2c190b",x"29170b",x"2a180b",x"29180b",x"201309",x"201309",x"1f1208",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"221409",x"191008",x"191008",x"180f08",x"180f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"3b2311",x"150e07",x"271609",x"2b180a",x"2f1a0c",x"2d1a0b",x"381f0e",x"331d0d",x"2f1b0c",x"341c0c",x"301b0b",x"2f1a0b",x"321b0b",x"321c0c",x"341d0d",x"3a210f",x"3b220f",x"3a200f",x"38200e",x"351e0d",x"351e0d",x"371e0d",x"351d0c",x"361e0d",x"351d0c",x"381e0d",x"351d0d",x"2e1a0b",x"311b0c",x"371f0d",x"321c0b",x"301a0b",x"341d0c",x"2e190b",x"2e190b",x"341d0d",x"321d0d",x"331d0d",x"351e0e",x"351e0e",x"351e0d",x"341d0d",x"2f1b0b",x"341d0d",x"341d0c",x"331c0c",x"2f1a0b",x"2d180a",x"251207",x"241207",x"261207",x"301a0b",x"331c0c",x"301b0b",x"311b0b",x"2d190b",x"311b0b",x"2f1a0b",x"341d0c",x"311b0b",x"150e07",x"241409",x"2b180a",x"2e190b",x"2b170a",x"281609",x"3c210f",x"321d0d",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442712",x"2b241d",x"3f3125",x"3e3024",x"362a20",x"3c2c1f",x"3b2a1b",x"352516",x"362718",x"3e2c1d",x"342517",x"342619",x"3b2c1c",x"402f1e",x"362719",x"39291a",x"3c2b1b",x"3b2a1a",x"3f2d1d",x"402e1e",x"412f1e",x"3c2a1a",x"3e2c1c",x"402e1e",x"3c2a1b",x"3f2d1d",x"3c2a1b",x"43301e",x"43301f",x"412f1e",x"453221",x"453120",x"453120",x"422f1e",x"473321",x"453220",x"473321",x"412e1c",x"422f1e",x"402d1d",x"3f2d1d",x"443221",x"402e1e",x"3e2c1c",x"42301f",x"3d2b1c",x"412e1d",x"412e1d",x"3f2d1d",x"3f2d1d",x"3e2d1e",x"3f2e1f",x"3f2e1f",x"42301f",x"423020",x"423121",x"3f2f20",x"423021",x"3f2e1f",x"392a1c",x"463424",x"3f2e20",x"3c2d20",x"3f2f21",x"3b2d1f",x"3f2f21",x"3c2d20",x"3b2c1f",x"3f2e20",x"3e2e1f",x"3d2d1f",x"3a2b1d",x"3d2f21",x"3a2c20",x"3d2f21",x"392b1f",x"392b1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1308",x"1f1308",x"201308",x"321c0b",x"371e0c",x"482a12",x"28180a",x"26160a",x"28180a",x"26170a",x"27170a",x"371f0d",x"191007",x"1d1208",x"1d1208",x"1c1208",x"1d1308",x"1d1208",x"1b1108",x"181007",x"170f07",x"150e07",x"160e07",x"160e07",x"160e07",x"170f07",x"191007",x"190f07",x"180f07",x"190f07",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"44270f",x"301e0a",x"2f1e0a",x"2e1d0a",x"221608",x"1c1208",x"160e07",x"160f07",x"170f07",x"181007",x"1b1107",x"1b1008",x"1b1108",x"201309",x"201409",x"1f1208",x"1e1208",x"1e1208",x"1b1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"331d0d",x"29180a",x"231509",x"2c190b",x"2b190b",x"2d190b",x"37200e",x"341e0d",x"37200e",x"341d0c",x"341d0c",x"311c0c",x"351f0d",x"29170a",x"301b0b",x"311c0c",x"351d0d",x"341e0c",x"351e0b",x"321d0c",x"3a220c",x"43270e",x"43270f",x"40260f",x"482a11",x"26160a",x"241509",x"241509",x"241509",x"231509",x"221309",x"221409",x"221409",x"211309",x"211309",x"201308",x"1f1208",x"201309",x"201309",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"201208",x"211309",x"221409",x"221409",x"231409",x"231509",x"221409",x"231409",x"221409",x"231409",x"231409",x"221309",x"211308",x"201208",x"1c0f07",x"1c1007",x"1d1007",x"221409",x"231409",x"221409",x"201308",x"201208",x"201308",x"211309",x"201309",x"201208",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1e1108",x"1d1108",x"1d1108",x"1f1208",x"201309",x"201309",x"211409",x"201309",x"211409",x"211409",x"211309",x"211409",x"201309",x"201309",x"1f1208",x"1f1209",x"1f1209",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"1a1008",x"1a1008",x"180f07",x"170f07",x"170f07",x"170f07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"3f2511",x"150e07",x"2b180b",x"2f1b0c",x"25150a",x"29170a",x"341d0d",x"39200e",x"3c220f",x"3e220f",x"3b210f",x"3a200e",x"3f2310",x"341d0d",x"3a200e",x"3c210f",x"3d230f",x"3b220f",x"3c220f",x"3c220f",x"381f0e",x"3d220f",x"3c210f",x"371e0d",x"381f0d",x"3d220f",x"3a200e",x"3a210f",x"371f0e",x"381f0e",x"351d0d",x"3e2310",x"371f0e",x"331d0d",x"3c220f",x"351e0d",x"371f0e",x"3a210f",x"3b210f",x"3c230f",x"3e2411",x"381f0e",x"3d2310",x"3f2310",x"3c2310",x"422611",x"432712",x"432712",x"412511",x"3e2310",x"3f2411",x"351e0d",x"3a200e",x"381f0e",x"39200e",x"381e0d",x"3a200d",x"371e0d",x"371d0c",x"3b200e",x"3e230f",x"150e07",x"301b0c",x"311b0c",x"2e1a0b",x"2a180b",x"39200e",x"311c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442712",x"2a231c",x"3b2f24",x"3b2e22",x"382b21",x"33271a",x"392819",x"342517",x"3f2d1d",x"402d1d",x"39281a",x"3b2a1b",x"3c2b1c",x"3c2b1d",x"38281a",x"3c2a1c",x"412f1e",x"402d1d",x"412f1d",x"3d2b1b",x"412e1d",x"44301f",x"3d2c1c",x"43301f",x"43301f",x"463220",x"463320",x"412e1e",x"402e1d",x"42301f",x"463220",x"483423",x"483423",x"443120",x"43301f",x"4a3523",x"483322",x"443120",x"43301e",x"43311f",x"443120",x"3f2d1d",x"3f2e1d",x"42301f",x"433120",x"382819",x"342416",x"3f2c1c",x"3c2b1b",x"3c2b1c",x"3f2d1e",x"3b2a1b",x"3f2e1e",x"402e1f",x"3f2e1f",x"423020",x"433222",x"453222",x"453323",x"3f2f20",x"413022",x"463424",x"403021",x"413122",x"403022",x"463526",x"403022",x"413022",x"433223",x"392b1f",x"382a1d",x"3a2c1f",x"362a1e",x"3b2d20",x"382b1f",x"3d2e21",x"3d2e21",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"28180a",x"28180a",x"27170a",x"3b220e",x"412611",x"482a12",x"28180b",x"251609",x"28180a",x"2c1a0a",x"28180a",x"3f240f",x"1f1308",x"1d1308",x"231608",x"1c1208",x"191107",x"1f1408",x"1a1107",x"191007",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"170f07",x"191007",x"170f07",x"180f07",x"191008",x"1b1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"472910",x"2c1c09",x"311f0a",x"261809",x"261809",x"180f07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f07",x"1a0f08",x"1c1208",x"1d1208",x"1b1108",x"1c1108",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1b1008",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1b1108",x"351d0d",x"241509",x"231409",x"28170a",x"2c190b",x"2d190b",x"331d0d",x"311c0c",x"351e0c",x"351e0d",x"331d0d",x"361f0d",x"24150a",x"27160a",x"221409",x"2f1a0c",x"341d0c",x"37200d",x"311c0b",x"321d0c",x"38200d",x"3f250e",x"3f250f",x"472910",x"4b2c11",x"27170a",x"27170a",x"25160a",x"24150a",x"231409",x"231509",x"221409",x"211309",x"221409",x"221409",x"211409",x"221409",x"211309",x"201309",x"201309",x"211409",x"201309",x"211409",x"211309",x"211409",x"231509",x"231409",x"221409",x"24150a",x"24150a",x"231409",x"25160a",x"25160a",x"26160a",x"28170b",x"28170b",x"28170b",x"27170a",x"27170a",x"27170b",x"241409",x"241509",x"241509",x"231409",x"211309",x"221409",x"211309",x"201308",x"211409",x"211309",x"201309",x"211409",x"201309",x"201309",x"201309",x"201309",x"201308",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1d1108",x"1b1008",x"1b1108",x"1a1008",x"1a1008",x"180f07",x"180f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"170f07",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"29180b",x"402512",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1a0c",x"341e0e",x"402512",x"37200f",x"3c2310",x"3d2310",x"3a210f",x"3e2411",x"3c2310",x"3e2411",x"371f0e",x"371e0d",x"3b210f",x"3a210f",x"3c2210",x"38200e",x"3f2310",x"3d2310",x"3b2210",x"3a200f",x"3b210f",x"39200e",x"351d0d",x"39200f",x"3f2410",x"3a200e",x"3c2310",x"3a2210",x"3a210f",x"341d0d",x"311b0b",x"351d0d",x"38200e",x"3a210f",x"3c220f",x"361e0d",x"361e0d",x"39200e",x"3c220f",x"3c2310",x"3c220f",x"371f0e",x"3c2310",x"3e2310",x"3d220f",x"381f0d",x"371f0d",x"361e0d",x"351d0d",x"3a200e",x"331b0b",x"361d0c",x"3d220f",x"3a210e",x"371e0d",x"3d220e",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"371f0e",x"2a170a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"492913",x"382b20",x"523d2c",x"533e2c",x"5b4430",x"5e452f",x"644932",x"5f462e",x"634931",x"5c412c",x"60442e",x"644931",x"674b32",x"6a4d34",x"70553a",x"6a4d34",x"694c34",x"6c4f37",x"715239",x"6b4e35",x"725438",x"61452e",x"63482f",x"694b32",x"684c33",x"6f5136",x"644830",x"5d432c",x"5d432d",x"61452e",x"644931",x"62472f",x"553e29",x"553e29",x"59412b",x"553c27",x"5c432d",x"573f29",x"5d4530",x"5b432d",x"563f2a",x"533c27",x"4e3824",x"624630",x"674b33",x"654932",x"674c35",x"634931",x"604630",x"71543a",x"6e5238",x"644932",x"644931",x"624730",x"6c4f36",x"6b4e36",x"674b34",x"654b33",x"624731",x"5c432d",x"614831",x"654a33",x"6c4f37",x"5d4630",x"5d452f",x"5f4630",x"604731",x"57402c",x"614832",x"58412d",x"624833",x"5b442f",x"5a432f",x"563f2b",x"4f3927",x"4f3b29",x"4f3b29",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1b0b",x"2d1b0b",x"341f0c",x"40250f",x"3f230e",x"452610",x"261709",x"241509",x"251609",x"26170a",x"27160a",x"40240f",x"201408",x"231608",x"1e1308",x"1c1208",x"1c1208",x"1a1107",x"1d1308",x"181007",x"191007",x"160f07",x"180f07",x"170e07",x"160e07",x"160e07",x"180f07",x"190f07",x"190f07",x"1d1208",x"1c1107",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"1c1108",x"482b11",x"2b1b09",x"2c1c09",x"241708",x"1d1208",x"191007",x"160f07",x"160f07",x"170f07",x"180f07",x"180f08",x"1a1108",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1d1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"341e0d",x"28160a",x"24150a",x"28170a",x"2e1a0b",x"301c0c",x"301c0c",x"341f0e",x"36200f",x"341e0d",x"2e1a0b",x"2f1b0c",x"27160a",x"2e1b0c",x"331d0e",x"321d0d",x"331e0d",x"37200d",x"38200e",x"321d0d",x"341f0d",x"432810",x"422710",x"442910",x"4c2d13",x"27170a",x"27170a",x"24150a",x"24150a",x"241509",x"26170b",x"24150a",x"231409",x"231409",x"221409",x"211309",x"201309",x"221409",x"201309",x"211409",x"211409",x"211409",x"201309",x"1f1208",x"1f1208",x"211309",x"221409",x"221409",x"231409",x"211309",x"231409",x"24150a",x"25160a",x"26170a",x"26160a",x"26160a",x"26160a",x"26160a",x"25150a",x"241509",x"241509",x"231409",x"231409",x"211309",x"1f1108",x"211309",x"231409",x"211309",x"201308",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"201309",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"211409",x"211409",x"211409",x"201309",x"201309",x"1f1309",x"1f1208",x"1f1208",x"1f1309",x"1e1208",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"191008",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"191007",x"191007",x"1a1007",x"000000"),
(x"150e07",x"150e07",x"150e07",x"26160a",x"412511",x"331d0d",x"25150a",x"472914",x"3d2311",x"3e2411",x"3a2110",x"422612",x"422611",x"452914",x"482a14",x"452913",x"412611",x"422612",x"432712",x"412511",x"371e0d",x"361d0d",x"381e0d",x"361d0d",x"391f0e",x"371e0d",x"3d220f",x"432612",x"442713",x"442813",x"462813",x"432612",x"462913",x"422611",x"412611",x"402510",x"422612",x"3b200e",x"371e0d",x"3a210f",x"432712",x"442813",x"3d2411",x"3f2410",x"3a1f0e",x"3a1f0d",x"402410",x"412410",x"3f2310",x"402410",x"422510",x"422511",x"3a200e",x"3f230f",x"3e220f",x"3d220f",x"3b210f",x"3b220f",x"432611",x"3e220f",x"3d220f",x"3f230f",x"381f0e",x"381f0d",x"3b200e",x"2f1b0c",x"3c210f",x"150e07",x"321c0d",x"150e07",x"301b0c",x"251509",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4b2b14",x"2b2219",x"372a1e",x"382a1f",x"3b2c1e",x"382819",x"362617",x"39281a",x"342517",x"302215",x"2f2114",x"312216",x"37281a",x"37281a",x"39281a",x"322316",x"342517",x"342517",x"332416",x"342516",x"352517",x"322316",x"322316",x"322416",x"332416",x"312214",x"302114",x"302114",x"322315",x"322316",x"332416",x"362618",x"312315",x"352517",x"312316",x"352618",x"342517",x"322316",x"322315",x"322316",x"322316",x"332417",x"322316",x"332517",x"342517",x"352618",x"322316",x"322316",x"2f2114",x"2f2116",x"322317",x"302216",x"342519",x"332417",x"342518",x"332518",x"36271a",x"302318",x"332519",x"342619",x"36281c",x"36281c",x"35281c",x"34281b",x"34261b",x"33261b",x"392a1c",x"3d2d1f",x"3a2c1f",x"3a2b1e",x"35271a",x"38291c",x"382a1d",x"38291d",x"332519",x"302318",x"302318",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1d0b",x"2f1d0b",x"341e0c",x"40260e",x"482b12",x"563417",x"28180b",x"2a190b",x"2f1c0b",x"27170a",x"2a190a",x"472a11",x"261809",x"1c1208",x"1d1208",x"1c1208",x"1d1308",x"1c1208",x"1c1208",x"191007",x"181007",x"181007",x"191007",x"170f07",x"160f07",x"170f07",x"181007",x"1b1107",x"190f07",x"1a1007",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1b1108",x"472a12",x"2f1e0a",x"291a09",x"281909",x"201408",x"231608",x"191007",x"1a1107",x"181007",x"180f07",x"180f08",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"1c1108",x"1c1108",x"1d1208",x"1d1208",x"1d1108",x"1c1108",x"1d1108",x"1d1208",x"1d1108",x"38200d",x"2f1b0b",x"281709",x"28170a",x"2f1c0d",x"301c0d",x"311d0c",x"35200e",x"321c0c",x"311d0c",x"1f1309",x"201409",x"29180b",x"28180b",x"28170b",x"29180b",x"27160a",x"321d0d",x"38220f",x"35200e",x"3a220f",x"39220e",x"41280f",x"3f2610",x"4c2d13",x"211409",x"241509",x"211308",x"211309",x"211309",x"211309",x"231509",x"24150a",x"24160a",x"23150a",x"221409",x"211409",x"201309",x"201309",x"201309",x"201409",x"1f1309",x"1e1208",x"201309",x"221409",x"23150a",x"23150a",x"23150a",x"221409",x"201208",x"211309",x"24150a",x"231509",x"241509",x"241509",x"25150a",x"25160a",x"231409",x"241509",x"241509",x"241509",x"24150a",x"241509",x"241509",x"221409",x"221409",x"211309",x"201308",x"1e1208",x"1f1208",x"211309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"201309",x"211409",x"201309",x"201309",x"211309",x"201309",x"201309",x"201308",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"1a1008",x"190f08",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"190f07",x"191007",x"1b1107",x"1c1108"),
(x"150e07",x"150e07",x"150e07",x"2d1a0c",x"3e2310",x"150e07",x"27160a",x"2e1a0b",x"3a210f",x"412411",x"412411",x"402310",x"3d210f",x"432611",x"442712",x"452712",x"462812",x"442712",x"462813",x"462712",x"3d210e",x"3d210f",x"381e0d",x"3b200e",x"3f2310",x"3f2410",x"412510",x"402310",x"3e230f",x"40230f",x"3f220f",x"3f230f",x"422510",x"3c210f",x"452712",x"3f2410",x"3a200e",x"39200e",x"3e2411",x"3f2511",x"3e2411",x"492a14",x"442813",x"432712",x"452812",x"3f230f",x"3c210f",x"3d210f",x"3f230f",x"40230f",x"3f230f",x"3f2310",x"482913",x"452812",x"462812",x"422510",x"3c210e",x"351d0c",x"391e0d",x"391f0d",x"3a200e",x"3e220e",x"3c200e",x"40230f",x"412510",x"432511",x"3a210f",x"2d190b",x"3b210e",x"150e07",x"321c0c",x"2e190a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"492a14",x"1e1711",x"3a2b1e",x"342519",x"3a291b",x"3a291a",x"3d2c1c",x"3d2b1c",x"3e2d1d",x"3d2c1c",x"422f20",x"3f2d1d",x"402f1f",x"402e1e",x"423120",x"402e1e",x"402e1e",x"443221",x"3e2c1c",x"3f2c1c",x"3e2c1b",x"3c2a1a",x"3c2b1b",x"3d2c1c",x"3b2a1b",x"412f1e",x"3f2d1c",x"412f1f",x"3d2c1d",x"3c2a1a",x"382617",x"3c2b1b",x"412f1e",x"3d2c1c",x"3d2c1c",x"3a291a",x"3f2d1d",x"3d2c1c",x"3e2d1d",x"3d2b1c",x"402e1e",x"402e1e",x"422f20",x"412f1e",x"402f1f",x"423020",x"402f1f",x"3e2d1d",x"402e1e",x"412f20",x"3a291a",x"3b2a1a",x"3c2a1a",x"3b2a1a",x"3f2d1d",x"3e2d1d",x"3d2c1d",x"3e2e1e",x"402e1f",x"3f2e1f",x"3e2d1f",x"362618",x"362618",x"3f2d1d",x"3e2d1f",x"3d2d1d",x"3e2d1e",x"3a2a1b",x"402e1f",x"3d2d1d",x"3c2c1d",x"3b2b1c",x"3c2b1c",x"3b2a1b",x"39291b",x"322417",x"322417",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"36200b",x"36200b",x"39220c",x"442910",x"503014",x"533116",x"29180a",x"2b1a0b",x"2e1c0b",x"2f1c0b",x"2a190a",x"41260f",x"1c1208",x"1d1308",x"1c1208",x"201408",x"1f1408",x"1a1107",x"1a1107",x"191007",x"180f07",x"1a1107",x"170f07",x"160e07",x"160e07",x"160f07",x"1a1107",x"170f07",x"1b1107",x"180f08",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"462a10",x"2f1d0a",x"2e1d0a",x"2d1c09",x"2a1b09",x"241608",x"1d1308",x"211508",x"1c1208",x"191007",x"1a1108",x"1a1008",x"1a1008",x"1c1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"1c1108",x"1c1108",x"251709",x"261709",x"231509",x"221509",x"1f1308",x"1b1108",x"1c1208",x"201409",x"241609",x"1e1309",x"231609",x"231509",x"201308",x"2a190b",x"231509",x"2b190b",x"301c0b",x"2d1a0b",x"301c0c",x"331f0c",x"3f250f",x"40260f",x"43290f",x"492c11",x"4a2c11",x"221408",x"231509",x"211409",x"231409",x"231509",x"231409",x"241509",x"221409",x"221408",x"211408",x"211408",x"201408",x"1f1208",x"211408",x"211309",x"1f1208",x"1f1208",x"201209",x"211509",x"211509",x"221509",x"231409",x"231509",x"231509",x"231409",x"221409",x"211309",x"221409",x"211309",x"221409",x"231409",x"231509",x"25160a",x"25150a",x"24150a",x"231409",x"211309",x"1f1208",x"1f1208",x"201208",x"201308",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"1f1209",x"201309",x"201309",x"201309",x"1f1208",x"211409",x"211409",x"211409",x"201409",x"1f1208",x"1f1208",x"1f1208",x"201309",x"1f1309",x"1f1309",x"1e1208",x"1d1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"170e07",x"180f07",x"1c1108",x"1c1108"),
(x"150e07",x"150e07",x"150e07",x"1a1008",x"38200f",x"311c0c",x"29170b",x"2c190b",x"2d1a0b",x"2f1b0c",x"2c190b",x"2c190b",x"2d190b",x"2c190b",x"2b180b",x"2f1b0c",x"2d1a0b",x"2d190b",x"2f1b0c",x"2e1a0b",x"2c190b",x"2e1a0b",x"29170a",x"251509",x"29170a",x"2d190b",x"2b180b",x"2a180a",x"2b180a",x"29170a",x"28160a",x"2b180a",x"2a170a",x"261509",x"28160a",x"28160a",x"271609",x"29170a",x"27170a",x"261509",x"241509",x"251509",x"29170a",x"29170a",x"2a180a",x"28170a",x"28170a",x"2c190b",x"2c180b",x"281609",x"2b180a",x"2c190b",x"2a180a",x"2d190b",x"2b180a",x"29170a",x"2a180a",x"27160a",x"2c190b",x"2a170a",x"251509",x"2d190b",x"211308",x"251509",x"251509",x"27160a",x"29170a",x"2e1a0b",x"39200e",x"150e07",x"3d220f",x"2b180a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"452611",x"150e07",x"332517",x"382719",x"3a2a1b",x"39281a",x"392819",x"392819",x"342416",x"3a2819",x"3b2a1b",x"3a291a",x"3d2b1b",x"3a2919",x"3d2c1c",x"3f2d1d",x"3c2a1b",x"3f2d1c",x"3a2919",x"392819",x"402e1d",x"3f2d1c",x"3e2b1b",x"3d2b1b",x"3e2c1c",x"3e2c1c",x"3d2b1c",x"392819",x"392819",x"392819",x"3a2819",x"3c2a1b",x"3b2a1b",x"3d2b1b",x"3d2b1c",x"402e1d",x"3f2e1e",x"3f2c1c",x"3e2c1c",x"3c2a1b",x"3b291a",x"3d2b1b",x"3d2c1c",x"3c2b1b",x"3e2c1c",x"3b2a1a",x"3f2d1c",x"402e1d",x"3d2b1b",x"3f2d1d",x"3a2919",x"372618",x"3e2c1c",x"3d2b1b",x"3a2919",x"3d2b1b",x"3b291a",x"3e2c1c",x"382719",x"332315",x"392819",x"362617",x"382718",x"3c2a1b",x"3d2b1c",x"3d2b1b",x"3a291a",x"3d2b1c",x"3c2b1c",x"3b2a1a",x"3a291a",x"392819",x"382718",x"372618",x"342517",x"2f2114",x"2f2114",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c240d",x"3c240d",x"3e250d",x"452810",x"43270f",x"462810",x"231508",x"28180a",x"25160a",x"28170a",x"27170a",x"3d230e",x"1a1107",x"231608",x"1b1108",x"1e1308",x"201408",x"1b1208",x"170f07",x"1b1108",x"191007",x"1f1408",x"1d1208",x"1c1108",x"160e07",x"160e07",x"160f07",x"191107",x"170f07",x"170f07",x"180f07",x"190f08",x"191008",x"191008",x"191008",x"190f08",x"190f08",x"452811",x"32200a",x"33200a",x"2f1e0a",x"301f0a",x"2b1b09",x"221508",x"241608",x"1e1408",x"1a1107",x"1a1007",x"180f07",x"191008",x"1b1108",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1b1108",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1b1108",x"251609",x"2d1c0a",x"271809",x"29190a",x"2b1a0a",x"201308",x"1e1308",x"1c1108",x"1d1208",x"221609",x"1e1208",x"241609",x"27180a",x"28170a",x"2a180b",x"2f1b0b",x"2e1b0b",x"2f1b0b",x"3b230d",x"39220d",x"3f260e",x"3e250d",x"442a0f",x"472a10",x"492b11",x"29190a",x"291909",x"241609",x"291909",x"271709",x"271809",x"221508",x"221509",x"261709",x"261709",x"251709",x"201409",x"211409",x"1e1308",x"211409",x"1e1208",x"1f1208",x"1e1208",x"211408",x"201408",x"1d1208",x"1e1208",x"1e1208",x"1e1208",x"1f1208",x"201309",x"201309",x"201208",x"1e1208",x"1f1208",x"211309",x"211309",x"201308",x"201308",x"201308",x"211309",x"201309",x"1f1308",x"1f1309",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1e1208",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1a1008",x"1a1008",x"191008",x"180f07",x"170f07",x"180f07",x"170f07",x"170f07",x"160e07",x"180f07",x"170f07",x"191007",x"180f07",x"1c1108"),
(x"150e07",x"150e07",x"150e07",x"211409",x"39200f",x"150e07",x"412511",x"432612",x"462712",x"462712",x"432511",x"472712",x"452712",x"4c2c15",x"4d2c14",x"492a13",x"4b2c15",x"4b2c15",x"4a2b14",x"4d2d15",x"4a2b14",x"492a14",x"462813",x"462712",x"452611",x"452711",x"452711",x"442611",x"452711",x"432511",x"3e220f",x"432511",x"442611",x"412410",x"432611",x"422511",x"3b200e",x"432611",x"412510",x"412510",x"412411",x"402410",x"412410",x"3e230f",x"3e220f",x"3b200e",x"422611",x"412410",x"40230f",x"432611",x"462812",x"462813",x"492a14",x"412410",x"432611",x"3b200e",x"341b0b",x"361d0c",x"371c0c",x"3b200e",x"3a1f0d",x"3d210e",x"3e230f",x"3d220f",x"3d220f",x"3a1f0d",x"361e0d",x"3e220f",x"39200e",x"150e07",x"3f2411",x"38200e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422511",x"150e07",x"382819",x"322416",x"362618",x"3a291a",x"3a291a",x"3b2a1b",x"382719",x"3c2a1b",x"3f2d1c",x"3d2b1b",x"3f2d1d",x"3d2b1b",x"3c2a1b",x"402d1d",x"3f2d1d",x"3d2b1c",x"3f2d1d",x"3d2b1b",x"402e1e",x"382718",x"3e2c1c",x"3e2c1c",x"412f1f",x"433120",x"3f2d1e",x"3f2d1d",x"402e1e",x"453220",x"3d2b1b",x"3f2d1d",x"3c2a1b",x"3e2c1d",x"3f2d1d",x"3e2c1c",x"3e2c1c",x"3f2d1c",x"3e2c1c",x"3d2b1c",x"3b291a",x"3d2b1b",x"3e2c1c",x"3d2b1b",x"422f1f",x"3e2c1c",x"3e2b1c",x"3e2c1d",x"412e1e",x"402d1d",x"3f2d1d",x"3a291a",x"3e2c1c",x"352516",x"3b2a1b",x"3f2d1d",x"3f2e1e",x"3f2e1e",x"3c2b1c",x"3c2a1b",x"3d2b1c",x"3d2c1d",x"3c2a1b",x"412f1e",x"3c2a1b",x"3d2b1c",x"3f2d1d",x"3b2a1b",x"3b291a",x"3f2d1c",x"3c2a1b",x"3a291a",x"362617",x"372718",x"3b291a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39220c",x"39220c",x"41270f",x"482a11",x"4b2c12",x"533114",x"261609",x"271709",x"221409",x"241509",x"26160a",x"412610",x"1d1308",x"221608",x"1f1408",x"1d1208",x"1f1408",x"1a1107",x"170f07",x"1e1308",x"241708",x"211508",x"160e07",x"1b1108",x"160e07",x"160e07",x"160e07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f08",x"180f07",x"180f07",x"180f07",x"4b2d10",x"37230b",x"36230b",x"33200a",x"35220b",x"2d1c0a",x"291a09",x"2a1a09",x"201508",x"1a1107",x"1a1107",x"180f07",x"191008",x"1b1108",x"1a1008",x"1a1008",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1008",x"1b1108",x"1b1108",x"1b1008",x"1b1008",x"2b1a0a",x"321f0b",x"261709",x"261709",x"261709",x"201408",x"201308",x"1f1308",x"1c1108",x"1b1108",x"261709",x"1d1108",x"25160a",x"321d0c",x"26160a",x"2d1b0b",x"36200d",x"38210e",x"3f260f",x"41270f",x"452a10",x"482c11",x"452a10",x"482c11",x"4f2f13",x"28180a",x"2b1b0a",x"2e1c0b",x"2c1b0b",x"311e0b",x"2a1a09",x"281909",x"281809",x"261709",x"241609",x"261709",x"241609",x"221509",x"221509",x"201408",x"251709",x"211409",x"221509",x"1e1208",x"201308",x"1e1308",x"201308",x"231609",x"1d1208",x"1e1208",x"1e1208",x"201309",x"1f1309",x"201309",x"221409",x"221409",x"231509",x"221409",x"211309",x"201309",x"1d1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"180f07",x"180f07",x"170f07",x"180f07",x"181007",x"180f07",x"180f07",x"191007",x"180f07",x"180f07",x"180f07",x"1a1107",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231509",x"38200e",x"150e07",x"371f0e",x"351e0d",x"3c220f",x"371f0e",x"3a210f",x"361e0d",x"371f0d",x"381e0d",x"381f0d",x"351e0d",x"3b210f",x"3a210f",x"381f0e",x"381f0d",x"381f0e",x"381f0e",x"3c210f",x"381f0d",x"361e0d",x"402511",x"3d2310",x"422611",x"3d2310",x"3c2310",x"3b2210",x"3a2210",x"3e2411",x"3b210f",x"351e0d",x"351e0d",x"321b0b",x"301a0b",x"311b0b",x"321c0c",x"341d0d",x"3a210f",x"3d2310",x"3a220f",x"3c2210",x"371f0e",x"39200e",x"3b210f",x"38200e",x"351e0d",x"381f0e",x"341c0d",x"301b0c",x"321c0c",x"351d0d",x"311b0c",x"2f1a0b",x"2e1a0b",x"361e0d",x"371f0d",x"371f0d",x"331d0c",x"331c0c",x"351e0d",x"371e0d",x"39200e",x"341d0d",x"381f0d",x"3e230f",x"150e07",x"3e230f",x"38200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422511",x"150e07",x"362618",x"3a281a",x"3d2c1c",x"3d2c1c",x"3a291a",x"3d2b1c",x"3c2a1b",x"412f1f",x"402e1e",x"3d2c1c",x"3f2d1d",x"453222",x"412f1f",x"443121",x"3f2e1e",x"3f2d1d",x"433020",x"44301f",x"402d1d",x"3c2a1a",x"3e2b1b",x"43301f",x"44301f",x"3f2d1d",x"3f2d1d",x"3f2d1d",x"402e1e",x"422f1e",x"3e2c1c",x"3f2d1c",x"3e2b1c",x"412f1e",x"3f2d1c",x"402d1d",x"433020",x"42301f",x"422f1e",x"412f1f",x"422f1f",x"443120",x"402e1e",x"3f2d1d",x"3f2d1d",x"473323",x"433120",x"453222",x"443121",x"423020",x"433020",x"3f2d1d",x"3e2b1c",x"3c2a1a",x"3a2919",x"402e1d",x"3f2d1d",x"3f2d1d",x"3d2b1c",x"3b2a1a",x"402e1e",x"3f2d1d",x"3d2b1b",x"3e2c1c",x"3d2a1b",x"3d2b1c",x"3c2a1b",x"402d1d",x"402e1e",x"3f2d1d",x"3c2b1b",x"3e2c1d",x"3c2a1b",x"3e2c1d",x"3b2a1b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412710",x"412710",x"43260e",x"45280f",x"482911",x"502f13",x"503014",x"27170a",x"26160a",x"28180b",x"251609",x"3e2310",x"221508",x"221608",x"191007",x"1e1308",x"1c1208",x"211508",x"170f07",x"1d1208",x"1c1208",x"251809",x"211508",x"180f07",x"180f07",x"170f07",x"160e07",x"160e07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"42270e",x"37230b",x"37230b",x"38230b",x"35210b",x"32200a",x"2a1a09",x"2b1b09",x"231608",x"1e1308",x"1c1107",x"180f07",x"191008",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"1b1108",x"2c1b0a",x"311e0a",x"2a1a09",x"2c1b0a",x"281909",x"231509",x"241609",x"221509",x"1c1108",x"1a1008",x"231509",x"231509",x"28170b",x"26160a",x"28170a",x"301c0b",x"301b0b",x"331d0c",x"39220d",x"42270e",x"42270e",x"43290e",x"462a0f",x"41270e",x"46290f",x"301d0a",x"2f1e0a",x"2c1b0a",x"301e0a",x"301d0a",x"2c1b0a",x"261709",x"281809",x"2f1d0a",x"271809",x"2a1a0a",x"241709",x"29190a",x"241609",x"281909",x"1c1108",x"1c1208",x"1e1309",x"201409",x"1f1308",x"1f1308",x"221509",x"1d1208",x"1d1208",x"1f1308",x"1e1208",x"1f1209",x"1f1209",x"1f1209",x"1e1208",x"1f1309",x"1e1208",x"1f1208",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1b1008",x"1b1008",x"1b1008",x"1b1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1008",x"1a1008",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"191008",x"190f07",x"190f07",x"180f07",x"170f07",x"170f07",x"171007",x"1a1007",x"1a1107",x"1b1107",x"1a1107",x"170f07",x"180f07",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"402511",x"331d0d",x"26160a",x"341d0d",x"331c0c",x"331c0d",x"2f1a0c",x"311b0c",x"341d0d",x"321c0c",x"341d0d",x"311c0c",x"311b0c",x"311b0c",x"301b0b",x"331c0c",x"2f1a0b",x"351d0d",x"341d0d",x"351d0d",x"371f0d",x"341d0d",x"341d0d",x"351d0d",x"371f0e",x"361e0e",x"361f0e",x"341e0d",x"361f0e",x"351d0d",x"311c0c",x"321c0c",x"301b0b",x"311c0d",x"301b0c",x"351e0d",x"331c0c",x"351d0d",x"321c0c",x"301a0b",x"331c0c",x"2e1a0b",x"331d0d",x"321c0d",x"321c0d",x"331c0d",x"311b0c",x"301b0c",x"2c190b",x"2e190b",x"311b0c",x"341c0c",x"2c180a",x"29160a",x"29160a",x"2e190b",x"361e0d",x"321c0c",x"301b0b",x"341d0d",x"301b0b",x"2a170a",x"29170a",x"2d180a",x"331c0c",x"150e07",x"311b0c",x"38200e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"452712",x"150e07",x"3c2b1c",x"412f1f",x"3d2c1d",x"3a291a",x"3c2a1b",x"3c2a1b",x"402d1d",x"402e1e",x"412f1f",x"443220",x"443120",x"412f1f",x"412f1e",x"3c2a1a",x"3c2a1a",x"3c2a1a",x"3b2a1a",x"3c2919",x"3b2919",x"3b2919",x"372617",x"3b2a19",x"3a2818",x"382718",x"3f2d1d",x"3e2b1c",x"3d2b1c",x"402d1d",x"433120",x"433120",x"412e1e",x"423020",x"463321",x"493624",x"42301f",x"422f1e",x"3f2d1c",x"3f2c1c",x"402d1d",x"402e1e",x"433120",x"443220",x"433120",x"412f1f",x"453220",x"3c2a1a",x"3d2b1b",x"3d2b1b",x"3a291a",x"3c2919",x"382717",x"352516",x"362516",x"3d2b1a",x"352416",x"3c2a1a",x"412f1e",x"3d2b1c",x"3f2c1c",x"3d2b1b",x"433120",x"433120",x"402d1d",x"412f1f",x"443120",x"443221",x"412f1f",x"3f2c1c",x"3e2c1c",x"392819",x"3d2b1b",x"3d2c1c",x"3e2d1d",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c240e",x"402510",x"472911",x"512e15",x"4b2c12",x"4f2e13",x"4a2b12",x"26160a",x"26160a",x"29180a",x"29180b",x"3f230f",x"241509",x"1f1408",x"1a1107",x"1b1108",x"160f07",x"191007",x"1e1308",x"160e07",x"160e07",x"231608",x"191007",x"160e07",x"1e1308",x"1b1107",x"180f07",x"160e07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"42260e",x"36220b",x"36220b",x"34210b",x"35220b",x"301e0a",x"291a09",x"2d1c09",x"221508",x"1c1208",x"1c1107",x"180f07",x"190f07",x"1b1007",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"2c1b0a",x"311d0a",x"301d0a",x"311d0b",x"2f1c0b",x"281709",x"231408",x"29180a",x"1f1308",x"27170a",x"27170a",x"2d1a0b",x"2f1a0c",x"231409",x"28170a",x"301b0b",x"311c0b",x"36200c",x"39220d",x"3c240d",x"462910",x"452a0f",x"45290f",x"44290e",x"43270e",x"2a1a0a",x"2b1a0a",x"2e1d0a",x"311f0b",x"311e0b",x"2e1d0a",x"2f1d0a",x"291a0a",x"271809",x"2a1a0a",x"2b1b0a",x"2a1a0a",x"281909",x"221508",x"261709",x"201408",x"241609",x"251709",x"1d1208",x"1b1108",x"1e1208",x"1d1208",x"201409",x"1c1108",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"1a1008",x"191008",x"190f07",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"190f07",x"190f07",x"190f07",x"180f07",x"191008",x"191008",x"1a1008",x"1a1008",x"190f07",x"190f07",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"190f08",x"190f07",x"180f07",x"170f07",x"170f07",x"170f07",x"160f07",x"191007",x"1b1107",x"1c1108",x"1e1308",x"1e1208",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"24150a",x"412611",x"351f0e",x"2b190b",x"402511",x"2a190b",x"3f2411",x"402511",x"452813",x"422612",x"402512",x"432611",x"412410",x"3f230f",x"3a200e",x"402310",x"432510",x"3f230f",x"412411",x"432611",x"442712",x"472914",x"442711",x"412511",x"412410",x"412410",x"3c210f",x"391f0e",x"3c210e",x"402310",x"3d220f",x"3a200e",x"3b200e",x"331b0b",x"361d0c",x"351c0c",x"3a1f0d",x"381e0d",x"381e0c",x"321b0b",x"361d0c",x"3b200d",x"3c200e",x"3c210e",x"381f0e",x"3b210e",x"3a200e",x"341c0b",x"341b0b",x"371d0d",x"3e2310",x"3f2410",x"412511",x"3a200f",x"371e0d",x"3b200f",x"422510",x"3f230f",x"3d210f",x"3b200e",x"3f2310",x"402410",x"150e07",x"3e220f",x"27160a",x"361e0d",x"150e07",x"3d220f",x"371f0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b1108",x"190f08",x"190f07",x"180f07",x"180f07",x"191008",x"190f07",x"190f07",x"190f07",x"190f07",x"180f07",x"191007",x"170f07",x"180f08",x"1b1008",x"170f07",x"150e07",x"170f07",x"180f07",x"190f07",x"191008",x"190f07",x"191008",x"180f07",x"170f07",x"160e07",x"160e07",x"170f07",x"160f07",x"170f07",x"180f07",x"1a1008",x"191008",x"180f07",x"1a1008",x"191008",x"191008",x"1a1008",x"170f07",x"191008",x"1a1008",x"170f07",x"150e07",x"190f07",x"180f07",x"180f07",x"170f07",x"191008",x"160e07",x"190f07",x"170f07",x"180f07",x"190f07",x"170f07",x"150e07",x"170f07",x"180f07",x"1a1107",x"1b1108",x"1e1308",x"201409",x"231609",x"231608",x"281909",x"2b1b09",x"261808",x"201508",x"191007",x"150e07",x"170f07",x"180f07",x"180f07",x"190f07",x"180f07",x"180f07",x"180f07",x"180f07",x"190f08",x"181007",x"180f08",x"180f08",x"160e07",x"190f08",x"180f08",x"180f08",x"180f07",x"191007",x"170f07",x"170f07",x"160f07",x"170f07",x"180f08",x"160e07",x"160f07",x"160e07",x"170f07",x"160e07",x"150e07",x"190f08",x"170f07",x"1a1008",x"191007",x"1a1008",x"1b1108",x"1a1008",x"180f08",x"180f08",x"191008",x"180f07",x"170f07",x"211308",x"2a170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"462812",x"22180e",x"523c29",x"523c28",x"4d3825",x"4f3926",x"513b28",x"523c28",x"4f3a26",x"533d29",x"563f2a",x"543d29",x"533d29",x"513b28",x"533d29",x"4b3623",x"4c3622",x"4d3723",x"483320",x"473220",x"493320",x"4f3824",x"4e3723",x"513a25",x"4f3825",x"503925",x"4f3927",x"4e3825",x"513b28",x"513b27",x"523c28",x"543d29",x"553e2a",x"58412b",x"59422d",x"5d452f",x"583f2b",x"543d29",x"513b28",x"553e29",x"563e29",x"543e29",x"533d29",x"563f2a",x"573f2b",x"533c28",x"533d29",x"4a3422",x"4f3824",x"4f3924",x"493320",x"473220",x"483320",x"4c3622",x"4c3522",x"4d3723",x"4d3724",x"4f3825",x"513b28",x"513b28",x"523c28",x"4f3a25",x"4f3926",x"533c28",x"4f3927",x"533d29",x"56402b",x"4f3a27",x"503a26",x"533c28",x"523c28",x"503a27",x"4e3925",x"503b27",x"523c28",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442710",x"42260f",x"371f0b",x"45260f",x"44260e",x"492b12",x"492b12",x"311d0b",x"261709",x"301c0b",x"40240e",x"1f1308",x"1d1308",x"1d1308",x"1c1208",x"1d1308",x"42250f",x"311d0b",x"27170a",x"211409",x"1f1309",x"1f1309",x"181007",x"1a1008",x"1d130b",x"321e11",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"170f07",x"190f07",x"1b1008",x"1d1108",x"1d1208",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1108",x"1f1208",x"211409",x"241609",x"1c1108",x"422711",x"482c12",x"452a11",x"1d1209",x"1e1309",x"1d1208",x"1b1008",x"1c1108",x"1b1108",x"1a1008",x"261709",x"2c1b0a",x"2b1b0a",x"35210b",x"492b10",x"43280e",x"1e1308",x"1d1208",x"190f08",x"1c1108",x"1b1107",x"1c1208",x"1d1208",x"170f07",x"191007",x"1f1308",x"201408",x"291909",x"2d1c0a",x"311e0a",x"38220b",x"40270e",x"3c250d",x"3f260d",x"41260e",x"271709",x"37230b",x"37230b",x"301e0a",x"2e1c0a",x"2d1c0a",x"2f1d0b",x"281909",x"251708",x"281909",x"2a1b09",x"271909",x"261809",x"231608",x"2a1b09",x"1e1308",x"1b1107",x"221508",x"201408",x"281909",x"261808",x"1d1208",x"170f07",x"170f07",x"180f07",x"190f07",x"191008",x"191008",x"1a1008",x"191008",x"180f07",x"190f07",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"190f08",x"180f07",x"180f08",x"180f07",x"180f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"180f07",x"170f07",x"1a1007",x"1c1108",x"1a1107",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231509",x"412410",x"150e07",x"1d1208",x"3f230f",x"351c0c",x"381d0c",x"311b0c",x"341e0d",x"361f0e",x"39200f",x"371f0e",x"371f0e",x"39200e",x"371f0d",x"341d0c",x"341d0c",x"341d0d",x"361e0d",x"371f0e",x"341d0d",x"341d0d",x"341d0d",x"331c0d",x"331d0d",x"321c0d",x"321c0d",x"341d0d",x"351e0e",x"351e0d",x"361f0e",x"351e0d",x"331d0d",x"2f1a0b",x"311b0c",x"311b0c",x"321c0c",x"301a0b",x"321c0c",x"321c0c",x"321c0c",x"341c0c",x"341c0c",x"311b0c",x"2d190b",x"331c0c",x"351d0d",x"2f1a0b",x"2f1a0b",x"2e1a0b",x"301a0b",x"301a0b",x"301b0c",x"311b0c",x"321c0c",x"311b0b",x"331c0c",x"341d0c",x"371e0d",x"371f0d",x"311a0b",x"3f230f",x"3f240f",x"472812",x"2a180b",x"422511",x"150e07",x"422611",x"361e0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351e0d",x"351e0d",x"1b1108",x"190f08",x"190f07",x"180f07",x"180f07",x"191008",x"190f07",x"190f07",x"190f07",x"190f07",x"180f07",x"191007",x"170f07",x"180f08",x"1b1008",x"170f07",x"150e07",x"170f07",x"180f07",x"190f07",x"191008",x"190f07",x"191008",x"180f07",x"170f07",x"160e07",x"160e07",x"170f07",x"160f07",x"170f07",x"180f07",x"1a1008",x"191008",x"180f07",x"1a1008",x"191008",x"191008",x"1a1008",x"170f07",x"191008",x"1a1008",x"170f07",x"150e07",x"190f07",x"180f07",x"180f07",x"170f07",x"191008",x"160e07",x"190f07",x"170f07",x"180f07",x"190f07",x"170f07",x"150e07",x"170f07",x"180f07",x"1a1107",x"1b1108",x"1e1308",x"201409",x"231609",x"231608",x"281909",x"2b1b09",x"261808",x"201508",x"191007",x"150e07",x"170f07",x"180f07",x"180f07",x"190f07",x"180f07",x"180f07",x"180f07",x"180f07",x"190f08",x"181007",x"180f08",x"180f08",x"160e07",x"190f08",x"180f08",x"180f08",x"180f07",x"191007",x"170f07",x"170f07",x"160f07",x"170f07",x"180f08",x"160e07",x"160f07",x"160e07",x"170f07",x"160e07",x"150e07",x"190f08",x"170f07",x"1a1008",x"191007",x"1a1008",x"1b1108",x"1a1008",x"180f08",x"180f08",x"191008",x"180f07",x"170f07",x"211308",x"2a170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4b2b14",x"1d1208",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"371f0b",x"3d210d",x"3d230f",x"492911",x"512f15",x"3e240e",x"39200d",x"2a1a0a",x"371f0d",x"2c190b",x"2c190b",x"1d1308",x"47280f",x"482910",x"45260f",x"301c0b",x"2b1a0a",x"201308",x"211408",x"1e1208",x"1e1208",x"1e1208",x"1d120b",x"1d120a",x"2c1b0f",x"2c1b0f",x"160e07",x"160e07",x"170f07",x"1c1108",x"1a1008",x"1c1108",x"211409",x"201309",x"1c1108",x"1c1108",x"1e1108",x"1f1208",x"221309",x"221309",x"29170a",x"201308",x"26160a",x"211309",x"1e1208",x"1e1208",x"1e1108",x"1f1208",x"211409",x"241509",x"2c1a0b",x"3f2710",x"422812",x"472b12",x"3e2613",x"392516",x"352113",x"1b1008",x"1c1108",x"1b1108",x"1a1008",x"261709",x"38240b",x"37230b",x"34200a",x"301e0a",x"41270e",x"42280e",x"462712",x"29180a",x"2b180b",x"28170a",x"25150a",x"25160a",x"25150a",x"180f07",x"180f07",x"180f07",x"29180b",x"251509",x"28170a",x"26160a",x"241509",x"231509",x"211408",x"39210d",x"41250f",x"492c11",x"462910",x"4a2c11",x"46290f",x"482a11",x"452810",x"44270f",x"452810",x"452810",x"43270f",x"452710",x"482911",x"472911",x"432610",x"41250f",x"41250f",x"442710",x"3e230e",x"3f240f",x"3f240f",x"402510",x"452711",x"41250f",x"3c200e",x"3c210e",x"381f0d",x"3c210e",x"3b210e",x"3b220f",x"3e230f",x"3d210e",x"3a1f0d",x"391f0d",x"3a1f0d",x"371e0c",x"3d220f",x"3c210f",x"3b200e",x"3d220e",x"3d210f",x"3d220f",x"3c210e",x"3b200d",x"3b200d",x"3c210e",x"3a200e",x"3d220f",x"3f230f",x"3e230f",x"3f2310",x"3b210f",x"3d220f",x"3d220f",x"3c210f",x"3e220f",x"381f0d",x"3c220e",x"381f0d",x"3e220f",x"3d220f",x"3d220f",x"402410",x"452611",x"432611",x"412410",x"3e2310",x"432611",x"3d220f",x"3b210f",x"351d0d",x"160e07",x"1b1107",x"1a1107",x"1e1208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"26160a",x"3c210e",x"150e07",x"1d1108",x"211308",x"221409",x"251509",x"331c0c",x"3a210f",x"3b210f",x"3b200e",x"381f0e",x"3a200e",x"3f2410",x"402410",x"432611",x"3d220f",x"3e2310",x"3f2410",x"3f2310",x"3e220f",x"3b210f",x"3b210f",x"3b210e",x"3d220f",x"3d220f",x"3b210f",x"3c210f",x"371f0d",x"3b210f",x"3b210f",x"361e0d",x"351d0d",x"311b0b",x"351d0c",x"381f0d",x"361e0d",x"381f0d",x"3c210f",x"371e0d",x"361d0c",x"381f0d",x"381f0d",x"3b200e",x"321c0c",x"3a200e",x"3b210f",x"402410",x"3d220f",x"3d220f",x"3c210f",x"39200e",x"3a200e",x"381f0e",x"3c220f",x"3e2310",x"3e230f",x"3c220f",x"3f2310",x"3f230f",x"3b210f",x"482913",x"150e07",x"28170a",x"2c1a0b",x"301c0d",x"2b190b",x"3e2310",x"38200e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c220f",x"3c220f",x"2d190b",x"26150a",x"261509",x"231409",x"211309",x"26160a",x"251509",x"271509",x"251509",x"251509",x"211309",x"251509",x"1f1208",x"231409",x"231409",x"1e1108",x"170f07",x"1f1208",x"231409",x"241409",x"26160a",x"251509",x"27160a",x"211309",x"1e1208",x"1b1008",x"1a1008",x"1d1108",x"1c1108",x"1e1108",x"231509",x"29170a",x"27160a",x"221409",x"27160a",x"241509",x"241509",x"221409",x"1f1208",x"24150a",x"27160a",x"1f1209",x"150e07",x"241509",x"221409",x"241509",x"201309",x"26160a",x"1a1008",x"251509",x"1e1208",x"221409",x"241509",x"1e1208",x"150e07",x"1d1108",x"1c1008",x"1f1208",x"1e1208",x"221609",x"26160a",x"29190a",x"261709",x"2d1b0a",x"261809",x"2e1c0a",x"251709",x"1e1208",x"150e07",x"1f1208",x"231409",x"231509",x"251509",x"221409",x"211309",x"221409",x"211409",x"24150a",x"231509",x"201309",x"221409",x"180f07",x"1d1108",x"211409",x"211409",x"221409",x"241509",x"201309",x"1e1208",x"1b1108",x"201309",x"24150a",x"180f07",x"1c1108",x"180f07",x"1d1108",x"180f08",x"150e07",x"25150a",x"1f1309",x"28170a",x"241509",x"28170a",x"2c190b",x"271509",x"201309",x"231409",x"26160a",x"201308",x"1b1008",x"211308",x"29160a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"482912",x"482912",x"150e07",x"150e07",x"160e07",x"1c1008",x"1d1108",x"221309",x"241409",x"231409",x"211308",x"241409",x"241509",x"29170b",x"29180b",x"2c190b",x"2e1b0c",x"2f1b0d",x"2a190b",x"221409",x"27170a",x"251509",x"26160a",x"2d190b",x"2e1a0c",x"2c1a0b",x"2d1a0c",x"2e1a0c",x"2b190b",x"2b180a",x"2d190b",x"2b190b",x"27160a",x"28170a",x"2c190b",x"2e1a0b",x"2a170a",x"2a170a",x"27160a",x"221409",x"241409",x"221409",x"231409",x"28160a",x"241509",x"261509",x"231409",x"29170a",x"2e190b",x"2d190a",x"2c180b",x"2d190b",x"2f1a0b",x"301b0b",x"311b0c",x"301b0c",x"2d190b",x"2a170a",x"2e1a0b",x"301b0c",x"311b0c",x"341d0d",x"311c0d",x"311c0c",x"341d0d",x"321c0d",x"311c0d",x"321d0e",x"351f0f",x"331e0e",x"311c0d",x"2d1a0c",x"331d0d",x"331d0d",x"2d190b",x"2d190b",x"2e1a0b",x"2e1b0b",x"2a180b",x"26160a",x"1e1208",x"1b1108",x"1f1208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1007",x"1a1007",x"1b1107",x"4f2f15",x"543115",x"3b230e",x"37200d",x"2b1a0a",x"3a220e",x"38210e",x"000000",x"4d2c13",x"4b2b12",x"47280f",x"351f0d",x"2d1b0a",x"241609",x"251609",x"231509",x"1f1208",x"1f1309",x"1d1208",x"1f130b",x"1e130b",x"2c1b0f",x"2c1b0f",x"000000",x"000000",x"211509",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1f1209",x"1e1208",x"1c1108",x"1d1208",x"1f1309",x"1e1208",x"1f1309",x"201309",x"1f1309",x"1f1309",x"201309",x"201309",x"221409",x"26170a",x"211308",x"2b1a0a",x"28180b",x"402711",x"412710",x"3b240d",x"3c2616",x"352113",x"2f1e0f",x"2d1e13",x"000000",x"000000",x"000000",x"35220b",x"36220b",x"39240b",x"36220b",x"39240b",x"33200a",x"41270e",x"462712",x"29180a",x"2b180b",x"28170a",x"25150a",x"25160a",x"25150a",x"180f07",x"180f07",x"180f07",x"29180b",x"251509",x"28170a",x"26160a",x"241509",x"231509",x"211408",x"2a190a",x"29180a",x"241509",x"2a180a",x"221509",x"1b1008",x"1d1208",x"26160a",x"24150a",x"28170b",x"2c1a0b",x"2d190b",x"28170a",x"2c190b",x"311b0c",x"341d0d",x"40250e",x"231608",x"1d1208",x"3b210e",x"462711",x"40240f",x"3c210e",x"351d0c",x"351d0c",x"3a200e",x"40230f",x"3e220f",x"3f230f",x"3f230f",x"402410",x"422510",x"432511",x"422510",x"412410",x"3f230f",x"3a200e",x"3c210f",x"3c220f",x"3a210f",x"3a210f",x"3a220f",x"351e0d",x"361e0d",x"38200e",x"38200f",x"3a210f",x"39200e",x"37200e",x"38200f",x"2b190b",x"512e14",x"4d2d15",x"452711",x"482911",x"492a12",x"442711",x"4b2b14",x"482912",x"432611",x"412410",x"40230f",x"40230f",x"432611",x"3f230f",x"3c210f",x"3b200d",x"3d220f",x"3e230f",x"3d220f",x"341d0d",x"381e0d",x"160e07",x"1d1208",x"1b1107",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"3b210e",x"150e07",x"281609",x"341d0d",x"341e0d",x"321d0d",x"371f0e",x"38200e",x"38200e",x"3b220f",x"3b210f",x"3d2310",x"3d2310",x"38200f",x"39200f",x"3b210f",x"3f2410",x"3b220f",x"381f0e",x"321c0c",x"361e0d",x"3c220f",x"3b210f",x"351e0e",x"331d0d",x"381f0e",x"351d0d",x"321b0c",x"311b0b",x"341c0c",x"331c0c",x"321b0c",x"321b0c",x"331c0c",x"331c0c",x"311b0b",x"371e0d",x"341c0c",x"361d0c",x"311b0b",x"321b0b",x"371e0d",x"391f0e",x"341d0d",x"3b210f",x"3c220f",x"3a210f",x"351d0d",x"331c0c",x"371e0d",x"331c0c",x"331c0c",x"331d0d",x"381f0e",x"371f0e",x"351e0e",x"351d0d",x"3b210f",x"3d220f",x"3e2310",x"4a2a14",x"211409",x"38200f",x"3b210f",x"3c220f",x"321c0c",x"3f2410",x"39200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381c0c",x"381c0c",x"28170a",x"29170a",x"231409",x"2a180a",x"25160a",x"26160a",x"2a180a",x"27160a",x"201309",x"241509",x"221409",x"26160a",x"231409",x"29170a",x"201308",x"1c1108",x"1b1108",x"1b1108",x"231409",x"231409",x"251509",x"241509",x"211309",x"231409",x"221309",x"221308",x"241509",x"25150a",x"1a1008",x"231509",x"1f1309",x"241509",x"26160a",x"2a180b",x"24150a",x"27170b",x"25150a",x"231509",x"27160a",x"241509",x"1e1208",x"1d1108",x"1c1108",x"1d1108",x"201309",x"27170a",x"201309",x"241509",x"1f1309",x"1e1208",x"231409",x"201308",x"211309",x"211309",x"231409",x"1d1108",x"221409",x"211309",x"1a1008",x"1e1208",x"1d1108",x"241509",x"201308",x"1b1107",x"221409",x"231509",x"1f1208",x"231509",x"1f1309",x"241509",x"25150a",x"25150a",x"26160a",x"180f07",x"251509",x"261609",x"221409",x"26150a",x"211409",x"231509",x"261609",x"25160a",x"28170a",x"201309",x"221409",x"231509",x"1e1209",x"1d1208",x"1d1108",x"241509",x"1e1108",x"180f07",x"201208",x"201309",x"1d1208",x"190f08",x"1d1208",x"231409",x"201208",x"201308",x"251509",x"27160a",x"261509",x"27160a",x"221409",x"241509",x"27160a",x"25160a",x"231409",x"231409",x"1e1208",x"241509",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442611",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1008",x"1d1108",x"221309",x"241409",x"231409",x"211308",x"241409",x"241509",x"29170b",x"29180b",x"2c190b",x"2e1b0c",x"2f1b0d",x"2a190b",x"221409",x"27170a",x"251509",x"26160a",x"2d190b",x"2e1a0c",x"2c1a0b",x"2d1a0c",x"2e1a0c",x"2b190b",x"2b180a",x"2d190b",x"2b190b",x"27160a",x"28170a",x"2c190b",x"2e1a0b",x"2a170a",x"2a170a",x"27160a",x"221409",x"241409",x"221409",x"231409",x"28160a",x"241509",x"261509",x"231409",x"29170a",x"2e190b",x"2d190a",x"2c180b",x"2d190b",x"2f1a0b",x"301b0b",x"311b0c",x"301b0c",x"2d190b",x"2a170a",x"2e1a0b",x"301b0c",x"311b0c",x"341d0d",x"311c0d",x"311c0c",x"341d0d",x"321c0d",x"311c0d",x"321d0e",x"351f0f",x"331e0e",x"311c0d",x"2d1a0c",x"331d0d",x"331d0d",x"2d190b",x"2d190b",x"2e1a0b",x"2e1b0b",x"2a180b",x"26160a",x"1e1208",x"241509",x"251509",x"241409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1007",x"1a1007",x"1b1107",x"211508",x"1e1308",x"241708",x"231608",x"4b2910",x"39210d",x"3b220d",x"522f15",x"43260f",x"4e2d14",x"331f0c",x"301e0b",x"2d1c0a",x"281809",x"231609",x"1e1108",x"1f1209",x"1e1208",x"1e1208",x"1f140a",x"1f130b",x"21170f",x"21170f",x"000000",x"000000",x"1c1108",x"241609",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1c1108",x"1d1108",x"1e1108",x"201309",x"201309",x"201309",x"201309",x"1f1208",x"1d1108",x"1d1108",x"201308",x"211309",x"1f1208",x"241509",x"27170a",x"26170a",x"25150a",x"3e2512",x"3b220f",x"2f1c0d",x"312012",x"2f1d0d",x"332114",x"2a1f17",x"2a221a",x"241c15",x"311e0a",x"311f0a",x"35220b",x"37230b",x"3a250b",x"3c260c",x"34210b",x"34210b",x"452910",x"3a200e",x"2d180a",x"251409",x"2b180b",x"2b190b",x"2b190b",x"28170a",x"201309",x"170f07",x"3f2410",x"402511",x"422611",x"3f2411",x"3e2410",x"402410",x"3f240f",x"432610",x"3d230f",x"3f2410",x"3c200f",x"3c210f",x"3b220f",x"351e0e",x"3e2310",x"3c2310",x"3c220f",x"3b200e",x"391f0d",x"3a1f0d",x"41240f",x"3e220f",x"3a200d",x"1d1308",x"251809",x"221508",x"1d1208",x"442611",x"40230f",x"341c0c",x"341c0c",x"391e0d",x"351d0c",x"391f0d",x"3e220f",x"3d220f",x"3e2310",x"3e2310",x"3d220f",x"3b210f",x"3a200e",x"371f0d",x"391f0d",x"3c210e",x"3b210f",x"3f2310",x"3e2310",x"3c220f",x"3e230f",x"3b200e",x"3e230f",x"3f2310",x"412511",x"402511",x"3f2511",x"3f2310",x"3c210f",x"2c190b",x"4c2c13",x"3c210e",x"381f0c",x"3d230f",x"3c2310",x"3e2310",x"3c210f",x"3b230e",x"311b0b",x"2b180a",x"331c0b",x"361e0d",x"361e0d",x"331c0d",x"351d0d",x"331d0d",x"301b0c",x"2f1b0c",x"311c0c",x"2e1a0b",x"2b180b",x"28170a",x"25160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231509",x"412511",x"150e07",x"2f1b0c",x"361f0e",x"351e0d",x"2c180b",x"251509",x"3e220f",x"412310",x"3f230f",x"442611",x"3f2310",x"3f230f",x"422511",x"40230f",x"462711",x"4a2b14",x"492a14",x"472913",x"452812",x"462712",x"432611",x"412410",x"3b210e",x"432510",x"462711",x"432511",x"452712",x"462812",x"422510",x"3f230f",x"3d220e",x"3c210e",x"3f230f",x"3c210e",x"3d210e",x"3b200d",x"3f220e",x"3f220e",x"3f220e",x"3a1f0d",x"3f220f",x"42240f",x"3b200e",x"41230f",x"3d210e",x"412410",x"3a200e",x"3c210e",x"3a1e0d",x"3d210e",x"3c220f",x"3f2410",x"412511",x"3f2411",x"442712",x"4c2d16",x"482a14",x"4a2b15",x"533117",x"150e07",x"2f1b0c",x"39210f",x"38200f",x"3a210f",x"311b0c",x"3e2310",x"38210f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2912",x"4a2912",x"2d190b",x"271609",x"231409",x"231409",x"231509",x"231509",x"2b190b",x"2f1b0c",x"2e1b0c",x"2c1a0b",x"2d1a0b",x"2a180b",x"2a180b",x"28170a",x"29170a",x"251509",x"201309",x"26160a",x"27160a",x"26160a",x"27160a",x"231409",x"26160a",x"231409",x"251509",x"28170a",x"2b190b",x"2b190b",x"211309",x"271609",x"29170a",x"2c190b",x"2a180b",x"28160a",x"29180a",x"26160a",x"25150a",x"28170a",x"25150a",x"27170a",x"25150a",x"1e1208",x"241509",x"201309",x"241509",x"1d1108",x"2a180a",x"2a180b",x"231409",x"1c1108",x"241509",x"27160a",x"201309",x"1f1208",x"241409",x"281609",x"271609",x"241509",x"201409",x"271609",x"2a1809",x"241609",x"1f1308",x"251609",x"2a180a",x"28180a",x"26160a",x"231509",x"251609",x"231509",x"261609",x"251609",x"241609",x"251508",x"28170a",x"28170a",x"26160a",x"2c1a0b",x"2f1b0c",x"25160a",x"27170a",x"2c1a0b",x"29190b",x"28180a",x"29180b",x"25160a",x"27170b",x"1d1108",x"26160a",x"241509",x"211308",x"201208",x"1a1008",x"1c1108",x"231409",x"211309",x"1c1108",x"231409",x"211308",x"261609",x"211308",x"281609",x"221308",x"251509",x"27160a",x"29170a",x"29170a",x"2b190b",x"2b190b",x"28170b",x"231509",x"27170a",x"23150a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422510",x"472811",x"452711",x"221409",x"211309",x"2a170a",x"301b0c",x"311c0c",x"2d190b",x"2f1a0b",x"2f1b0c",x"2d1a0b",x"2e1a0b",x"2b180b",x"2c190b",x"2f1b0c",x"301b0c",x"311b0c",x"311b0c",x"321c0c",x"2d190b",x"321c0d",x"321c0c",x"361e0d",x"371f0e",x"341e0e",x"341e0d",x"38200e",x"361f0e",x"341d0d",x"351d0d",x"2f1a0b",x"2f1b0c",x"2f1a0c",x"331d0d",x"311c0d",x"331d0d",x"301b0c",x"2c190b",x"2d190b",x"2e190b",x"2c190b",x"2d190a",x"2b180a",x"2e190a",x"2b180a",x"2e1a0a",x"2e190a",x"321c0b",x"311c0b",x"2f1a0b",x"2e1a0b",x"311b0b",x"311b0c",x"321c0c",x"341d0c",x"2e190b",x"2a170a",x"2d190b",x"321c0c",x"331d0d",x"361f0f",x"37200f",x"341d0e",x"351f0f",x"36200f",x"321d0d",x"37200f",x"341e0e",x"341e0e",x"37200e",x"341e0e",x"2d190b",x"2c190b",x"2d190b",x"2a170a",x"291609",x"291509",x"2b180a",x"301b0c",x"381f0e",x"3a1f0c",x"553319",x"5c381c",x"5c381c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"190f07",x"191007",x"191007",x"1f1308",x"211408",x"201408",x"231608",x"38200c",x"3c230d",x"3a220d",x"533015",x"512e14",x"37200c",x"2d1b0b",x"311e0a",x"2c1b0a",x"311d0a",x"231509",x"1d1108",x"1f1309",x"1f1209",x"201309",x"1f1309",x"20140b",x"20140c",x"2e1c10",x"2e1c10",x"000000",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1b1008",x"1c1008",x"1c1108",x"1f1208",x"1e1208",x"1f1208",x"201208",x"1e1208",x"201308",x"1e1208",x"231508",x"231508",x"231509",x"27170a",x"27170a",x"28170a",x"3b2312",x"321d0e",x"2a1a0c",x"2d1c0f",x"291a0e",x"251c14",x"33261c",x"292019",x"231b13",x"281809",x"2d1c0a",x"2f1e0a",x"37230b",x"35210b",x"38230b",x"35210b",x"32200a",x"291a09",x"2c190b",x"2d190b",x"241509",x"27170a",x"29180b",x"1f1208",x"170f07",x"191008",x"170f07",x"361f0e",x"381f0e",x"39200e",x"381f0d",x"351d0d",x"3f230f",x"371f0d",x"3e220f",x"402411",x"38200e",x"3b220f",x"3c220f",x"3b210f",x"2b180b",x"351d0d",x"371e0e",x"381f0e",x"331c0c",x"3a210f",x"402411",x"522f16",x"3b220d",x"211508",x"1a1107",x"181007",x"160f07",x"191007",x"201408",x"422511",x"3d210e",x"381e0c",x"361d0c",x"361d0c",x"381f0d",x"371e0d",x"311b0b",x"351d0d",x"371e0d",x"371e0d",x"381e0d",x"361d0d",x"361d0c",x"3b210e",x"3f2410",x"412611",x"402511",x"412512",x"3f2411",x"412612",x"422612",x"442813",x"452813",x"422612",x"422512",x"452813",x"402411",x"2d190b",x"2f1a0c",x"442610",x"301a0a",x"341d0b",x"2f190a",x"38200d",x"3c220f",x"3a210e",x"381f0d",x"281609",x"311b0b",x"321b0b",x"2f1a0b",x"2e1a0b",x"331c0c",x"351d0d",x"321d0d",x"311b0c",x"351e0d",x"311c0c",x"351e0e",x"2b190b",x"1d1208",x"150e07",x"25150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"442813",x"150e07",x"28170a",x"321c0c",x"331d0d",x"2e1a0b",x"311c0c",x"381f0e",x"3a200e",x"351d0d",x"331d0d",x"331d0d",x"39200f",x"341d0d",x"2e1a0c",x"341d0d",x"361f0e",x"37200f",x"2d1a0b",x"311c0c",x"321c0d",x"301b0c",x"321c0c",x"2e1a0b",x"321c0c",x"341d0d",x"341e0d",x"2f1b0c",x"311c0c",x"2e1a0b",x"2b170a",x"2c180a",x"2c180a",x"2f1a0b",x"351d0d",x"321c0c",x"311c0c",x"2f1b0b",x"29160a",x"2b180a",x"29170a",x"301b0b",x"2a180a",x"2c180b",x"2d190b",x"28160a",x"2d190b",x"301b0c",x"301b0c",x"27160a",x"27160a",x"29170a",x"2e1a0b",x"361f0e",x"361f0e",x"331d0d",x"361f0e",x"3c2310",x"402511",x"422612",x"27170b",x"2a180b",x"361f0e",x"39200f",x"361f0e",x"301c0c",x"3f2411",x"371f0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29170a",x"29170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1107",x"191007",x"1a1107",x"1c1208",x"1b1108",x"1d1308",x"1c1208",x"1c1208",x"1f1408",x"201508",x"201508",x"201508",x"1f1408",x"201508",x"1e1308",x"1f1408",x"1c1208",x"1c1208",x"181007",x"1a1107",x"1b1108",x"1c1208",x"181007",x"181007",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"a8a8a8",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"492912",x"472811",x"3e220f",x"371e0d",x"3e210e",x"452611",x"482811",x"3d210e",x"3c210e",x"3b200e",x"3e220e",x"3d210e",x"3f230f",x"3c210e",x"3f230f",x"402410",x"432611",x"492a14",x"482b14",x"492a15",x"4a2b15",x"4b2c15",x"492a14",x"472813",x"462812",x"4a2b14",x"4a2a14",x"492a14",x"4a2b14",x"4b2c15",x"492a14",x"482913",x"452812",x"442611",x"462812",x"492a14",x"452813",x"412410",x"442711",x"412410",x"422611",x"452812",x"442711",x"442711",x"422611",x"442712",x"452812",x"452711",x"452812",x"422510",x"412410",x"432611",x"442711",x"422611",x"442712",x"452712",x"462813",x"492a14",x"452712",x"442612",x"412410",x"40230f",x"3f230f",x"442611",x"422511",x"412410",x"412410",x"40230f",x"3f230f",x"402410",x"442712",x"432611",x"432611",x"432611",x"412511",x"442712",x"452812",x"432712",x"452712",x"472913",x"492914",x"482a14",x"57341a",x"5c381c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"191007",x"1d1308",x"1e1308",x"211608",x"1f1408",x"251709",x"28180a",x"452810",x"3f250e",x"4c2a11",x"513015",x"371f0c",x"35200b",x"2a1a0a",x"2c1b0a",x"2f1d0b",x"2b1b0a",x"1e1208",x"1f1209",x"1d1108",x"1f1309",x"201309",x"1f1309",x"1e1209",x"20140b",x"291a10",x"291a10",x"000000",x"1b1108",x"1a1008",x"1e1208",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1f1208",x"1f1209",x"1f1208",x"1e1208",x"201309",x"1f1208",x"1e1208",x"201308",x"1d1108",x"221409",x"231409",x"231509",x"231508",x"291909",x"28180a",x"2e1c0b",x"3b2211",x"351f10",x"28190e",x"27180d",x"1f150e",x"282018",x"2c241d",x"251e16",x"211911",x"2c1b09",x"2e1d0a",x"311f0a",x"35210b",x"37230b",x"301e0a",x"321f0a",x"2d1c0a",x"251709",x"291909",x"311b0c",x"271609",x"271509",x"29170a",x"25150a",x"201309",x"191008",x"170f07",x"391f0d",x"3c210f",x"3c220f",x"3d2310",x"472910",x"432711",x"412611",x"432611",x"422611",x"3d2410",x"3b210e",x"402510",x"3d220f",x"321c0c",x"371f0d",x"351d0d",x"3d230f",x"3c2310",x"412511",x"502d14",x"351d0c",x"2c180a",x"1b1108",x"2b1b09",x"1a1107",x"181007",x"170f07",x"1d1308",x"1f1308",x"432511",x"381e0d",x"371d0c",x"3a200e",x"3b210e",x"371e0d",x"39200e",x"391f0d",x"391f0d",x"3f2410",x"3d220f",x"422611",x"412410",x"3c210e",x"3c210f",x"422611",x"422611",x"3f2411",x"3e2410",x"3e2411",x"422712",x"3a2210",x"432712",x"452813",x"432711",x"462812",x"29170a",x"2a180b",x"452811",x"452811",x"42260f",x"3d220f",x"3e230f",x"38200d",x"351e0c",x"3c210f",x"381f0d",x"351d0c",x"351d0c",x"2c180a",x"331c0b",x"311b0b",x"321c0b",x"321c0c",x"2f1a0b",x"2c190b",x"2e1a0b",x"341d0d",x"311c0c",x"311c0c",x"201309",x"20140a",x"1f130a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"452813",x"150e07",x"251409",x"281609",x"261509",x"271509",x"291509",x"281609",x"2f190a",x"2d180a",x"351d0c",x"361e0d",x"391f0d",x"341c0b",x"271408",x"271308",x"271308",x"281307",x"2a1508",x"391f0d",x"381e0d",x"391f0d",x"381f0d",x"412410",x"3d220f",x"3b210f",x"381f0e",x"3d220f",x"3b200e",x"3b200e",x"3a200e",x"3d220f",x"381f0d",x"3a200e",x"3d220f",x"3b210e",x"3a200e",x"402410",x"3c220f",x"351d0c",x"331b0b",x"351d0c",x"381e0d",x"391f0e",x"3b210e",x"361e0d",x"3b200e",x"3e2310",x"38200f",x"39210f",x"37200e",x"39200e",x"3a210f",x"3b220f",x"38200e",x"361e0d",x"3b210f",x"3f230f",x"3a200e",x"3c210f",x"432611",x"150e07",x"2d190b",x"2d1a0b",x"2d1a0b",x"2b190b",x"3a200e",x"2e1a0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f190b",x"2f190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1107",x"1b1108",x"1c1208",x"1d1308",x"1e1308",x"221508",x"201508",x"211508",x"1e1308",x"1e1308",x"1c1208",x"211508",x"201408",x"241708",x"1a1107",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"a8a8a8",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"472813",x"472813",x"3e220f",x"3d210e",x"3e210e",x"452611",x"482811",x"3d210e",x"3c210e",x"3b200e",x"3e220e",x"3d210e",x"3f230f",x"3c210e",x"3f230f",x"402410",x"432611",x"492a14",x"482b14",x"492a15",x"4a2b15",x"4b2c15",x"492a14",x"472813",x"462812",x"4a2b14",x"4a2a14",x"492a14",x"4a2b14",x"4b2c15",x"492a14",x"482913",x"452812",x"442611",x"462812",x"492a14",x"452813",x"412410",x"442711",x"412410",x"422611",x"452812",x"442711",x"442711",x"422611",x"442712",x"452812",x"452711",x"452812",x"422510",x"412410",x"432611",x"442711",x"422611",x"442712",x"452712",x"462813",x"492a14",x"452712",x"442612",x"412410",x"40230f",x"3f230f",x"442611",x"422511",x"412410",x"412410",x"40230f",x"3f230f",x"402410",x"442712",x"432611",x"432611",x"432611",x"412511",x"442712",x"452812",x"432712",x"452712",x"472913",x"492914",x"482a14",x"513018",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1308",x"1c1208",x"1c1108",x"241708",x"261809",x"211508",x"2c1b0a",x"452810",x"3c240d",x"4d2c13",x"4c2b13",x"36200c",x"291909",x"301d0a",x"2d1c0a",x"301e0a",x"2c1a0b",x"1f1309",x"1d1108",x"1f1309",x"1f1209",x"1f1209",x"1f1309",x"1e1209",x"1d1108",x"1e130a",x"2d1c0f",x"2d1c0f",x"1c1008",x"1c1208",x"1c1108",x"1b1008",x"1d1208",x"1d1108",x"1e1209",x"1e1209",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"201309",x"1d1108",x"1e1108",x"211408",x"241609",x"241608",x"261609",x"221408",x"251609",x"281809",x"2d1a0b",x"382011",x"2f1c0f",x"29190c",x"20140a",x"21160d",x"261e16",x"2b231c",x"241c15",x"211912",x"221508",x"2d1c0a",x"2b1b09",x"321f0a",x"2f1e0a",x"301f0a",x"2f1e0a",x"2e1d0a",x"261809",x"201408",x"29170a",x"2d190b",x"271509",x"251509",x"231409",x"1e1208",x"1d1107",x"180f07",x"160e07",x"321b0b",x"361e0d",x"381f0d",x"3c220c",x"3c210c",x"2f1809",x"2b1609",x"271307",x"261207",x"321a0b",x"351d0c",x"1d1108",x"331c0c",x"371e0d",x"381f0e",x"3e230f",x"3d220f",x"4c2a13",x"361e0d",x"371f0c",x"1a1107",x"170f07",x"150e07",x"1f1408",x"1e1308",x"1c1208",x"1b1108",x"150e07",x"462711",x"452611",x"381e0d",x"321a0b",x"361d0d",x"361d0d",x"371e0d",x"3d210f",x"391f0e",x"3e230f",x"3c230f",x"422612",x"432712",x"442711",x"422510",x"402411",x"412511",x"3e220f",x"3c220f",x"3b210f",x"3f230f",x"3e230f",x"3a210f",x"3c210f",x"412410",x"301b0c",x"2e1a0b",x"432812",x"432813",x"4a2a13",x"39200d",x"3a210d",x"381f0d",x"331d0b",x"361d0d",x"371f0e",x"361e0c",x"331c0c",x"351d0c",x"331c0c",x"311b0b",x"351d0c",x"311b0b",x"331c0c",x"2d190b",x"2d190b",x"2a180b",x"2c190b",x"2d190b",x"2c190b",x"2b1a0c",x"22150b",x"24160b",x"1a110a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231409",x"3d2310",x"150e07",x"351e0d",x"311b0c",x"301b0c",x"3e2310",x"3a210f",x"361e0d",x"381f0d",x"2e190b",x"371f0e",x"3a200e",x"381f0d",x"371e0c",x"361d0c",x"331b0b",x"381f0d",x"3b200e",x"3e230f",x"3f2410",x"3c220f",x"3f2410",x"3a210f",x"39200f",x"361f0e",x"391f0e",x"341d0c",x"361d0c",x"371e0d",x"3b210f",x"3b200e",x"381f0d",x"3a210e",x"402410",x"3b210f",x"3e230f",x"3b210f",x"3d220f",x"3c220f",x"3d2310",x"3c220f",x"3d230f",x"39200e",x"391f0e",x"301a0b",x"3c230f",x"3b2210",x"3a210f",x"39200e",x"311c0d",x"37200f",x"331d0d",x"351f0e",x"3d2411",x"3f2410",x"361f0e",x"38200e",x"3c220f",x"3f2410",x"3e230f",x"41230f",x"2c180a",x"321c0c",x"3a200f",x"150e07",x"150e07",x"391f0e",x"2d190b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432410",x"432410",x"432510",x"321c0b",x"341d0d",x"38200e",x"351d0d",x"351d0d",x"351d0d",x"321c0c",x"341d0d",x"341d0d",x"321c0c",x"321c0c",x"2f1a0b",x"311b0c",x"331c0c",x"341d0d",x"311c0c",x"311c0c",x"311b0c",x"311b0c",x"311b0b",x"301b0c",x"341d0d",x"331c0c",x"331c0d",x"311b0c",x"311c0c",x"311c0c",x"311c0c",x"361f0e",x"341d0d",x"2f1a0b",x"2e190b",x"2d190b",x"2b180b",x"2e190b",x"2a170a",x"2b170a",x"28160a",x"2a170a",x"2b180a",x"2b180b",x"2e1a0b",x"2f1b0c",x"2f1b0c",x"2e1a0b",x"2a190b",x"2f1b0c",x"2f1b0c",x"2c180b",x"29170a",x"301a0b",x"2e1a0b",x"29170a",x"28170a",x"2b180b",x"29180b",x"2f1c0c",x"2c190a",x"29180b",x"301b0b",x"2c1a0b",x"36200e",x"37200e",x"35200c",x"341e0c",x"341e0c",x"2f1c0b",x"2f1a0b",x"2f1c0c",x"311c0d",x"2f1b0c",x"27170a",x"2b190b",x"2e1b0c",x"2a180b",x"2b190b",x"2a190b",x"2c1a0b",x"29180b",x"25160a",x"29180b",x"29170a",x"29170a",x"27160a",x"2b180a",x"2e1a0b",x"2e1a0c",x"2a180b",x"2e1a0b",x"2d190b",x"2a180a",x"28160a",x"261609",x"29180a",x"241509",x"251509",x"2a180b",x"251509",x"241509",x"281709",x"1f1208",x"2d190a",x"281609",x"29170a",x"28170a",x"2c190b",x"2b180b",x"29170a",x"2b180b",x"28170a",x"27160a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"452712",x"452712",x"150e07",x"150e07",x"150e07",x"28170a",x"2e1a0b",x"2d190b",x"2e190b",x"2c180a",x"2d190a",x"2a180a",x"311b0c",x"301b0c",x"321c0c",x"331d0d",x"351e0e",x"331d0d",x"351e0d",x"351f0e",x"341e0e",x"351f0e",x"351f0e",x"36200f",x"321d0d",x"37200e",x"361f0e",x"37200f",x"331d0d",x"301b0c",x"29170a",x"331d0d",x"2f1b0c",x"341d0d",x"29180b",x"331c0c",x"331d0d",x"361f0e",x"341e0e",x"37200e",x"361f0e",x"27160a",x"331c0c",x"321c0c",x"37200f",x"351e0e",x"321c0d",x"2e1a0b",x"311c0d",x"361f0e",x"341e0e",x"331c0d",x"351f0e",x"331d0d",x"2e1a0b",x"2f1b0c",x"2b180b",x"2c190b",x"2c190b",x"28170b",x"2c190b",x"2e1a0b",x"2f1a0b",x"2b180b",x"2d190b",x"2d190b",x"321c0c",x"321c0d",x"311c0d",x"311c0c",x"321c0d",x"2f1b0c",x"2e1a0b",x"2c180b",x"27160a",x"29170a",x"28170a",x"2d1a0b",x"27160a",x"1d1108",x"150e07",x"150e07",x"1a1008",x"391f0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"191007",x"1a1107",x"1c1207",x"211508",x"221508",x"201408",x"2d1b0b",x"35200c",x"36200c",x"492912",x"452610",x"29190b",x"2f1d0b",x"2b1a0a",x"2f1d0a",x"2d1c0b",x"2d1c0b",x"211309",x"1f1208",x"1f1309",x"000000",x"201309",x"201309",x"201309",x"1f1209",x"1f1308",x"1e1208",x"2c1b0f",x"2c1b0f",x"191008",x"1a0f08",x"1b1108",x"1b1008",x"1d1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1d1108",x"1f1309",x"1f1208",x"1e1208",x"201309",x"211308",x"201308",x"221409",x"221409",x"2a1a09",x"251609",x"27170a",x"2a1a0a",x"2a190a",x"382011",x"311e0f",x"25170b",x"21160d",x"231911",x"29211a",x"221a12",x"241c15",x"1d1208",x"261809",x"241708",x"251708",x"291a09",x"291a09",x"261809",x"281909",x"2d1c09",x"271809",x"1f1308",x"170f07",x"27160a",x"341c0c",x"301c0b",x"2d1b0b",x"191008",x"1d1208",x"180f07",x"170e07",x"1a1107",x"3c210e",x"40240f",x"3a1f0d",x"371d0c",x"381e0c",x"3a1f0d",x"3b200e",x"3e220f",x"3c210f",x"27170a",x"331d0d",x"39200e",x"3d2310",x"3c230f",x"361e0d",x"432612",x"381f0e",x"311c0b",x"160e07",x"160e07",x"160e07",x"180f07",x"181007",x"170f07",x"1a1107",x"150e07",x"150e07",x"191007",x"472812",x"4d2c14",x"3e2310",x"402410",x"3b210e",x"351d0c",x"3a200e",x"422611",x"412511",x"3e2410",x"3f2511",x"442712",x"442712",x"452811",x"462912",x"442712",x"432711",x"3a210f",x"3e2310",x"412511",x"3e2310",x"3e220f",x"3b200e",x"311b0b",x"331c0d",x"482c12",x"492c13",x"432812",x"462811",x"3f240e",x"3b210e",x"39210d",x"3a210e",x"3d230e",x"39200d",x"3b220f",x"39210e",x"361e0c",x"311b0b",x"2c180a",x"2f1a0b",x"321c0b",x"311b0b",x"331c0c",x"311c0c",x"321c0c",x"331c0c",x"2d190b",x"2f1c0d",x"2e1b0d",x"26170b",x"1a110a",x"1d130a",x"1f130a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211309",x"381f0e",x"2b180a",x"1d1108",x"432510",x"2a180a",x"3c210e",x"38200e",x"432611",x"432611",x"412510",x"442711",x"482a13",x"452813",x"462913",x"452813",x"402712",x"412511",x"402511",x"442712",x"462813",x"402411",x"3d220f",x"3e210e",x"3e2410",x"3f2410",x"462711",x"432711",x"40240f",x"422510",x"422712",x"482a13",x"452813",x"432712",x"412511",x"432610",x"442611",x"442712",x"442712",x"452712",x"432511",x"412410",x"452812",x"462913",x"422611",x"452813",x"452812",x"3f2310",x"3a210e",x"3d220f",x"3f230f",x"3d2310",x"381f0e",x"39200f",x"3f2410",x"3e230f",x"391f0e",x"371f0d",x"402410",x"3e230f",x"442711",x"4b2b14",x"2f1b0c",x"412511",x"150e07",x"39200e",x"150e07",x"341c0c",x"311b0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351b0b",x"351b0b",x"422410",x"311b0c",x"3c230f",x"2e1a0b",x"321c0c",x"311b0c",x"361e0d",x"341d0d",x"331d0d",x"371f0e",x"3a200f",x"351e0d",x"301b0b",x"331c0c",x"311b0c",x"331c0c",x"311b0c",x"2d190b",x"2e190b",x"311a0b",x"351d0d",x"341d0d",x"331c0c",x"301a0b",x"2f1a0b",x"301a0b",x"2e1a0b",x"311c0c",x"351e0d",x"371f0d",x"371f0e",x"321c0d",x"311c0c",x"2e1a0b",x"311d0d",x"351e0e",x"331d0d",x"39210f",x"35200e",x"301c0d",x"311c0d",x"311c0d",x"2f1c0c",x"2a180b",x"2c190b",x"29180a",x"2c190b",x"2e1a0b",x"2f1a0b",x"321d0d",x"2f1a0c",x"2d190b",x"301b0c",x"2e1b0c",x"341e0e",x"2c1a0c",x"2f1b0c",x"2d1a0b",x"311c0b",x"341f0d",x"351f0d",x"301c0c",x"331e0c",x"321d0c",x"2e1b0b",x"2f1c0b",x"331f0d",x"341e0d",x"2f1a0c",x"28170a",x"2f1a0b",x"2f1b0c",x"2c190b",x"2e1a0c",x"351e0e",x"2d1a0b",x"2e1a0b",x"29170a",x"241509",x"26160a",x"27160a",x"28170a",x"27170a",x"2a180b",x"2c1a0b",x"2f1b0c",x"2d1a0b",x"321c0d",x"2c190b",x"2c190b",x"2e1a0b",x"2e1a0b",x"2c190b",x"2e1a0c",x"2c190b",x"29170a",x"251509",x"1c1108",x"2c190b",x"27170a",x"29170b",x"2b180b",x"2a180a",x"2a180a",x"2f1b0c",x"29170a",x"2d190b",x"2a180a",x"29170a",x"2e1a0b",x"2c190b",x"2a180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"472812",x"150e07",x"150e07",x"150e07",x"150e07",x"29170a",x"2f1a0b",x"2d190b",x"2e190b",x"2c180a",x"2d190a",x"29170a",x"321c0c",x"301b0c",x"311c0c",x"341d0d",x"341d0d",x"311c0c",x"361f0e",x"341e0d",x"341e0e",x"351f0e",x"341f0e",x"36210f",x"301c0c",x"37200e",x"361f0e",x"361f0e",x"331d0d",x"341d0d",x"321c0c",x"331d0d",x"331d0d",x"341d0d",x"341d0d",x"331c0c",x"341d0d",x"331e0e",x"351f0e",x"37200f",x"361e0e",x"351e0d",x"321c0c",x"311c0c",x"341e0e",x"351e0e",x"321c0d",x"2e1a0b",x"2f1b0c",x"351e0e",x"341e0d",x"331d0d",x"331e0e",x"341e0d",x"2e1a0b",x"2f1b0c",x"2d190b",x"2d1a0b",x"2a180b",x"27160a",x"2d1a0b",x"2e1a0c",x"2f1a0b",x"2a170a",x"2f1a0b",x"2d190b",x"321c0c",x"321c0d",x"321d0d",x"311c0c",x"321c0d",x"2e1a0b",x"2d1a0b",x"2b180b",x"2a180a",x"29170a",x"29170a",x"2f1b0c",x"2a180b",x"1f1208",x"150e07",x"1a1008",x"28170a",x"391f0e",x"391f0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1107",x"1b1107",x"1d1208",x"201408",x"201408",x"251708",x"271809",x"513015",x"37210c",x"472b15",x"341e0c",x"2c1a0a",x"2d1b0a",x"311e0b",x"311e0b",x"2c1b0a",x"29190a",x"2a1909",x"271809",x"281909",x"000000",x"1d1208",x"1d1208",x"1e1208",x"1d1208",x"201308",x"231609",x"2f1d0f",x"2f1d0f",x"190f08",x"1a1008",x"1c1108",x"1c1208",x"1c1108",x"1d1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1f1309",x"201309",x"1e1208",x"1f1308",x"1f1208",x"1f1208",x"201308",x"201309",x"25160a",x"251609",x"28190a",x"2a1a09",x"2a1a0a",x"27170a",x"2e1b0b",x"3a2312",x"2f1c0f",x"28180d",x"271c13",x"2e231b",x"271e16",x"241c15",x"1a1007",x"1c1107",x"1c1107",x"1f1408",x"251709",x"221508",x"231608",x"2e1d0a",x"281909",x"1f1408",x"241708",x"1a1107",x"160e07",x"160f07",x"201309",x"3a200d",x"29180a",x"201309",x"201408",x"160e07",x"180f07",x"1d1208",x"201408",x"452712",x"482b13",x"452813",x"482b13",x"4c2c14",x"452712",x"3e240f",x"24160a",x"321d0d",x"321d0d",x"331d0d",x"2f1a0b",x"3c210f",x"3f2311",x"432612",x"341d0c",x"170f07",x"170f07",x"191007",x"180f07",x"181007",x"170f07",x"180f07",x"160e07",x"150e07",x"181007",x"1b1108",x"170f07",x"452611",x"4a2a13",x"422611",x"412611",x"3e2310",x"432712",x"3e2310",x"3b210e",x"3c230f",x"412510",x"3f230f",x"42250f",x"432610",x"3f2410",x"40240f",x"38200d",x"3b200e",x"3c210f",x"3f240f",x"3f230f",x"422611",x"3f2410",x"331c0d",x"432811",x"472a12",x"442a12",x"382310",x"4a2b12",x"3b220e",x"402510",x"3e240f",x"3b220e",x"39210d",x"381f0d",x"38200d",x"371e0d",x"361f0d",x"351e0d",x"351e0d",x"371f0e",x"341d0c",x"351d0d",x"301a0b",x"311c0c",x"331c0c",x"351d0d",x"331c0c",x"341d0e",x"311c0e",x"2f1c0d",x"1e130b",x"1f130a",x"22150b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"201309",x"391f0e",x"150e07",x"271609",x"311c0c",x"351e0e",x"3a200e",x"361e0d",x"381e0d",x"371e0d",x"391f0d",x"3a1f0d",x"3a1f0d",x"3a1f0d",x"3c210e",x"3d210e",x"3a200e",x"3a200d",x"3b200e",x"381e0d",x"331c0c",x"381f0d",x"3d220f",x"3b210e",x"3b200e",x"3a200e",x"391f0e",x"341d0c",x"3a200e",x"3f230f",x"3e220f",x"3d220f",x"3a200e",x"3c210e",x"381f0d",x"3b200e",x"412410",x"3e230f",x"3a200e",x"391f0d",x"351c0c",x"381e0d",x"381f0d",x"371e0d",x"391f0d",x"391f0d",x"3d220f",x"3d220f",x"3d220f",x"3f2410",x"3d220f",x"422611",x"38200f",x"3b210f",x"3c210f",x"3f2411",x"422611",x"3c2310",x"3f2410",x"3d220f",x"3c210e",x"3a200e",x"3c220f",x"28160a",x"311b0b",x"3f220f",x"150e07",x"331c0c",x"301a0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"321a0b",x"321a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191007",x"1a1107",x"1d1308",x"1f1408",x"1f1408",x"1f1408",x"1f1408",x"1f1408",x"221608",x"221508",x"211508",x"251708",x"231608",x"201508",x"221508",x"221608",x"231608",x"221508",x"1e1308",x"1d1308",x"201408",x"201508",x"1e1308",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"462712",x"442610",x"432510",x"39200e",x"2e1a0b",x"241509",x"261509",x"251509",x"251509",x"28170a",x"261509",x"2a180a",x"2a180b",x"29180a",x"27160a",x"271609",x"1d1108",x"2b180a",x"2b180a",x"281609",x"29170a",x"26160a",x"28170a",x"27160a",x"2a180a",x"2a180a",x"2b180a",x"29170a",x"251509",x"301b0c",x"2b180b",x"29170a",x"29170a",x"29170a",x"28160a",x"2c190b",x"2d190b",x"2a180a",x"2b180a",x"2f1a0c",x"29170a",x"2b180a",x"2d1a0b",x"2a180b",x"2e1a0b",x"2f1a0b",x"271609",x"261509",x"29170a",x"251509",x"261509",x"28160a",x"28170a",x"2c190b",x"29170a",x"2c190b",x"27160a",x"2d1a0b",x"2d1a0c",x"28170b",x"27160a",x"28170a",x"2c1a0c",x"2c1a0b",x"2f1b0c",x"29170b",x"2d190b",x"2a180a",x"2c190b",x"2f1a0b",x"301b0c",x"2b180b",x"2b180b",x"2c190b",x"2c190b",x"2a180a",x"2c190b",x"2b190b",x"221409",x"1d1108",x"180f07",x"3a200e",x"3d210e",x"3b200e",x"3b200e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"191008",x"1c1107",x"1b1107",x"201408",x"1d1208",x"221508",x"321e0c",x"3b220e",x"39220d",x"39210d",x"4a2c15",x"472a13",x"4e2f15",x"331e0c",x"2e1c0a",x"2c1b0a",x"291909",x"291909",x"261709",x"261709",x"2b1b0a",x"291909",x"281909",x"201308",x"1f1308",x"201408",x"281809",x"2d1c0a",x"3e2611",x"180f07",x"180f07",x"190f08",x"1b1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1d1208",x"1d1108",x"1e1208",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1f1208",x"231509",x"211308",x"251609",x"241609",x"2a1909",x"2b1b0a",x"24160a",x"211408",x"241509",x"2a190a",x"392212",x"2c1b10",x"25180e",x"2f2117",x"282019",x"261e17",x"1b1007",x"191008",x"201408",x"1a1107",x"1e1308",x"170e07",x"241608",x"1f1308",x"211508",x"201408",x"1f1308",x"1f1408",x"170e07",x"160e07",x"160f07",x"170f07",x"201309",x"351f0d",x"28170a",x"281809",x"211509",x"160e07",x"181007",x"181007",x"160f07",x"391f0d",x"3c210e",x"42260f",x"3e230f",x"39200d",x"2f1b0b",x"2d190b",x"301b0b",x"351e0d",x"351d0d",x"311b0c",x"3a200f",x"512f16",x"361e0d",x"1a1007",x"1d1208",x"1c1108",x"191008",x"190f08",x"191008",x"191007",x"170f07",x"170f07",x"181007",x"1b1107",x"160e07",x"1b1107",x"170f07",x"512f16",x"3f220f",x"381e0d",x"381e0d",x"3d220e",x"3b210e",x"3f240f",x"3f240f",x"412510",x"432511",x"442711",x"452811",x"3d210f",x"3f230f",x"452812",x"432711",x"412611",x"3d230f",x"3e230f",x"38200d",x"331d0d",x"3b2515",x"3c2616",x"351f0d",x"3a2510",x"3e2710",x"4a2a13",x"3c220f",x"3a210e",x"3b210e",x"351d0c",x"331e0c",x"3c210d",x"3b220e",x"3b210d",x"301b0b",x"371f0d",x"351d0d",x"321c0c",x"2e190b",x"341d0d",x"321c0c",x"301a0b",x"2f1a0b",x"2d190b",x"311c0d",x"2a190c",x"2e1b0d",x"311c0d",x"21150b",x"20140b",x"19110a",x"1a110a",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"251509",x"3f2410",x"150e07",x"1f1309",x"211409",x"201309",x"26160a",x"221409",x"231409",x"29180a",x"2c190b",x"261609",x"27160a",x"29170a",x"251509",x"2b180a",x"28170a",x"29170a",x"28170a",x"28160a",x"241409",x"231409",x"241509",x"27160a",x"251509",x"251509",x"2a180b",x"241509",x"2c190b",x"2a190b",x"2e1b0c",x"2c1a0c",x"2e1b0c",x"2a180b",x"27160a",x"29170a",x"27160a",x"28160a",x"2a180a",x"28170a",x"29170a",x"221309",x"29170a",x"27170a",x"27170a",x"29170a",x"2a180a",x"29180a",x"29170a",x"241509",x"251509",x"24150a",x"27170a",x"29180b",x"29180b",x"29180b",x"2a180b",x"27160a",x"27160a",x"2a180b",x"28170a",x"27160a",x"2b180b",x"28170a",x"2c190b",x"39200e",x"150e07",x"381f0e",x"301b0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f230f",x"3f230f",x"261509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"221508",x"241708",x"221508",x"221608",x"211508",x"221608",x"221608",x"271809",x"271909",x"271909",x"251809",x"261809",x"231608",x"201408",x"201408",x"201408",x"201508",x"201408",x"1f1408",x"1c1208",x"1a1107",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442611",x"150e07",x"150e07",x"150e07",x"150e07",x"25160a",x"301b0c",x"2e1a0b",x"2e1a0b",x"2d190b",x"29170a",x"2e1a0b",x"2f1a0b",x"2e1a0b",x"2f1a0b",x"2e1a0b",x"2e1a0b",x"331c0c",x"2f1a0b",x"2e190b",x"2d190b",x"2d190a",x"2f1a0b",x"311b0b",x"301b0c",x"301b0b",x"2e190b",x"2f1a0b",x"2d180a",x"2c180a",x"2c180a",x"2c180b",x"2d190b",x"331d0c",x"2f1b0c",x"301c0c",x"211409",x"37200e",x"351f0e",x"36200e",x"301c0d",x"321d0d",x"331e0d",x"37200e",x"331d0d",x"341e0e",x"351e0e",x"331d0d",x"311c0c",x"2e1a0b",x"311b0c",x"351d0d",x"2f1b0c",x"2e1a0b",x"2a170a",x"2a180b",x"2d1a0b",x"2f1c0c",x"2d1a0c",x"2f1b0c",x"301c0c",x"2c1a0b",x"2a180b",x"2c190b",x"2d1b0b",x"2d1a0b",x"301c0c",x"2f1b0b",x"2f1a0b",x"2b190b",x"2d1a0b",x"2a170a",x"2b180a",x"2d190a",x"2b180b",x"271609",x"2a180b",x"2a180b",x"28170a",x"1d1209",x"150e07",x"150e07",x"261609",x"311b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"191008",x"191008",x"1c1208",x"1b1108",x"1d1207",x"2a190b",x"2e1b0b",x"482711",x"39210c",x"39220d",x"472a13",x"462a13",x"4b2d15",x"4f2f16",x"4c2d14",x"341f0c",x"281809",x"291909",x"2f1c0b",x"281909",x"271809",x"241709",x"241709",x"1e1208",x"1f1308",x"251709",x"2f1d0a",x"37230b",x"402711",x"180f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1e1209",x"1f1309",x"1d1108",x"1f1309",x"1e1208",x"221408",x"201308",x"261709",x"1f1308",x"241609",x"251709",x"251609",x"231509",x"201409",x"2b1a0b",x"412615",x"2f1e13",x"2f1d11",x"2f1d12",x"2c1f15",x"191007",x"1b1108",x"1c1208",x"1a1007",x"1c1207",x"1d1208",x"1d1308",x"221508",x"201408",x"221508",x"1e1308",x"1d1208",x"1f1308",x"1b1207",x"170f07",x"180f07",x"1b1107",x"1a1007",x"25160a",x"321d0c",x"2a170a",x"211308",x"170f07",x"150e07",x"150e07",x"160e07",x"391f0d",x"3d230e",x"45280f",x"3e220f",x"3f230f",x"251609",x"2c180b",x"321b0c",x"311a0b",x"3b200e",x"3b200e",x"512e16",x"3c2110",x"37200e",x"1f1208",x"1c1108",x"1d1208",x"1d1108",x"1d1208",x"1c1108",x"1b1108",x"1a1008",x"1a0f07",x"1b1107",x"170f07",x"160f07",x"160f07",x"271809",x"1b1108",x"502e15",x"472a13",x"41240f",x"41250f",x"3e220e",x"3e230f",x"41240f",x"3e220f",x"412510",x"452911",x"432711",x"432511",x"412410",x"452911",x"412610",x"432610",x"3e230f",x"462712",x"321c0c",x"311e10",x"382110",x"2d2216",x"2b1d0f",x"34210f",x"352110",x"4e2d14",x"3e230f",x"412610",x"432810",x"442910",x"3e2410",x"3a220e",x"38200d",x"321c0b",x"371f0d",x"301b0b",x"2c170a",x"2d180a",x"321c0c",x"331c0c",x"37200e",x"371f0e",x"341d0d",x"341d0d",x"301b0c",x"321d0e",x"2f1a0d",x"2b1a0d",x"2a1a0c",x"1f130b",x"20140a",x"1a110a",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"201309",x"3d2310",x"150e07",x"39200e",x"38200e",x"331c0c",x"321a0b",x"361d0c",x"3c210f",x"3b210f",x"3a200d",x"3b1f0d",x"381e0c",x"3a1f0d",x"361d0c",x"361d0c",x"381e0c",x"3e210e",x"351c0b",x"361c0b",x"341b0b",x"361d0c",x"351d0c",x"331c0b",x"381e0d",x"391f0d",x"391e0c",x"371e0c",x"361d0c",x"371d0c",x"391f0d",x"3f220f",x"3a200e",x"3a200d",x"3c200e",x"3b200d",x"3b200e",x"3a200d",x"3b200d",x"381e0d",x"391f0d",x"391f0d",x"3a200e",x"3c210e",x"3c210e",x"3d210e",x"3c210e",x"432510",x"3f2310",x"432611",x"3a200e",x"3d210f",x"3e220f",x"39200e",x"412510",x"422611",x"422511",x"3c210e",x"361e0d",x"3b200d",x"3c210e",x"381f0d",x"371d0c",x"391f0d",x"361c0b",x"321a0b",x"150e07",x"361f0d",x"2f1b0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351d0c",x"351d0c",x"2c180a",x"3d220f",x"4d2b13",x"522f15",x"4f2d15",x"4c2a13",x"462711",x"472711",x"472711",x"442510",x"4e2c14",x"512f16",x"4b2912",x"4f2d14",x"4e2c14",x"512e15",x"502d15",x"4e2c14",x"4f2d15",x"482812",x"492812",x"4b2a13",x"4f2c14",x"4b2a13",x"4d2b14",x"482812",x"4a2912",x"4a2912",x"40200d",x"43240f",x"472812",x"4a2912",x"452610",x"42240f",x"40220e",x"41230e",x"3d210d",x"41220e",x"43240f",x"42240e",x"41220e",x"3d1f0c",x"3c1f0d",x"40220e",x"41230f",x"43240f",x"3d210d",x"442510",x"3d210d",x"3b200d",x"42230e",x"42230e",x"46270f",x"4a2a11",x"4b2b11",x"482910",x"462710",x"43260f",x"47280f",x"492910",x"492a10",x"46270f",x"44270f",x"45270f",x"482910",x"4b2a11",x"4a2911",x"4c2b12",x"4c2b12",x"4d2c12",x"4c2c12",x"512f15",x"4f2d14",x"462711",x"462711",x"452611",x"472712",x"452712",x"472912",x"472712",x"3c210e",x"41230f",x"3d210e",x"3f230f",x"3d210e",x"3e220e",x"391e0d",x"391e0c",x"3b1e0c",x"3c1f0c",x"3b1f0c",x"3b1e0c",x"381c0c",x"40230e",x"40230e",x"3d1f0d",x"3e220e",x"482812",x"482812",x"482711",x"472711",x"482812",x"4b2a13",x"472711",x"492812",x"4a2913",x"492912",x"4b2a13",x"492912",x"492812",x"432510",x"452611",x"28170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3f220f",x"2a190c",x"3c220f",x"381f0e",x"29170a",x"241509",x"26160a",x"231509",x"241509",x"241509",x"231409",x"29180a",x"201208",x"201208",x"231409",x"241509",x"1e1208",x"1f1208",x"1e1208",x"211308",x"211309",x"211308",x"211308",x"211308",x"221309",x"221308",x"231308",x"231309",x"221409",x"231409",x"211308",x"150e07",x"221409",x"1f1208",x"1d1108",x"1f1208",x"211309",x"241409",x"26150a",x"261509",x"201208",x"241509",x"1f1208",x"261509",x"231409",x"231409",x"221409",x"231409",x"1d1108",x"1e1208",x"1b1108",x"27160a",x"201309",x"1c1108",x"211409",x"221409",x"201309",x"1f1208",x"211409",x"1f1208",x"241509",x"1d1108",x"191008",x"1a1008",x"1c1108",x"1d1108",x"1e1108",x"201308",x"1d1108",x"241509",x"201208",x"1f1208",x"1c1008",x"1a1008",x"1b1008",x"1f1208",x"1b1008",x"221309",x"170f07",x"150e07",x"150e07",x"1a1008",x"341d0d",x"331c0c",x"331c0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c1108",x"1e1209",x"190f07",x"1b1107",x"1a1007",x"1a1007",x"211308",x"371f0b",x"351f0d",x"37210d",x"000000",x"000000",x"000000",x"513116",x"4f3015",x"4e2d14",x"523015",x"3c230d",x"34200c",x"2d1c0a",x"281909",x"281809",x"261809",x"261809",x"1e1208",x"1f1408",x"271809",x"301e0b",x"34200b",x"442811",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f07",x"190f07",x"190f07",x"1a0f07",x"190f07",x"1a1008",x"1c1108",x"1c1108",x"1a1008",x"1d1108",x"201408",x"1f1408",x"251609",x"241609",x"221409",x"271709",x"231509",x"281809",x"221509",x"2f1b0c",x"462a17",x"342113",x"2a1b10",x"20170f",x"1a0f08",x"1b1108",x"1b1108",x"191008",x"1b1108",x"1a1007",x"170f07",x"160f07",x"190f07",x"201408",x"1e1308",x"201408",x"1a1007",x"1f1308",x"160f07",x"191007",x"1d1208",x"181007",x"191007",x"1a1107",x"361d0b",x"351e0b",x"2a190a",x"201308",x"160e07",x"170f07",x"160f07",x"170f07",x"3a210c",x"3a210d",x"381e0c",x"371e0c",x"221308",x"291609",x"2f190b",x"341d0c",x"2e190b",x"41220e",x"3f2210",x"3b230f",x"1c1108",x"231509",x"231509",x"221509",x"1c1108",x"1d1108",x"1c1108",x"1b1008",x"1a1008",x"1b1108",x"180f07",x"170f07",x"1b1107",x"251808",x"1e1308",x"1b1107",x"1c1108",x"432510",x"3d210e",x"3e230e",x"3c210e",x"40230f",x"442711",x"442611",x"41240f",x"3f240f",x"3e230f",x"42250f",x"402510",x"472812",x"40240f",x"3e220e",x"40250e",x"3a200e",x"32251c",x"291e16",x"221a12",x"2d231b",x"251b13",x"291b0d",x"27190e",x"503015",x"39210b",x"371f0b",x"41260d",x"3f260e",x"3a220d",x"38210c",x"3f250e",x"331e0c",x"37200d",x"37200d",x"331d0b",x"351d0c",x"351d0d",x"351d0d",x"361e0d",x"361e0d",x"331d0d",x"331d0d",x"2f1a0b",x"331d0e",x"301d0e",x"2b1a0c",x"2f1c0d",x"2a190d",x"19110a",x"29190c",x"25160b",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1f1208",x"381f0e",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"1d1208",x"201309",x"170f07",x"1d1208",x"1d1108",x"1a1008",x"1d1108",x"1c1108",x"180f07",x"1a1008",x"180f07",x"150e07",x"170f07",x"180f07",x"150e07",x"170f07",x"1d1208",x"201309",x"1f1208",x"1c1108",x"1c1108",x"1f1208",x"1c1108",x"211309",x"221409",x"201309",x"221409",x"1b1108",x"1b1108",x"1c1108",x"1a1008",x"1b1108",x"1b1008",x"170f07",x"170f07",x"150e07",x"150e07",x"180f07",x"180f07",x"150e07",x"180f07",x"191008",x"1c1108",x"170f07",x"180f07",x"1d1108",x"1d1108",x"150e07",x"150e07",x"190f07",x"170f07",x"191008",x"201308",x"201308",x"1f1208",x"311a0b",x"150e07",x"371f0e",x"361f0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351d0c",x"351d0c",x"2c180a",x"41240f",x"3e220f",x"3a200d",x"341d0c",x"3d210f",x"3e230f",x"3a200e",x"3b210f",x"412410",x"442711",x"442712",x"462813",x"442712",x"422511",x"452812",x"422611",x"3e220f",x"412410",x"432511",x"432611",x"412411",x"432611",x"432712",x"412511",x"402410",x"40240f",x"432510",x"432611",x"3a1f0d",x"371d0c",x"3d210e",x"412410",x"442711",x"432611",x"432711",x"412410",x"3c210e",x"3b1f0d",x"3d210e",x"432610",x"3d210e",x"3d220f",x"3d210e",x"3a200e",x"3e220f",x"371e0c",x"3b200d",x"3c210f",x"3f2410",x"432610",x"40240f",x"442610",x"3f250f",x"432710",x"442710",x"442710",x"432510",x"41260f",x"43260f",x"42260f",x"42260e",x"43280f",x"462811",x"462811",x"432711",x"452811",x"432710",x"442710",x"442610",x"42260f",x"462810",x"3f230f",x"3a210d",x"381f0d",x"361e0d",x"361e0d",x"371e0d",x"371d0c",x"331b0b",x"221107",x"281207",x"2a1408",x"361d0c",x"3a1f0d",x"371e0d",x"361d0c",x"371d0c",x"361d0c",x"361d0c",x"2e190b",x"381e0d",x"381f0d",x"3a200e",x"3c210f",x"3c210e",x"3c210f",x"3a200e",x"3e230f",x"3f230f",x"432510",x"422511",x"422611",x"442611",x"3f230f",x"3c200e",x"3e220f",x"3c210e",x"3e220f",x"3f230f",x"3e220f",x"422511",x"241509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3f220f",x"3e230f",x"391e0d",x"3f230f",x"412410",x"412410",x"3e2310",x"3b210e",x"3e220f",x"3d220f",x"3c210e",x"3c200e",x"39200e",x"381e0d",x"371e0c",x"381e0d",x"381e0d",x"381f0d",x"381e0d",x"3a200e",x"3b200e",x"3c210e",x"391f0e",x"3a200e",x"381f0e",x"361d0d",x"351d0d",x"3b210e",x"391f0d",x"361d0c",x"3b200e",x"361d0c",x"3a200d",x"3e220f",x"3f230f",x"3c210e",x"3e220f",x"3f230f",x"3d210e",x"3c200e",x"3d220f",x"3d220e",x"3f220f",x"402410",x"3b210e",x"3c210f",x"3f230f",x"3c210f",x"3a200e",x"361e0d",x"3a200e",x"381f0d",x"371f0d",x"3c210e",x"3b200e",x"3a210e",x"391f0e",x"361d0d",x"361d0d",x"381f0e",x"391f0d",x"361d0c",x"311a0b",x"321a0b",x"30190a",x"30180a",x"2e170a",x"331b0b",x"321a0b",x"2b1509",x"321a0b",x"331b0b",x"341c0b",x"341c0b",x"351c0b",x"331b0b",x"331b0b",x"381d0c",x"371d0c",x"391f0d",x"3c200e",x"412410",x"472711",x"432511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201309",x"201309",x"201409",x"1a1008",x"191008",x"2d190b",x"361d0d",x"422611",x"2d1a0b",x"2e1b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"512f14",x"4d2c12",x"512f15",x"4e2d13",x"37200d",x"2e1c0b",x"281909",x"261808",x"261809",x"211509",x"1d1108",x"201308",x"311f0a",x"452810",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f07",x"190f08",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1f1308",x"231609",x"231509",x"291909",x"2a1909",x"2a1a0a",x"281809",x"271809",x"2b1a0b",x"472b17",x"322014",x"251910",x"1a1008",x"1a1008",x"201308",x"1b1108",x"1d1208",x"1b1108",x"180f07",x"170f07",x"160f07",x"160e07",x"180f07",x"1d1208",x"1f1408",x"1d1208",x"170f07",x"1e1308",x"180f07",x"181007",x"191007",x"1b1107",x"1a1008",x"1b1108",x"301b0b",x"301b0a",x"1f1308",x"1a1008",x"160f07",x"191007",x"191007",x"271709",x"3c210e",x"2f1a0b",x"29170a",x"2c180b",x"311c0c",x"341d0c",x"361e0d",x"3d210e",x"402311",x"331d0d",x"1e1208",x"261709",x"231508",x"241509",x"241509",x"201308",x"1f1208",x"1f1208",x"1e1208",x"1d1108",x"1b1008",x"191008",x"180f07",x"231608",x"1f1408",x"1c1107",x"1c1107",x"181007",x"542f15",x"492812",x"40240f",x"3f240f",x"3f240e",x"42250f",x"3e230e",x"3c210d",x"391f0d",x"39210d",x"3d220e",x"3f240e",x"3a200d",x"371d0b",x"2b1507",x"371e0d",x"291f16",x"2a221b",x"2b221b",x"2e251d",x"2b221b",x"261d16",x"21150c",x"20160d",x"4a2a11",x"44290f",x"40250e",x"3e240e",x"40260e",x"3d230e",x"3d220d",x"39210e",x"3a210d",x"39210e",x"351e0c",x"351e0c",x"351e0e",x"351e0d",x"331c0c",x"301b0b",x"2f1a0b",x"331c0c",x"311b0c",x"321c0c",x"321c0c",x"321c0e",x"2f1b0d",x"301c0e",x"2e1c0e",x"27180c",x"25170d",x"20140a",x"1d130a",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1b1108",x"391f0e",x"1b1108",x"341e0d",x"3a210f",x"39200f",x"361f0e",x"371f0e",x"3c220f",x"381f0d",x"3a200e",x"361e0d",x"3c210e",x"3b200e",x"3b200e",x"3d210e",x"3f230f",x"3b210e",x"3b200e",x"351d0d",x"38200e",x"3a200e",x"3c210f",x"3f2410",x"3c220f",x"38200e",x"3e220f",x"3b210e",x"3c210e",x"3b210f",x"3f2410",x"381f0e",x"3c210e",x"3f230f",x"412511",x"422511",x"422510",x"412511",x"412511",x"412511",x"3f2410",x"3d2310",x"3e2310",x"3e2310",x"3c210f",x"3d220f",x"3d220f",x"3a200e",x"381f0d",x"3a200e",x"3a200e",x"3c210f",x"39200e",x"3c220f",x"381f0d",x"3a200e",x"391f0d",x"381e0d",x"381f0d",x"351d0d",x"321c0c",x"331c0c",x"381f0d",x"341d0d",x"351e0d",x"412510",x"150e07",x"3c220f",x"36200e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"41230e",x"41230e",x"402410",x"422611",x"3f2410",x"3c210f",x"3d220f",x"3d210f",x"371e0d",x"381f0d",x"3e220f",x"412410",x"3f2410",x"3e230f",x"3f230f",x"3a200e",x"3c210f",x"3f2410",x"3b200e",x"3e230f",x"402310",x"3e2310",x"422611",x"432611",x"402511",x"452712",x"482a13",x"412511",x"462813",x"422611",x"432611",x"3c210e",x"3c220f",x"3f220f",x"40230f",x"3e220e",x"3e220e",x"3f220f",x"41240f",x"3f220f",x"3f230f",x"3e230f",x"432511",x"3f230f",x"3c220f",x"432611",x"452812",x"422511",x"3f230f",x"3f240f",x"402410",x"452711",x"442711",x"452710",x"3f230f",x"3d220f",x"432611",x"432610",x"452811",x"492b12",x"4a2c12",x"4a2b12",x"482a12",x"492b12",x"482a12",x"472912",x"472911",x"432610",x"42260f",x"41240f",x"40230f",x"3e220f",x"3d220f",x"3f230f",x"3e220f",x"3c220f",x"41240f",x"3a200e",x"3c210e",x"391f0e",x"371e0d",x"391f0d",x"3a200e",x"361e0d",x"3b200e",x"3c210e",x"3d220f",x"3b210f",x"381f0e",x"3b200e",x"3c210e",x"3b200e",x"3a200e",x"391f0e",x"3e230f",x"3b210e",x"3c220f",x"381f0e",x"3e230f",x"462712",x"3f2310",x"422611",x"422611",x"422611",x"452712",x"432611",x"442712",x"402410",x"3f230f",x"3f230f",x"3d210f",x"3c210e",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3d210e",x"1f1309",x"150e07",x"1f1208",x"1a1008",x"25160a",x"2b190b",x"331d0d",x"2d1a0c",x"311c0d",x"311c0d",x"2d1a0c",x"2f1c0c",x"2d1a0c",x"311c0c",x"301b0c",x"301b0c",x"251509",x"2c180a",x"2f1a0b",x"341d0c",x"341c0c",x"371e0d",x"2e190b",x"371f0d",x"391f0e",x"39200e",x"3b210f",x"3a200e",x"3b210f",x"3e2310",x"3a200f",x"39200e",x"3a200e",x"3a200e",x"39200e",x"39200e",x"3b200e",x"381f0d",x"39200e",x"3d230f",x"3d230f",x"412411",x"422611",x"402511",x"402511",x"3d2310",x"422611",x"3d2310",x"3b210f",x"341d0d",x"2c190b",x"371e0e",x"361f0d",x"2f1a0b",x"29170a",x"2a180a",x"231509",x"170f07",x"1c1108",x"201309",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"1d1208",x"23150a",x"23150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231509",x"231509",x"412611",x"412610",x"452710",x"4c2e17",x"432d16",x"482b15",x"4d2d14",x"422711",x"442711",x"442811",x"452812",x"402410",x"3c220f",x"000000",x"000000",x"512e15",x"533016",x"522f14",x"523116",x"301d0b",x"211509",x"221508",x"1b1108",x"201308",x"160f07",x"160f07",x"150e07",x"160e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1d1208",x"1d1208",x"241609",x"231609",x"241609",x"281909",x"2c1b0a",x"311f0b",x"2b1b0a",x"301c0c",x"472b17",x"472b17",x"1a1008",x"1a1008",x"1c1108",x"1c1108",x"1b1008",x"201409",x"1b1008",x"180f07",x"170f07",x"160e07",x"160e07",x"160e07",x"170f07",x"190f07",x"1a1007",x"180f07",x"170f07",x"180f07",x"170f07",x"180f07",x"1a1008",x"191008",x"1c1108",x"201409",x"311c0b",x"2b190a",x"241509",x"191007",x"170f07",x"150e07",x"191007",x"311c0c",x"331c0c",x"2e1a0b",x"361e0d",x"331c0c",x"38200e",x"3b200e",x"4d2b13",x"331d0d",x"1f1208",x"1f1208",x"221408",x"231509",x"221509",x"211409",x"25160a",x"201208",x"201208",x"201309",x"1f1309",x"1d1208",x"1b1108",x"1e1208",x"1a1008",x"231608",x"1c1207",x"1f1408",x"160f07",x"160e07",x"502e15",x"4b2a12",x"452711",x"40230f",x"41250f",x"442610",x"41250f",x"42260f",x"432711",x"442610",x"41250f",x"422610",x"3f230f",x"331c0b",x"201811",x"221a12",x"261e16",x"2c241d",x"271f18",x"2a211a",x"292019",x"20170e",x"24190f",x"4c2c12",x"3d230d",x"3a220d",x"41260e",x"432810",x"3d240e",x"3c230e",x"3a210e",x"361f0d",x"39210d",x"39220e",x"39210e",x"371f0d",x"341e0d",x"341e0d",x"351e0e",x"341d0d",x"321c0c",x"2f1a0c",x"351d0d",x"331c0c",x"2f1c0d",x"2e1b0d",x"2d1a0d",x"2f1c0d",x"28180c",x"20140a",x"291a0d",x"29190d",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"241509",x"3a200e",x"37200f",x"2b190b",x"4b2b14",x"28180b",x"3b2210",x"3e2410",x"412511",x"412511",x"3d220f",x"3c210f",x"3e220f",x"3a200e",x"391f0d",x"3b200d",x"381e0c",x"381f0d",x"361e0d",x"361e0d",x"321c0b",x"3a200d",x"371e0d",x"391f0d",x"381f0d",x"371e0d",x"361e0d",x"361e0d",x"381e0d",x"391f0d",x"371d0c",x"331c0b",x"311a0a",x"351b0b",x"361d0c",x"381d0c",x"381e0d",x"3a200d",x"3a200e",x"391f0d",x"361d0c",x"30180a",x"30190a",x"331b0b",x"3b200e",x"432611",x"402411",x"412511",x"3e2310",x"3c210f",x"3c210e",x"391f0d",x"3c210e",x"3c220f",x"381f0e",x"3f2310",x"3f2310",x"3d210e",x"3d230f",x"38200e",x"3d230f",x"422510",x"311b0c",x"442711",x"150e07",x"3a210f",x"150e07",x"402410",x"351e0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462711",x"462711",x"462a14",x"482b14",x"412511",x"3d2310",x"422612",x"452914",x"3f2511",x"412512",x"442712",x"3d220f",x"3f2410",x"3e2310",x"412612",x"402410",x"3b210f",x"3d230f",x"391f0e",x"3e2310",x"412612",x"3d2311",x"412511",x"3d2310",x"3c2310",x"3d2310",x"402511",x"3d2310",x"402511",x"412511",x"3a220f",x"39200e",x"3c210f",x"3b210e",x"3c210e",x"381e0d",x"371e0c",x"361d0c",x"351d0c",x"371d0c",x"381e0d",x"371e0d",x"361e0d",x"321b0b",x"361e0d",x"351d0c",x"381f0d",x"361e0d",x"361e0d",x"381f0d",x"351d0c",x"361d0c",x"331c0b",x"331c0b",x"31190a",x"2e180a",x"311a0b",x"321b0b",x"391f0c",x"371e0c",x"3c220d",x"39210d",x"3b210d",x"361e0b",x"361e0b",x"3b210c",x"3f240e",x"3f240f",x"3c210f",x"3e2310",x"3a210e",x"3a200f",x"3c210f",x"3a200e",x"371e0d",x"351d0d",x"3b210f",x"3b210f",x"3a210f",x"351d0c",x"3a200e",x"3a200e",x"39210f",x"3f2410",x"371f0d",x"3b210f",x"38200e",x"361f0e",x"361e0d",x"3c220f",x"3d230f",x"3c220f",x"3f2410",x"3e2411",x"3a210f",x"432812",x"3a210f",x"3d2411",x"412612",x"452913",x"412612",x"472a14",x"442813",x"472a14",x"472a14",x"4b2d16",x"472a14",x"3f2310",x"3f2411",x"462914",x"442713",x"422611",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3d210e",x"391f0e",x"4f2f16",x"482a14",x"432712",x"3f2411",x"3f2511",x"3c2210",x"3f2410",x"3f2511",x"3c2310",x"3b220f",x"3b220f",x"3a210f",x"351e0e",x"3a210f",x"351e0d",x"381f0e",x"361f0d",x"311c0c",x"2c180a",x"2f1a0b",x"311b0b",x"301a0b",x"29170a",x"311b0b",x"311b0c",x"2f1a0b",x"351d0d",x"351d0c",x"351d0d",x"321c0c",x"331c0c",x"311c0c",x"331c0c",x"311b0c",x"2f190b",x"321c0b",x"30190b",x"2d170a",x"2c170a",x"30190a",x"2f190b",x"311b0b",x"331c0c",x"331c0c",x"331c0c",x"2d180a",x"271509",x"2a1609",x"2a170a",x"311b0c",x"341d0d",x"38200e",x"341d0d",x"371f0e",x"331d0d",x"2f1a0b",x"311b0b",x"331c0c",x"361e0d",x"371f0e",x"381f0e",x"2f1b0b",x"2e1a0b",x"351e0d",x"351e0d",x"361f0e",x"321c0c",x"2e1b0b",x"361f0e",x"39200f",x"341d0d",x"39200e",x"321c0c",x"321c0d",x"301c0c",x"2f1b0c",x"2e1a0c",x"341f0e",x"38210f",x"4d2d15",x"462913",x"4f2e16",x"4f2e16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432611",x"442812",x"4f3118",x"472a13",x"4a2b14",x"462711",x"3f230e",x"3c230f",x"3e240f",x"442811",x"452812",x"3a210e",x"3c2310",x"38200f",x"27170a",x"2e1b0c",x"2d1a0b",x"553317",x"513116",x"43250f",x"331e0c",x"231609",x"1b1107",x"170e07",x"160e07",x"161009",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f08",x"180f08",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1c1208",x"201409",x"201409",x"221609",x"2c1b0a",x"2c1c0a",x"2b1b0a",x"2e1d0a",x"221509",x"2e1b0b",x"2e1b0b",x"1b1008",x"1a1008",x"1e1209",x"21150a",x"201408",x"1c1108",x"1d1208",x"191008",x"1a1008",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"170e07",x"170e07",x"191107",x"180f07",x"180f07",x"1b1007",x"1c1108",x"1b1108",x"1f1409",x"201409",x"1f1409",x"261609",x"2d190a",x"2d1a0b",x"211409",x"1b1107",x"181007",x"181007",x"29180a",x"2e1a0a",x"311c0b",x"321c0c",x"321c0c",x"2d190a",x"452611",x"4e2c14",x"1a1008",x"211509",x"1d1108",x"1d1208",x"211408",x"1f1308",x"251609",x"201308",x"1d1108",x"1c1008",x"1d1108",x"1c1108",x"1c1108",x"1b1008",x"190f08",x"191007",x"170f07",x"160e07",x"1c1108",x"160e07",x"160e07",x"191008",x"563318",x"4c2c13",x"482911",x"452811",x"452811",x"42250f",x"3f240f",x"462811",x"472911",x"442711",x"452711",x"442710",x"331d0c",x"201811",x"211911",x"211912",x"261d16",x"231b14",x"2c241d",x"292018",x"20160e",x"20160d",x"4d2d13",x"3f250e",x"3f250f",x"412710",x"452911",x"472c11",x"472b13",x"442911",x"412710",x"412811",x"402611",x"3f2611",x"3d2411",x"3b2310",x"402612",x"412713",x"402612",x"361e0e",x"371f0e",x"38200f",x"38210f",x"37200f",x"372111",x"341f0f",x"301c0e",x"28180c",x"29190c",x"1b120a",x"28190d",x"19110a",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"28170a",x"371e0d",x"150e07",x"39200e",x"321c0c",x"301b0c",x"3c220f",x"311c0c",x"2e1a0b",x"311b0b",x"2a1709",x"281509",x"29170a",x"2f1a0b",x"331c0c",x"361e0d",x"39200e",x"311c0c",x"39200e",x"381f0e",x"351e0d",x"331c0c",x"311b0c",x"351d0d",x"2d190b",x"2c190b",x"2d180a",x"2d190b",x"2e1a0b",x"301b0c",x"351d0d",x"381f0e",x"371f0d",x"371e0c",x"341c0c",x"331c0c",x"351d0c",x"311b0b",x"301a0b",x"301a0b",x"311b0b",x"2e1a0b",x"2e190b",x"2f190b",x"2b180a",x"301b0b",x"361e0d",x"331d0d",x"351d0d",x"301a0b",x"331c0c",x"341d0c",x"361f0e",x"361e0e",x"311c0d",x"38200f",x"3e2410",x"3a210e",x"381f0e",x"38200e",x"3e2410",x"462813",x"311c0d",x"402511",x"452712",x"150e07",x"1b1108",x"3e2310",x"311c0d",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b1f0d",x"3b1f0d",x"452812",x"422612",x"402511",x"482a14",x"432712",x"462812",x"402511",x"3f230f",x"402410",x"412511",x"402411",x"402410",x"361e0d",x"3d220f",x"3b200e",x"3f230f",x"3d220f",x"3d220f",x"3c210f",x"3c210f",x"3f230f",x"3f230f",x"3a200e",x"3e220f",x"3c210e",x"412410",x"422510",x"3e220f",x"3f230f",x"361d0d",x"361c0c",x"31190a",x"351b0b",x"3a1f0d",x"391f0d",x"3d210e",x"402410",x"432611",x"432611",x"3f2310",x"432611",x"412410",x"3b200e",x"3d210f",x"3b200e",x"3b200d",x"321b0b",x"381f0d",x"381e0d",x"3e230f",x"402410",x"402410",x"3f240f",x"3b200e",x"391f0d",x"3f230f",x"3c220e",x"3d220e",x"381f0d",x"39200c",x"3b210e",x"3d220e",x"3f240e",x"3b220c",x"3f230d",x"40240e",x"41250f",x"452811",x"412510",x"41240e",x"41250f",x"3f230e",x"40240f",x"432611",x"482a13",x"472913",x"452812",x"472912",x"41250f",x"41250f",x"422611",x"422612",x"412511",x"442712",x"422511",x"432612",x"452812",x"3d2310",x"412511",x"432611",x"442712",x"442813",x"452813",x"462813",x"402410",x"3b200e",x"3d210f",x"3d220f",x"432611",x"472914",x"472913",x"452712",x"442712",x"472914",x"462913",x"462913",x"482a14",x"452713",x"442712",x"422511",x"2a180a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3f230f",x"3f230f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181008",x"191008",x"1d1108",x"191008",x"170f07",x"1a1008",x"1a1008",x"1c1108",x"1b1008",x"1b1008",x"1a1008",x"1c1108",x"170f07",x"1b1108",x"190f07",x"191008",x"1c1108",x"1b1008",x"1e1208",x"1f1208",x"1b1108",x"241509",x"1f1309",x"1d1108",x"221409",x"1c1108",x"1e1209",x"201309",x"1e1209",x"1d1208",x"170f07",x"23150a",x"231409",x"201309",x"160e07",x"160e07",x"1d1208",x"1c1108",x"1a1008",x"160e07",x"160e07",x"160e07",x"170f07",x"150e07",x"150e07",x"150e07",x"170f07",x"2a180b",x"2a180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452813",x"452813",x"361e0c",x"271809",x"261709",x"281809",x"2a1909",x"261609",x"281809",x"251609",x"201208",x"2c180a",x"27170a",x"2e1b0c",x"2d1a0b",x"2a180b",x"361f0e",x"211409",x"44260f",x"45260f",x"201308",x"2a180b",x"150e07",x"181109",x"171009",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"180f08",x"180f08",x"180f08",x"191008",x"191008",x"191008",x"191008",x"190f08",x"180f07",x"211409",x"1b1107",x"231609",x"2d1d0a",x"28190a",x"291a0a",x"221609",x"28190a",x"2d1b0a",x"1c1108",x"1c1108",x"1e1209",x"1d1208",x"1d1208",x"1c1208",x"1c1108",x"1a1008",x"180f08",x"1a1107",x"170f07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"160e07",x"180f07",x"1f1408",x"1d1208",x"201408",x"1c1107",x"1f1308",x"211409",x"1f1409",x"201409",x"201509",x"2d1b0b",x"361e0c",x"271509",x"231509",x"251509",x"2c190b",x"2b1a0b",x"341e0c",x"3e240f",x"3d240f",x"3c220f",x"4a2a13",x"472711",x"311c0d",x"1f1309",x"1d1208",x"1c1108",x"1e1208",x"271709",x"241609",x"29190a",x"211309",x"211409",x"211309",x"1f1208",x"1f1208",x"1d1108",x"1b1008",x"190f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"191008",x"533016",x"4a2a12",x"41250f",x"42250e",x"472a10",x"472911",x"4c2d12",x"4e2f13",x"492b14",x"4f2f15",x"3b220d",x"331d0c",x"331d0c",x"211912",x"211913",x"211811",x"221912",x"292019",x"2a221a",x"231911",x"21170e",x"502d14",x"442810",x"452911",x"452911",x"422811",x"432812",x"422610",x"381f0d",x"3a210d",x"351e0d",x"321d0c",x"37200f",x"39210f",x"37200f",x"3a200f",x"3d2310",x"37200f",x"37200f",x"37200f",x"351f0e",x"361f0e",x"331d0d",x"2e1a0b",x"301d0e",x"2f1c0e",x"2a190c",x"28180c",x"21150b",x"19110a",x"20140c",x"25180c",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"361d0c",x"150e07",x"211409",x"2f1a0b",x"321c0d",x"321d0d",x"381f0e",x"381f0e",x"391f0e",x"331c0c",x"341d0c",x"351d0c",x"331c0c",x"381f0d",x"3a200e",x"39200d",x"301a0b",x"341c0c",x"321b0b",x"301a0b",x"361e0d",x"381f0d",x"301a0b",x"301a0b",x"2f190b",x"361d0c",x"341c0c",x"341c0c",x"381f0d",x"351d0c",x"321b0b",x"311a0b",x"2f190a",x"30180a",x"331b0b",x"361d0c",x"341d0d",x"3c220f",x"3a200e",x"3a200e",x"3b210f",x"3b210f",x"3c220f",x"3b220f",x"3f2410",x"412511",x"3e2310",x"391f0e",x"361d0d",x"351d0d",x"391f0e",x"381f0e",x"3e2310",x"3c2210",x"3e220f",x"3c210f",x"39200e",x"391f0d",x"3b200e",x"3c220f",x"462812",x"150e07",x"39210f",x"321c0c",x"301c0d",x"341e0d",x"371f0d",x"37200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f230f",x"3f230f",x"452812",x"432712",x"432712",x"432612",x"452814",x"482a14",x"462914",x"462914",x"492a14",x"452813",x"432612",x"462913",x"412612",x"412511",x"432712",x"462913",x"402410",x"3e2310",x"432712",x"412611",x"422611",x"3e2310",x"3d220f",x"3d210e",x"3c210e",x"412510",x"432712",x"432611",x"452712",x"3d210e",x"3b200e",x"3a200e",x"3a200e",x"391f0d",x"3d210f",x"3d210e",x"3f220f",x"3e220f",x"391f0d",x"3b200e",x"371d0c",x"3b200d",x"3d210f",x"3b200e",x"371e0c",x"391f0d",x"381e0d",x"351c0b",x"3a1f0d",x"3a200d",x"3a200d",x"381e0d",x"391e0d",x"351c0b",x"351b0a",x"371d0b",x"3d220d",x"41240f",x"41260f",x"41250f",x"41250f",x"432610",x"40240f",x"3f240f",x"412510",x"402510",x"462811",x"452911",x"442810",x"3c210e",x"3d220e",x"3e230e",x"42260f",x"482912",x"482912",x"432611",x"422510",x"3f230f",x"3f230f",x"3c210d",x"40230f",x"3d230f",x"412610",x"3d230f",x"412510",x"442713",x"3f2410",x"432711",x"422612",x"3f2411",x"422612",x"432612",x"482913",x"452712",x"422611",x"452812",x"412511",x"432611",x"472914",x"432712",x"482a14",x"492a14",x"452712",x"482a14",x"492a14",x"492a14",x"482a14",x"472914",x"482a15",x"4c2c15",x"2a180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3c210e",x"25150a",x"150e07",x"221409",x"38200f",x"29180b",x"231509",x"231409",x"201309",x"1e1208",x"180f07",x"1f1208",x"201309",x"150e07",x"1a1008",x"1c1108",x"1e1208",x"1a1008",x"1b1108",x"180f07",x"1d1108",x"1c1108",x"1a1008",x"201308",x"251509",x"221409",x"201208",x"211308",x"241509",x"211309",x"261509",x"221309",x"281609",x"261509",x"271609",x"2c180a",x"2a170a",x"261509",x"29160a",x"271509",x"251408",x"231308",x"251409",x"27160a",x"1e1208",x"231509",x"26160a",x"27160a",x"29170a",x"27160a",x"201309",x"25160a",x"28170a",x"26160a",x"221409",x"241509",x"231409",x"28170a",x"221409",x"241509",x"2b190b",x"26160a",x"26160a",x"27160a",x"241509",x"211309",x"201309",x"1f1309",x"1e1208",x"1d1208",x"1f1209",x"150e07",x"211409",x"211409",x"1e1209",x"150e07",x"1b1108",x"191008",x"150e07",x"150e07",x"150e07",x"180f08",x"3a210f",x"3c210e",x"3c210e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b2b1f",x"3b2b1f",x"201308",x"261609",x"29190a",x"29190a",x"27170a",x"2b1a0a",x"29180a",x"27170a",x"251609",x"241509",x"221409",x"231509",x"211409",x"201309",x"1f1208",x"211309",x"211309",x"492811",x"43240e",x"3f220e",x"150e07",x"191109",x"181009",x"171009",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"1f1308",x"1b1108",x"251708",x"28190a",x"261708",x"261808",x"261708",x"2c1b0b",x"1c1108",x"1e1209",x"1e1209",x"1e1209",x"211508",x"201408",x"201409",x"1b1008",x"1a0f08",x"180f08",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"170e07",x"180f07",x"1c1108",x"221608",x"271909",x"231608",x"1e1308",x"231509",x"211509",x"221509",x"231609",x"221509",x"201409",x"2f1c0a",x"311c0b",x"2b180a",x"2d190b",x"2d1a0b",x"321c0b",x"3e250e",x"351e0c",x"38200d",x"42240e",x"4a2912",x"251509",x"191008",x"190f07",x"1c1108",x"1f1308",x"1d1108",x"231409",x"201308",x"1f1208",x"1f1208",x"1f1208",x"1e1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"170f07",x"191008",x"502f14",x"472a10",x"472910",x"4f2f12",x"4e2d11",x"4e2f12",x"4d2e13",x"492a12",x"331d0b",x"361f0c",x"231608",x"261809",x"201508",x"1f1408",x"180f07",x"211911",x"271b13",x"231911",x"231911",x"20160e",x"362010",x"452912",x"462a11",x"3f2610",x"442910",x"3e230f",x"361e0d",x"3f2510",x"39200f",x"3c220e",x"3a210f",x"38200f",x"3d2310",x"3a220f",x"371f0e",x"3a210f",x"3a210f",x"38200f",x"361f0e",x"351f0e",x"351f0f",x"2a190b",x"2f1c0d",x"301c0d",x"311d0f",x"29190c",x"2d1b0e",x"24170c",x"1f140b",x"22150b",x"25170b",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25150a",x"391f0d",x"150e07",x"2d190b",x"3a210f",x"371f0e",x"311c0d",x"331d0d",x"38200e",x"361e0d",x"371f0d",x"3b210f",x"371f0e",x"39200e",x"371f0d",x"351d0d",x"341d0d",x"321c0c",x"361e0d",x"341c0c",x"2e1a0b",x"331c0c",x"361e0d",x"341c0c",x"351d0d",x"341d0c",x"361e0d",x"321c0b",x"321b0b",x"381f0d",x"371e0d",x"351d0c",x"351d0c",x"331c0c",x"341c0c",x"351d0c",x"341c0c",x"361e0c",x"3c210e",x"39200e",x"381f0e",x"331c0c",x"391f0d",x"3c210f",x"331c0c",x"3b220f",x"3b210f",x"3a200f",x"381f0e",x"381f0e",x"39200e",x"39200e",x"3a200e",x"39200e",x"331c0c",x"311b0b",x"3b220f",x"3c220f",x"3a200e",x"402411",x"3e2410",x"331e0e",x"24150a",x"331c0c",x"3c2210",x"3c2310",x"351f0e",x"39210f",x"3b2210",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b1508",x"2b1508",x"452611",x"412410",x"412410",x"3f230f",x"422410",x"3f220f",x"422410",x"3f230f",x"3d220f",x"3f230f",x"492912",x"472812",x"462913",x"512f16",x"502f16",x"512f16",x"4f2e16",x"492912",x"4b2b13",x"4b2a13",x"4a2a13",x"4b2a13",x"4b2a13",x"4b2b13",x"512e15",x"502e15",x"4b2b14",x"502f16",x"4d2c14",x"4a2913",x"4b2a12",x"4b2a13",x"4b2a12",x"4a2913",x"4c2b13",x"472812",x"4a2912",x"4f2c13",x"4a2912",x"452610",x"462610",x"452510",x"482811",x"482811",x"482711",x"4a2811",x"492811",x"4a2912",x"43240f",x"472710",x"4a2912",x"452610",x"472610",x"472710",x"452510",x"482711",x"482610",x"492810",x"472710",x"4d2c13",x"4c2a12",x"4d2c13",x"4b2a12",x"502d14",x"492811",x"4c2b13",x"4b2a14",x"4c2b14",x"4a2913",x"462711",x"4d2c14",x"4e2c15",x"492812",x"4a2912",x"432510",x"472611",x"4a2912",x"4f2d14",x"4a2812",x"4a2912",x"4c2b14",x"523017",x"553318",x"43230e",x"4e2c14",x"4b2b14",x"4b2b14",x"4b2c14",x"4b2b13",x"482812",x"4d2c15",x"4e2d15",x"4a2913",x"4a2913",x"4b2912",x"4a2912",x"4e2c14",x"452611",x"492912",x"452610",x"462711",x"4b2a13",x"4b2a12",x"492812",x"482712",x"492812",x"482811",x"442510",x"442510",x"452510",x"2b180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200e",x"502e15",x"482913",x"492a14",x"3e230f",x"331d0d",x"361e0d",x"371f0e",x"371f0e",x"381f0e",x"341d0d",x"341e0d",x"351e0e",x"321d0d",x"2f1c0c",x"341d0d",x"331d0d",x"38200e",x"371f0e",x"341d0d",x"341d0d",x"39200e",x"3b200e",x"3b210f",x"3a200e",x"3c210e",x"391f0d",x"381f0d",x"371e0d",x"3f230f",x"3b200d",x"3c210f",x"3a200d",x"3d220f",x"3b200d",x"3b200d",x"432510",x"3f230f",x"3b200d",x"361d0c",x"3a200e",x"3c210d",x"3b200e",x"3e220e",x"381f0d",x"422510",x"442611",x"3c210f",x"3f220f",x"422510",x"402410",x"3d220f",x"462812",x"3d220f",x"381e0d",x"351d0c",x"361d0c",x"3a1f0d",x"361d0c",x"371d0d",x"391f0d",x"3b200d",x"3c210e",x"3d220e",x"3a200d",x"3c210e",x"3c210f",x"3d230f",x"391f0d",x"3e220f",x"412511",x"3f230f",x"40230f",x"3f230f",x"3b1f0d",x"3c210f",x"3d220f",x"3d210e",x"3b200e",x"3d220e",x"3d210e",x"3b200e",x"3d210e",x"3d220e",x"3d220e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b2118",x"2b2118",x"371e0d",x"201308",x"211309",x"211309",x"261709",x"27170a",x"231509",x"25160a",x"241609",x"201308",x"221409",x"221409",x"221409",x"211309",x"211409",x"201308",x"201308",x"29170a",x"41230e",x"432610",x"3a2110",x"341e0e",x"382010",x"412512",x"412512",x"422512",x"442712",x"422510",x"412410",x"432510",x"452712",x"452611",x"432511",x"442510",x"412410",x"442610",x"442510",x"462611",x"442611",x"442611",x"422410",x"41240f",x"462710",x"482811",x"452710",x"472810",x"452610",x"4d2c13",x"4e2c13",x"502f14",x"1b1108",x"1c1108",x"1b1008",x"1b1008",x"1b1108",x"1a1108",x"191008",x"1a1108",x"201408",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"180f07",x"1a1007",x"271809",x"251808",x"221508",x"211508",x"2d1c09",x"241709",x"221609",x"271809",x"281909",x"241609",x"281909",x"281809",x"37200d",x"3b220f",x"361f0d",x"361f0d",x"371e0c",x"3d220e",x"472a10",x"442610",x"502d15",x"2a180b",x"1c1108",x"1d1208",x"191008",x"1b1008",x"1e130a",x"20140b",x"1d1108",x"1e1208",x"201309",x"201208",x"201208",x"201308",x"1f1208",x"1f1208",x"1d1108",x"1c1108",x"1a1008",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"522e13",x"563314",x"523113",x"503013",x"4e2e12",x"4a2b11",x"3b220d",x"1c1207",x"1f1408",x"1f1408",x"201408",x"251708",x"1d1208",x"1c1208",x"170f07",x"160e07",x"23190f",x"231911",x"21170e",x"331e10",x"3f240f",x"492b12",x"452812",x"422610",x"3c220e",x"3c220e",x"3f240f",x"3a200e",x"371e0d",x"371e0d",x"341c0c",x"351d0d",x"3d220f",x"3c220f",x"381f0e",x"2d190b",x"341d0d",x"311c0c",x"321c0c",x"321c0c",x"29170a",x"2e1a0b",x"2f1a0b",x"29170a",x"2e1c0d",x"2c1a0d",x"2a1a0d",x"28190c",x"27180c",x"371f0f",x"452813"),
(x"150e07",x"150e07",x"150e07",x"28170a",x"3a200d",x"150e07",x"271509",x"2f1a0b",x"331c0d",x"2d1a0b",x"150e07",x"3c210f",x"3e220f",x"3d220f",x"3d220f",x"3e220f",x"3d220f",x"3f230f",x"432611",x"412410",x"402410",x"3c220f",x"422511",x"3d220f",x"402310",x"3f2410",x"452812",x"462913",x"3e2310",x"3d210e",x"3d220f",x"422510",x"422510",x"41230f",x"422510",x"3a1f0d",x"391e0c",x"422510",x"422510",x"432511",x"422510",x"422510",x"432611",x"432610",x"3b210f",x"432711",x"462712",x"462812",x"462913",x"452812",x"432612",x"472913",x"452812",x"432611",x"442712",x"432611",x"422511",x"412410",x"3e2310",x"40230f",x"3f220f",x"422510",x"442611",x"40210e",x"150e07",x"28160a",x"2f1a0b",x"371e0d",x"351c0c",x"2a170a",x"3d2310",x"3a210f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39200d",x"39200d",x"3c210e",x"3b210e",x"341d0d",x"351d0d",x"301b0c",x"351d0d",x"351d0d",x"311b0c",x"361e0d",x"331c0c",x"341d0d",x"492912",x"2b180b",x"1c1108",x"1c1108",x"150e07",x"170f07",x"150e07",x"150e07",x"190f08",x"1c1108",x"1b1008",x"190f07",x"190f07",x"190f07",x"1a1008",x"180f07",x"1a1008",x"1a1008",x"170f07",x"1a1008",x"150e07",x"1c1108",x"170f07",x"150e07",x"180f08",x"1d1208",x"1a1008",x"1f1309",x"190f08",x"170f07",x"1f1209",x"170f07",x"150e07",x"150e07",x"1d1108",x"1e1208",x"1a1008",x"1b1008",x"1d1108",x"1d1108",x"150e07",x"150e07",x"1a1008",x"170f07",x"1d1208",x"170f07",x"180f08",x"150e07",x"150e07",x"150e07",x"1b1108",x"201309",x"1b1108",x"221608",x"1f1308",x"201409",x"2a1a09",x"201408",x"281909",x"1a1107",x"150e07",x"180f08",x"150e07",x"1a1008",x"180f08",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"1d1208",x"1f1208",x"150e07",x"1b1108",x"1f1309",x"221409",x"1b1108",x"150e07",x"1f1309",x"1f1209",x"1d1108",x"1d1108",x"201309",x"1c1108",x"1a1008",x"371f0e",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"29170a",x"2b180a",x"2d190b",x"2b170a",x"2b170a",x"221107",x"29160a",x"2c180a",x"2a170a",x"2d1a0b",x"2c190b",x"29170b",x"2f1a0b",x"311b0c",x"341d0d",x"2c190b",x"311c0c",x"371f0e",x"381f0e",x"321c0c",x"351d0d",x"38200e",x"28170a",x"26160a",x"301b0c",x"38200e",x"361f0e",x"311c0d",x"1c1108",x"27160a",x"301b0b",x"2f1a0c",x"2b180b",x"241509",x"1d1108",x"261509",x"251509",x"26160a",x"25150a",x"180f07",x"180f07",x"190f07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f08",x"1a1008",x"160e07",x"180f08",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"1b1008",x"2d1a0c",x"2d1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b180a",x"2b180a",x"1f1208",x"27170a",x"231409",x"231409",x"231409",x"231409",x"231509",x"231509",x"241609",x"231509",x"24150a",x"24150a",x"24150a",x"24150a",x"231409",x"29180b",x"27160b",x"29170a",x"27160a",x"2e1a0b",x"311c0c",x"331d0e",x"311b0c",x"2e1a0b",x"2f1a0b",x"3a200e",x"3f2310",x"341e0d",x"271809",x"211408",x"221409",x"1f1208",x"432511",x"442510",x"412410",x"211309",x"231509",x"211409",x"211309",x"201309",x"2a190b",x"41240f",x"211409",x"201309",x"211409",x"28180a",x"2a190a",x"2c1b0a",x"1d1108",x"1a1008",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1b1008",x"1a1008",x"1c1208",x"1a1008",x"180f07",x"170f07",x"160e07",x"160e07",x"190f07",x"191007",x"1b1107",x"1a1007",x"1c1208",x"251708",x"231608",x"2c1b09",x"261808",x"281909",x"35210b",x"311e0a",x"28190a",x"271809",x"29190a",x"28190a",x"281809",x"291909",x"3f240f",x"381f0d",x"3a210d",x"39210e",x"3e240e",x"3f240f",x"522f15",x"23150a",x"221409",x"1a1008",x"1e1308",x"1d1308",x"1e130a",x"1d130a",x"1e130b",x"20140a",x"1f1309",x"1f1309",x"201308",x"1f1208",x"1d1108",x"1e1208",x"1f1308",x"1e1208",x"1d1108",x"1a1008",x"180f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"543114",x"573315",x"4f2f13",x"513013",x"4f2f12",x"43270f",x"3b220c",x"321c0b",x"2b190b",x"1e1308",x"1c1208",x"211508",x"251809",x"201408",x"201408",x"170e07",x"160f07",x"211810",x"23170f",x"2d1a0d",x"432610",x"38200d",x"3c220e",x"44270f",x"3e230e",x"371f0d",x"3b220e",x"40230f",x"391f0e",x"381f0e",x"3f230f",x"3f2310",x"3e2310",x"3d2310",x"432712",x"412511",x"3c210f",x"3b200e",x"412511",x"412511",x"3f2511",x"3b220f",x"3b200e",x"3c220f",x"3d2310",x"3e2311",x"371f0f",x"3a2010",x"361f0f",x"25160c",x"25160c"),
(x"150e07",x"150e07",x"150e07",x"241509",x"3a1f0d",x"150e07",x"201308",x"2e1a0b",x"311b0b",x"29170a",x"2d1a0b",x"311b0c",x"2e1a0b",x"321c0c",x"301b0b",x"321c0c",x"321c0c",x"341d0c",x"321c0c",x"381f0e",x"381f0e",x"301b0c",x"2f1a0b",x"351d0d",x"361e0d",x"311b0b",x"2d190b",x"2a170a",x"2c180a",x"29170a",x"2f1a0b",x"321c0c",x"311b0c",x"301a0b",x"321c0c",x"341d0d",x"331c0c",x"331c0c",x"2d190b",x"301a0b",x"301a0b",x"301a0b",x"311b0b",x"321c0c",x"351d0d",x"321c0c",x"301a0b",x"2d170a",x"2b1609",x"251208",x"231107",x"221006",x"221006",x"211106",x"211006",x"2e180a",x"301a0b",x"2f190b",x"2f190b",x"341c0c",x"341d0c",x"381f0e",x"3c220f",x"371f0e",x"422511",x"231509",x"38200e",x"39200e",x"38200f",x"301b0c",x"39200f",x"3b2210",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39200d",x"3c210e",x"3b210e",x"341d0d",x"351d0d",x"301b0c",x"351d0d",x"351d0d",x"311b0c",x"361e0d",x"331c0c",x"2a180b",x"2a180b",x"341e0d",x"25150a",x"241509",x"241509",x"1f1309",x"191008",x"1b1108",x"201308",x"1d1108",x"231409",x"221409",x"251509",x"1c1108",x"211309",x"1c1108",x"201309",x"201309",x"1b1108",x"231409",x"211309",x"201309",x"201309",x"1c1108",x"1d1108",x"1e1208",x"241509",x"241509",x"221409",x"1c1108",x"1d1208",x"1e1208",x"1c1108",x"170f07",x"170f07",x"1e1208",x"1b1108",x"1e1208",x"211309",x"1c1108",x"211309",x"1d1208",x"1b1108",x"1d1108",x"1b1008",x"1d1108",x"1b1008",x"1b1008",x"1d1108",x"1b1008",x"1d1108",x"1e1308",x"29180a",x"2a1a0a",x"2c1b0a",x"291a09",x"2a1909",x"291909",x"271809",x"1f1208",x"160e07",x"170f07",x"1a1008",x"1b1008",x"1b1008",x"180f07",x"191008",x"1a1008",x"1d1108",x"1b1108",x"1f1309",x"150e07",x"1f1309",x"1f1309",x"211409",x"1c1108",x"211309",x"1a1008",x"1d1108",x"1e1208",x"211309",x"211309",x"1c1108",x"221409",x"241509",x"1f1209",x"211409",x"25160a",x"25160a",x"231509",x"241509",x"24150a",x"24150a",x"1d1208",x"211309",x"221409",x"27170a",x"231509",x"150e07",x"150e07",x"160f07",x"170f07",x"180f08",x"191008",x"150e07",x"150e07",x"422510",x"412410",x"301b0b",x"28170a",x"2d190b",x"2c180a",x"2b180a",x"2b180a",x"29170a",x"2a170a",x"29170a",x"2d190b",x"261509",x"29180a",x"2a170a",x"28170a",x"2a180b",x"2a180a",x"2d190b",x"2c190b",x"2c180b",x"2f1a0b",x"301b0c",x"301b0c",x"2f1b0c",x"311c0c",x"2d190b",x"2e1a0b",x"2a180a",x"2c190a",x"2c180a",x"29170a",x"2e190b",x"301b0b",x"301a0b",x"2d190b",x"2c180b",x"301b0b",x"301b0b",x"301a0b",x"2d190b",x"2c190b",x"2a170a",x"281609",x"281609",x"2b180a",x"27160a",x"2b180b",x"2a170a",x"261509",x"241409",x"1f1108",x"1d1007",x"1f1007",x"1d0f06",x"1d0f07",x"1d0f07",x"1f1107",x"261509",x"28160a",x"261509",x"271509",x"2a170a",x"2b180b",x"2d1a0b",x"2c190b",x"27160a",x"2a180b",x"2b190b",x"29180b",x"28170a",x"29180b",x"29170a",x"2d1a0b",x"29170a",x"26160a",x"231409",x"241509",x"2d190b",x"321c0c",x"3c210f",x"3c210f",x"2d1a0c",x"2d1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1208",x"231409",x"211309",x"211308",x"211309",x"211309",x"211309",x"211309",x"211309",x"231509",x"231509",x"24150a",x"24150a",x"24150a",x"24150a",x"180e07",x"1a0f07",x"1e0f06",x"2b170a",x"281609",x"1b1008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"4b2b13",x"41250f",x"2f1c0b",x"25160a",x"201309",x"201309",x"211409",x"23150a",x"231509",x"1f1208",x"1f1208",x"201208",x"201309",x"211309",x"412510",x"25160a",x"23150a",x"23150a",x"23150a",x"29190a",x"28190a",x"41250f",x"1b1008",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"191008",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"170e07",x"190f07",x"1a1007",x"1e1408",x"191007",x"221508",x"231608",x"261809",x"33200b",x"291a09",x"2a1a09",x"2f1d0a",x"291909",x"281809",x"2a1a09",x"2c1b0a",x"261809",x"251709",x"261709",x"40250f",x"3c220e",x"40250f",x"3c220e",x"4f2d14",x"553315",x"241509",x"1a1008",x"191008",x"1d1207",x"1a110a",x"1a110a",x"1b1209",x"1d120a",x"1d130a",x"1d130a",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"1a1008",x"190f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"593415",x"42260b",x"47290e",x"43270e",x"3c240c",x"41230f",x"361e0d",x"351d0c",x"2a190a",x"201508",x"201408",x"211508",x"221608",x"201508",x"1b1108",x"190f07",x"170f07",x"170f07",x"20170f",x"432610",x"371f0e",x"472711",x"563117",x"4e2c14",x"472611",x"492812",x"4b2a14",x"533017",x"432612",x"4c2b15",x"432511",x"43250f",x"462610",x"4a2812",x"472811",x"432510",x"492912",x"43240f",x"4e2c13",x"4f2d13",x"553213",x"4f2d14",x"502d14",x"4f2e14",x"492911",x"371f0f",x"1b1108",x"361f0f",x"25160c",x"25160c"),
(x"150e07",x"150e07",x"150e07",x"28170a",x"3c210e",x"150e07",x"211409",x"2b190b",x"2a180b",x"2f1c0c",x"371f0e",x"301c0c",x"381f0e",x"351e0e",x"361f0e",x"3a210f",x"3a2210",x"331c0d",x"341d0d",x"39200e",x"361e0d",x"371f0e",x"351d0c",x"38200e",x"361e0d",x"331c0c",x"341d0d",x"351e0d",x"381f0d",x"311b0c",x"311c0c",x"331d0c",x"381f0e",x"341d0d",x"351e0d",x"381f0e",x"371f0e",x"331c0c",x"361e0d",x"391f0e",x"331c0c",x"371e0d",x"351d0d",x"341d0d",x"2f190b",x"331c0c",x"361f0e",x"321b0b",x"331c0b",x"331c0b",x"2f1a0b",x"371e0d",x"351c0c",x"3b210f",x"351e0d",x"38200e",x"38200e",x"39200f",x"3b220f",x"3b210f",x"3e230f",x"361d0d",x"301a0b",x"3a200e",x"381f0e",x"150e07",x"2d190b",x"2f1a0b",x"2f1b0c",x"27160a",x"371e0d",x"37210f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341d0c",x"482912",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1408",x"1f1408",x"221508",x"251809",x"271909",x"241708",x"241708",x"201508",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f08",x"191008",x"150e07",x"150e07",x"452711",x"412510",x"3f2310",x"412310",x"412410",x"402410",x"4d3729",x"594436",x"564132",x"402310",x"3f230f",x"3c210e",x"3a210f",x"3f2310",x"402410",x"3e2310",x"422611",x"3a200e",x"371d0d",x"3b200e",x"402310",x"432611",x"432611",x"3f230f",x"442611",x"452712",x"432611",x"422510",x"40230f",x"452711",x"462812",x"452611",x"442610",x"432510",x"432510",x"452711",x"432611",x"442611",x"432510",x"432511",x"422410",x"452711",x"442611",x"3f230f",x"3b200e",x"3a1f0d",x"3c200e",x"41230f",x"3c210e",x"3b200e",x"3e220f",x"3e210e",x"40230f",x"422410",x"422410",x"422410",x"432510",x"43240f",x"42240f",x"432510",x"432510",x"43240f",x"3e210e",x"3c200e",x"3d210e",x"3c210e",x"3f220f",x"40230f",x"3c200e",x"3e220e",x"3e210f",x"412510",x"442611",x"452813",x"452813",x"412611",x"3d2310",x"3b210f",x"3d210e",x"422511",x"432611",x"452812",x"432511",x"432511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231409",x"211309",x"211308",x"211309",x"211309",x"211309",x"211309",x"211309",x"231509",x"231509",x"24150a",x"24150a",x"24150a",x"1f1208",x"201309",x"211409",x"211309",x"211409",x"211409",x"211409",x"211409",x"211409",x"201309",x"1f1208",x"1e1208",x"201208",x"472712",x"371f0c",x"231508",x"231409",x"211309",x"211308",x"1f1208",x"231509",x"231509",x"201309",x"211409",x"211309",x"25160a",x"211409",x"211409",x"221509",x"231509",x"25160a",x"251609",x"28180a",x"29180a",x"452812",x"1d1108",x"1d1108",x"1c1108",x"1b1108",x"211309",x"211409",x"1c1108",x"2b180b",x"22150b",x"32251c",x"170f07",x"160f07",x"381f0e",x"39200d",x"371f0d",x"472911",x"37200c",x"3a210d",x"3f2510",x"442810",x"40270f",x"3a220d",x"351f0b",x"321d0a",x"301b0b",x"28170a",x"261609",x"28180a",x"2f1c0c",x"2c1b0a",x"28180a",x"29190a",x"29190a",x"41260f",x"3a210e",x"452810",x"573315",x"512f15",x"1c1108",x"1a1008",x"1a1008",x"191008",x"1a1008",x"1a110a",x"1a1109",x"1d120a",x"1c120b",x"1d120b",x"1d130a",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1a1008",x"1a1008",x"180f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"191007",x"512e12",x"502f13",x"3f260d",x"2b190b",x"2c190b",x"1b1108",x"1c1208",x"221509",x"1e1408",x"2b190a",x"221608",x"231608",x"1c1208",x"1b1108",x"1b1107",x"160e07",x"170f07",x"170f07",x"180f08",x"3c220f",x"2e190b",x"2c180b",x"2d190b",x"2d190b",x"321c0e",x"331d0e",x"351e0f",x"331c0e",x"351d0e",x"381f0f",x"3d2210",x"391f0e",x"371e0e",x"40230f",x"3f230f",x"3e220f",x"452711",x"492911",x"472911",x"42240f",x"40230f",x"40240e",x"4c2811",x"442811",x"1a1008",x"1a1008",x"362920",x"362920",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"3b200e",x"150e07",x"150e07",x"3e220f",x"341d0d",x"351d0d",x"331d0d",x"371e0e",x"381f0e",x"351d0d",x"321c0c",x"321c0d",x"2e1a0b",x"2c190b",x"28170a",x"351e0d",x"341d0d",x"331d0d",x"301b0c",x"301a0b",x"2c180b",x"2d1a0b",x"341d0d",x"2e190b",x"2d190b",x"2c180b",x"301b0c",x"2e1a0b",x"2d190b",x"2c190b",x"2d190b",x"331c0c",x"331c0c",x"361e0d",x"351d0d",x"331c0d",x"321c0c",x"331c0d",x"341d0d",x"331c0c",x"2f1b0c",x"321b0c",x"331d0d",x"321d0d",x"341d0d",x"341d0d",x"38200e",x"311c0c",x"341d0d",x"301b0b",x"2f190b",x"2e180a",x"2e180a",x"2f1a0b",x"331c0c",x"331c0c",x"341c0c",x"361d0c",x"3c210e",x"381f0d",x"381f0d",x"301a0b",x"371d0c",x"29170a",x"311b0c",x"150e07",x"331b0b",x"39200f",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b200e",x"442610",x"3e220f",x"371e0c",x"341c0c",x"351c0c",x"321b0b",x"3c210f",x"3d210f",x"3f2310",x"412410",x"422510",x"3e2310",x"412511",x"442611",x"3b200e",x"3a200e",x"3a200e",x"3b210e",x"3d220f",x"3e220f",x"3e230f",x"3d220f",x"3a200e",x"391f0e",x"39200e",x"3a200e",x"3e2310",x"432611",x"3b210f",x"3a200d",x"3b200e",x"3e230f",x"3d220f",x"3d210f",x"381e0c",x"381f0d",x"3b210e",x"3a200e",x"3b200e",x"3e220e",x"3d210f",x"3b210e",x"3d220f",x"3a200e",x"3d230f",x"422510",x"422510",x"3c210f",x"3b210e",x"3a200e",x"3a200e",x"3d220f",x"3d220f",x"432711",x"3e240f",x"3e230f",x"3b220e",x"371f0c",x"422610",x"3b200d",x"42250f",x"3c220d",x"3a200c",x"361e0b",x"39200c",x"361d0c",x"3a200d",x"351d0c",x"361e0d",x"3b200e",x"381f0d",x"381f0d",x"361d0c",x"381e0c",x"371e0d",x"3a200d",x"391f0d",x"371d0c",x"391f0e",x"361d0c",x"2e180a",x"321b0b",x"341c0c",x"3a200e",x"39200e",x"3b210e",x"3d210f",x"3d210e",x"371d0c",x"391f0d",x"391f0e",x"3d210f",x"3d210f",x"3f220f",x"432510",x"3f240f",x"412410",x"3e230f",x"482812",x"170f07",x"898989",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2310",x"422510",x"412410",x"402410",x"4d3729",x"594436",x"564132",x"402310",x"3f230f",x"3c210e",x"3a210f",x"3f2310",x"402410",x"3e2310",x"422611",x"3a200e",x"371d0d",x"3b200e",x"402310",x"432611",x"432611",x"41240f",x"442611",x"452712",x"432611",x"422510",x"40230f",x"452711",x"462812",x"452611",x"442610",x"432510",x"432510",x"452711",x"432611",x"442611",x"432510",x"432511",x"422410",x"452711",x"442611",x"3f230f",x"3b200e",x"3a1f0d",x"3c200e",x"41230f",x"3c210e",x"3b200e",x"3f220e",x"3e210e",x"40230f",x"422410",x"422410",x"422410",x"432510",x"43240f",x"42240f",x"432510",x"432510",x"43240f",x"3e210e",x"3c200e",x"3d210e",x"3c210e",x"3f220f",x"40230f",x"3c200e",x"3e220e",x"3e210f",x"412510",x"442611",x"452813",x"452813",x"412611",x"3d2310",x"3b210f",x"3d210e",x"422511",x"432611",x"452812",x"482913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1108",x"1e1108",x"1f1208",x"1f1208",x"1e1108",x"1e1108",x"1f1208",x"211309",x"201308",x"201308",x"201208",x"201309",x"27160a",x"3c210f",x"432811",x"3a230e",x"38200e",x"351f0d",x"2d1b0b",x"2e1c0a",x"271909",x"201308",x"1d1108",x"1d1108",x"1e1108",x"1f1208",x"201309",x"221408",x"231509",x"251609",x"281609",x"28170a",x"331d0b",x"2d1b0b",x"2f1b0b",x"28180a",x"271709",x"27160a",x"27190d",x"191008",x"191008",x"1e1208",x"39200e",x"33261c",x"352c24",x"4a392d",x"3b210f",x"3b210f",x"3a210d",x"291809",x"2d1b0a",x"36210c",x"35200b",x"36200c",x"36210c",x"37210d",x"3a220d",x"351e0d",x"3b230e",x"301b0b",x"28170a",x"2d1a0b",x"28180a",x"2f1c0c",x"2b190b",x"28180a",x"29190a",x"39220e",x"3a220e",x"492a12",x"4a2a12",x"5e3617",x"533115",x"1c1108",x"221608",x"211508",x"1f1408",x"39200e",x"26160a",x"261509",x"2e190b",x"26160a",x"27160a",x"231509",x"231509",x"1d1108",x"1d1108",x"3a2210",x"331d0d",x"24160a",x"26170a",x"261709",x"180f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1207",x"1c1207",x"1c1107",x"1a1007",x"1b1008",x"1c1107",x"4e2d11",x"231509",x"1f1309",x"160f07",x"160e07",x"181007",x"1d1308",x"221608",x"211508",x"251508",x"1e1308",x"1c1208",x"181007",x"170f07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f07",x"190f07",x"221409",x"201208",x"22150b",x"27180c",x"27180c",x"24160b",x"2a190c",x"2a190c",x"2c1a0c",x"2f1b0d",x"311c0d",x"381f0f",x"392010",x"3d2211",x"412512",x"442711",x"422610",x"41250f",x"3c220f",x"432710",x"40240f",x"442610",x"3e240f",x"1a1008",x"191008",x"351d0d",x"351d0d",x"000000"),
(x"150e07",x"150e07",x"150e07",x"251509",x"3c220f",x"2c190b",x"211409",x"432611",x"26160a",x"462813",x"432713",x"412511",x"3d2210",x"37200e",x"3b210f",x"341d0d",x"341d0d",x"361f0e",x"37200e",x"3b210f",x"3c210f",x"3c210f",x"38200e",x"39200e",x"3f2410",x"3e230f",x"3a210f",x"3a200e",x"371f0d",x"381f0e",x"381f0e",x"341d0c",x"361e0d",x"351d0d",x"361d0d",x"351d0d",x"351d0c",x"341c0c",x"341c0c",x"321c0c",x"301b0b",x"311b0b",x"341c0c",x"371f0e",x"38200f",x"3d220f",x"3d220f",x"3b210e",x"361e0c",x"3d220e",x"331c0b",x"3b210f",x"321b0b",x"341c0c",x"341c0b",x"2e170a",x"2e1709",x"2f180a",x"2f180a",x"2b1609",x"30190a",x"351c0c",x"331b0b",x"351c0c",x"331b0b",x"1f1208",x"391f0d",x"150e07",x"2d190b",x"150e07",x"2e180a",x"341c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39200d",x"39200d",x"351d0c",x"3b210e",x"351e0c",x"331c0c",x"2e1a0b",x"311b0c",x"2f1b0c",x"2d190b",x"361f0e",x"361f0e",x"321c0c",x"331d0d",x"351f0e",x"38200e",x"341d0d",x"331d0d",x"331d0d",x"37200f",x"351e0e",x"331d0d",x"321c0d",x"2f1b0c",x"301b0c",x"2e1a0b",x"311c0c",x"341d0d",x"2f1b0c",x"301b0c",x"2e1a0c",x"2d1a0b",x"2b180b",x"28160a",x"29170a",x"2a170a",x"2c190b",x"301a0b",x"2f1a0b",x"28160a",x"29170a",x"27160a",x"261509",x"241509",x"251509",x"211309",x"231409",x"271709",x"2b180a",x"2c190a",x"271609",x"2a180a",x"2c190a",x"2e1b0a",x"2d1a0a",x"29180a",x"251509",x"2a180a",x"2c1a0a",x"2e1b0b",x"301c0b",x"321c0b",x"2f1b0b",x"2e1b0b",x"301c0c",x"2f1b0b",x"2e1a0b",x"2b190b",x"2c190b",x"2c190b",x"2a180b",x"29170a",x"27160a",x"27160a",x"29180b",x"28170a",x"28170a",x"2b190b",x"2b190b",x"27160a",x"301c0c",x"301c0d",x"2e1b0b",x"2b190b",x"27170b",x"29180b",x"25160a",x"28170a",x"2d1a0c",x"301c0d",x"351f0e",x"36200f",x"37200f",x"351f0e",x"452813",x"422612",x"3c2210",x"3d2310",x"402511",x"422611",x"3a210f",x"3e220f",x"3e220f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1209",x"1e1209",x"1f1309",x"1e1208",x"1c1108",x"1b1108",x"1b1008",x"1b1108",x"1f1209",x"211509",x"231509",x"2a1a0a",x"261809",x"251708",x"231608",x"1e1108",x"1f1208",x"1f1208",x"1f1208",x"1f1108",x"1f1108",x"1f1208",x"1f1208",x"1d1108",x"1e1108",x"1e1108",x"1a1108",x"432810",x"432811",x"351f0c",x"331f0b",x"2d1b0a",x"281809",x"271709",x"2a1a09",x"1b1108",x"201308",x"201309",x"201309",x"211309",x"201309",x"211309",x"201309",x"201309",x"26170a",x"26170a",x"27180a",x"25160a",x"29180a",x"2a180a",x"331c0c",x"321c0c",x"3d2f25",x"1d150e",x"1b110b",x"351e0e",x"26160a",x"3f362d",x"40362c",x"463b32",x"534135",x"361f0d",x"29180a",x"2f1c0b",x"321d0b",x"2e1b0a",x"35200c",x"39230d",x"36210b",x"35200c",x"311d0b",x"2b1a0b",x"2b1a0b",x"2c1a0b",x"28170a",x"28160a",x"2c1a0b",x"26160a",x"27180a",x"2a190a",x"27170a",x"2f1c0a",x"3a220e",x"4a2a12",x"452811",x"522f15",x"1d1208",x"1a1107",x"251609",x"472911",x"3c220e",x"341d0d",x"39200e",x"361e0d",x"3d200e",x"211309",x"201309",x"201308",x"2d190b",x"23140a",x"221409",x"24150a",x"1d1108",x"1c1108",x"1c1108",x"29190a",x"29180a",x"231409",x"1b1107",x"1d1208",x"211508",x"1a1108",x"1c1308",x"1e1308",x"1c1208",x"1d1208",x"201408",x"1d1208",x"211509",x"221509",x"251c14",x"261e16",x"150e07",x"150e07",x"160e07",x"1a1107",x"221508",x"1e1308",x"1d1308",x"221508",x"29170a",x"2d1b0c",x"1c1208",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"191008",x"180f07",x"1d1208",x"20140b",x"20140b",x"21150b",x"23160b",x"26170b",x"2d1b0d",x"311c0e",x"2f1b0d",x"2e1b0d",x"331d0e",x"38200f",x"39200f",x"3d2211",x"412611",x"402412",x"432611",x"442712",x"4a2b12",x"422610",x"4f2d14",x"39200d",x"1f1309",x"1b1008",x"27160a",x"27160a",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231409",x"341c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"150e07",x"2c170a",x"301a0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b210f",x"351d0d",x"4c2b14",x"432612",x"462812",x"3f2310",x"402410",x"412511",x"432712",x"482a14",x"432712",x"402410",x"3f230f",x"3e220f",x"402410",x"412410",x"3e230f",x"3f230f",x"422510",x"3f2410",x"452812",x"412511",x"3e2411",x"412511",x"422612",x"432611",x"402310",x"452712",x"422611",x"412511",x"452712",x"432611",x"3d230f",x"412511",x"412511",x"3f2310",x"3d220f",x"422611",x"412511",x"402511",x"432611",x"482a14",x"442611",x"472a14",x"462813",x"3d2310",x"3b220e",x"422711",x"462912",x"452912",x"3e240d",x"412711",x"462911",x"46280f",x"43270f",x"3c220c",x"3e230d",x"43260f",x"40240e",x"402510",x"412510",x"41240f",x"3f250f",x"43260f",x"3c220e",x"3a200e",x"371e0d",x"351c0c",x"341c0c",x"331c0c",x"331c0c",x"301a0b",x"351c0c",x"351c0b",x"381e0d",x"361e0d",x"371e0d",x"3b200e",x"3c210f",x"412410",x"3d220f",x"3e2310",x"3e220f",x"3c220f",x"3f2310",x"3d220f",x"3b200e",x"3d220f",x"412411",x"432611",x"402411",x"3e2310",x"402411",x"422511",x"412511",x"402411",x"412411",x"432611",x"402410",x"482912",x"1d1208",x"29170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1209",x"1e1209",x"1f1309",x"1e1208",x"1c1108",x"1b1108",x"1b1008",x"1b1108",x"1f1209",x"211509",x"231509",x"2a1a0a",x"261809",x"251708",x"231608",x"211509",x"201408",x"1f1408",x"29180a",x"2f1c0b",x"2f1b0b",x"2e1a0b",x"29190a",x"231608",x"28190a",x"442a0f",x"37230b",x"321f0a",x"311f0a",x"311f0a",x"301e0a",x"271809",x"241708",x"2b1b09",x"221608",x"361f0d",x"211309",x"211409",x"211309",x"211409",x"211309",x"201309",x"211409",x"201309",x"251509",x"251609",x"241609",x"211409",x"27170a",x"2a180b",x"321b0d",x"351e0e",x"43362d",x"29211a",x"221a13",x"3c200e",x"29190e",x"3c3229",x"453b32",x"4c4137",x"4e4339",x"371f0e",x"28170a",x"29180b",x"2c1a0b",x"341f0c",x"38220d",x"3a230d",x"38220c",x"341f0c",x"301d0b",x"2f1c0b",x"2a190b",x"2c1a0b",x"29180a",x"251609",x"251509",x"26160a",x"26160a",x"29190a",x"29190a",x"27180a",x"171007",x"1a1107",x"1a1107",x"191007",x"4b2c14",x"442812",x"3a210f",x"3d2410",x"37200e",x"3b220f",x"3b220f",x"301b0c",x"180f07",x"221409",x"231509",x"221409",x"221409",x"24150a",x"221409",x"1f1208",x"1f1309",x"1f1309",x"201309",x"241509",x"29190b",x"1b1107",x"1b1107",x"1d1308",x"221608",x"221508",x"221508",x"231708",x"291a09",x"231608",x"271808",x"201309",x"201409",x"1f1308",x"2e241a",x"22160d",x"150e07",x"150e07",x"150e07",x"1b1108",x"221608",x"1e1308",x"221608",x"211508",x"1e1408",x"211509",x"2a180b",x"2c190b",x"160e07",x"160f07",x"170f07",x"180f07",x"191008",x"180f07",x"34210b",x"40260f",x"452a11",x"20140b",x"21150b",x"27170c",x"22150b",x"2a190d",x"311d0e",x"321d0f",x"372010",x"361f10",x"3d2311",x"3d2312",x"3f2412",x"412513",x"3f2412",x"432711",x"482a13",x"432612",x"492b13",x"4b2b13",x"422813",x"1d1208",x"1c1108",x"211408",x"211408",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211309",x"2d190b",x"301a0b",x"341d0d",x"371f0e",x"3b2210",x"3c2310",x"3d2310",x"3d2310",x"3b220f",x"351e0e",x"2f1a0b",x"3b210f",x"321c0d",x"361f0e",x"39200e",x"3d2310",x"331d0d",x"39200f",x"351e0d",x"3d2310",x"3c2310",x"38200f",x"3a2210",x"351e0e",x"371f0e",x"3d2310",x"38200f",x"3c2311",x"3a210f",x"3d2310",x"432713",x"3f2411",x"39200f",x"3f2512",x"402511",x"3e2411",x"3e2411",x"3b2210",x"351e0d",x"3d2310",x"361d0d",x"341c0b",x"311b0b",x"3b210e",x"3b200e",x"381e0c",x"361d0c",x"3b210f",x"311c0c",x"341d0d",x"321c0c",x"341d0c",x"351d0d",x"3a200f",x"3b200f",x"331c0c",x"301a0b",x"341c0c",x"2a1509",x"281408",x"281408",x"251308",x"261308",x"241308",x"2f180a",x"321b0c",x"301a0b",x"2c190a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200e",x"321c0c",x"472912",x"4b2a13",x"462712",x"4c2a13",x"472812",x"462711",x"4a2913",x"4b2a13",x"4d2c14",x"4a2912",x"4e2c14",x"4e2d14",x"4d2b14",x"4f2d15",x"4d2b13",x"4b2a13",x"482711",x"492912",x"4d2b14",x"4b2a13",x"4c2b13",x"482812",x"4a2a13",x"442410",x"42240f",x"462711",x"4a2913",x"472711",x"42240f",x"43240f",x"41230f",x"41220e",x"44250f",x"41230e",x"42240f",x"3f200e",x"3d200d",x"452610",x"432510",x"42240f",x"442510",x"3e220f",x"41230f",x"43240f",x"44260f",x"482910",x"4b2b12",x"482911",x"472810",x"45270f",x"472810",x"4a2a10",x"44260f",x"46280f",x"46280f",x"482910",x"492911",x"4b2a12",x"492911",x"4b2a12",x"4f2d13",x"4d2d14",x"4c2b13",x"442611",x"462711",x"412410",x"432611",x"472812",x"452611",x"391f0d",x"3d210e",x"3b200d",x"3a1f0d",x"3d210e",x"3b1f0d",x"391f0c",x"3c1f0d",x"3c1f0c",x"3b1f0c",x"3b1e0c",x"3c200d",x"42240f",x"40230e",x"3d210e",x"462611",x"482812",x"462711",x"482811",x"4b2b13",x"492912",x"482812",x"4a2913",x"4a2a13",x"4a2913",x"492812",x"462611",x"462711",x"331c0c",x"180f08",x"1c1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1208",x"1d1208",x"211509",x"26170a",x"201409",x"241509",x"1f1309",x"1e1208",x"1e1208",x"241508",x"2c190b",x"301c0a",x"27170a",x"2c1a0b",x"2f1a0b",x"331d0c",x"311c0b",x"311b0b",x"331d0b",x"37200d",x"351f0d",x"331d0e",x"201408",x"1c1107",x"3e270e",x"37230b",x"3a250b",x"33200a",x"34210b",x"35210b",x"2f1e0a",x"281909",x"241708",x"271909",x"291a09",x"221608",x"201309",x"27160a",x"29170a",x"28170a",x"29160a",x"2d1a0b",x"311c0c",x"2e1b0b",x"311c0c",x"331e0c",x"331d0c",x"361e0d",x"39200d",x"3d2210",x"492a13",x"452812",x"504135",x"3e3127",x"302720",x"1c1108",x"301b0c",x"38271c",x"352c23",x"3b3027",x"382e25",x"1f1309",x"2c190a",x"29180a",x"321e0b",x"301c0a",x"311e0b",x"331f0b",x"311d0b",x"321e0b",x"2c1a0a",x"2c1a0a",x"29180a",x"2e1b0b",x"29180a",x"29180a",x"28180a",x"26160a",x"251609",x"27170a",x"28180a",x"1b1108",x"1a1107",x"311c0c",x"492912",x"3c2310",x"38210e",x"3a210e",x"3c220f",x"422711",x"422611",x"361f0e",x"211409",x"231509",x"211409",x"150e07",x"231509",x"221409",x"221409",x"24150a",x"24150a",x"160e07",x"170e07",x"160f07",x"170f07",x"180f07",x"1b1107",x"201408",x"1e1308",x"221508",x"241608",x"271809",x"241608",x"281909",x"261808",x"221508",x"261809",x"261709",x"221509",x"1f1308",x"291d14",x"1e1208",x"2c1b0a",x"150e07",x"150e07",x"181007",x"1b1108",x"1c1208",x"251809",x"281a09",x"1d1208",x"1e1308",x"1c1208",x"29170a",x"27160a",x"160e07",x"170f07",x"170f07",x"211509",x"261809",x"311f0b",x"3b240d",x"432811",x"1e130b",x"23150b",x"24150c",x"1d130a",x"20140b",x"28180c",x"27180c",x"2c1a0d",x"321d0e",x"392111",x"3f2512",x"432613",x"402412",x"3c2211",x"462913",x"432812",x"472b13",x"432811",x"482a13",x"3d230f",x"1c1108",x"251609",x"201308",x"1f1208",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1a1008",x"241409",x"28160a",x"2f1a0b",x"2d190b",x"2a170a",x"311c0c",x"311c0c",x"341d0d",x"2a180a",x"2c180b",x"311b0c",x"321c0c",x"29180b",x"2a180b",x"331d0d",x"351e0e",x"331d0d",x"311c0d",x"2f1b0c",x"351e0e",x"361f0e",x"311c0d",x"39210f",x"37200f",x"301b0c",x"341d0d",x"331c0d",x"351e0e",x"311c0c",x"39200f",x"392110",x"39200f",x"37200e",x"36200f",x"321c0d",x"381f0e",x"351e0d",x"351f0e",x"311c0c",x"2f1a0b",x"2f1a0a",x"2e190a",x"2e1a0b",x"2b170a",x"351d0c",x"271509",x"2f1a0b",x"321c0c",x"311c0d",x"331d0d",x"321c0d",x"351f0e",x"321c0d",x"331d0d",x"38200e",x"331c0d",x"331c0c",x"2f1a0c",x"301b0c",x"351d0d",x"341d0d",x"361f0e",x"351e0e",x"331d0d",x"331d0d",x"361f0e",x"331d0e",x"221409",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c210f",x"472912",x"4b2a13",x"462712",x"4c2a13",x"472812",x"462711",x"4a2913",x"4b2a13",x"4d2c14",x"4a2912",x"4e2c14",x"4e2d14",x"4d2b14",x"4f2d15",x"4d2b13",x"4b2a13",x"482711",x"492912",x"4d2b14",x"4b2a13",x"4c2b13",x"482812",x"4a2a13",x"442410",x"42240f",x"462711",x"4a2913",x"472711",x"42240f",x"43240f",x"41230f",x"41220e",x"44250f",x"41230e",x"42240f",x"3f200e",x"3d200d",x"452610",x"432510",x"42240f",x"442510",x"3e220f",x"41230f",x"43240f",x"44260f",x"482910",x"4b2b12",x"482911",x"472810",x"45270f",x"472810",x"4a2a10",x"44260f",x"46280f",x"46280f",x"482910",x"492911",x"4b2a12",x"492911",x"4b2a12",x"4f2d13",x"4d2d14",x"4c2b13",x"442611",x"462711",x"412410",x"432611",x"472812",x"452611",x"391f0d",x"3d210e",x"3b200d",x"3a1f0d",x"3d210e",x"3b1f0d",x"391f0c",x"3c1f0d",x"3c1f0c",x"3b1f0c",x"3b1e0c",x"3c200d",x"42240f",x"40230e",x"3d210e",x"462611",x"482812",x"462711",x"482811",x"4b2b13",x"492912",x"482812",x"4a2913",x"4a2a13",x"4a2913",x"492812",x"462611",x"462711",x"331c0c",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1308",x"1e1308",x"1d1208",x"1e1208",x"1f1309",x"201309",x"1e1208",x"211309",x"201308",x"28180a",x"241609",x"26170a",x"271709",x"291809",x"2b1a0a",x"2d1b0b",x"301d0b",x"2a190b",x"2f1c0c",x"2f1c0b",x"361e0d",x"312113",x"20150c",x"1b1008",x"311f0b",x"33200a",x"37230b",x"37230b",x"301f0a",x"2b1b09",x"251809",x"1d1308",x"1e1308",x"241708",x"191007",x"211508",x"301c0d",x"26170a",x"29180b",x"2d1a0c",x"2d1a0b",x"2e1a0b",x"2e1b0b",x"301d0c",x"2f1c0b",x"2f1c0b",x"321d0c",x"38200d",x"3b220e",x"402510",x"482a12",x"442811",x"4e3f34",x"2e251d",x"211912",x"22150a",x"3e2310",x"2d1a0b",x"21150a",x"1f1208",x"2d1a0c",x"2d1a0c",x"27170a",x"27170a",x"2d1b0a",x"311e0b",x"35200b",x"341f0c",x"331f0b",x"301d0b",x"41270f",x"43280f",x"42270f",x"3f240f",x"2b190b",x"27170a",x"29180a",x"27170a",x"191007",x"191007",x"180f07",x"4a2a12",x"3d230f",x"3a220e",x"38200e",x"3e2310",x"402510",x"412510",x"432610",x"39200e",x"341d0d",x"2d1a0c",x"211409",x"351f0e",x"221409",x"1c1108",x"181007",x"180f07",x"170f07",x"1e1308",x"170f07",x"170f07",x"170f07",x"160f07",x"170f07",x"1b1107",x"1f1309",x"201409",x"241608",x"291909",x"38210d",x"43260e",x"34200c",x"36200b",x"38210d",x"3f2310",x"2b190b",x"3c230f",x"3d230f",x"3d240f",x"2b1f14",x"23160a",x"25160a",x"150e07",x"150e07",x"150e07",x"191007",x"1a1107",x"1d1208",x"1f1408",x"1a1107",x"1a1107",x"1c1207",x"1a1107",x"27160a",x"201309",x"170f07",x"1e1208",x"1d1208",x"241609",x"2e1c0a",x"3b240d",x"452913",x"452913",x"23150b",x"23150b",x"20140b",x"1e140b",x"17110a",x"25170b",x"24170b",x"2f1c0d",x"382010",x"3b2211",x"402513",x"412712",x"432713",x"462914",x"432712",x"442713",x"432911",x"462912",x"3a220f",x"241509",x"381e0b",x"1f1208",x"1f1209",x"1f1209"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"201308",x"2f1a0b",x"39200e",x"361d0d",x"3b210f",x"361e0d",x"381f0e",x"331d0d",x"311c0c",x"2f1b0c",x"241509",x"150e07",x"24150a",x"1a1008",x"1a1008",x"201309",x"1d1108",x"1b1108",x"150e07",x"2d1a0c",x"2e1b0c",x"331d0e",x"331d0e",x"361f0f",x"3d2411",x"3d2410",x"3c2310",x"3e2310",x"3a2110",x"361f0f",x"351f0e",x"351e0e",x"351f0e",x"25160a",x"1b1108",x"1b1108",x"170f07",x"241509",x"231409",x"170f07",x"150e07",x"251509",x"201208",x"1f1208",x"241509",x"29170a",x"2c190b",x"2f1b0c",x"301b0c",x"331d0d",x"321c0c",x"321c0c",x"341c0c",x"371f0e",x"3c220f",x"3b210f",x"351d0d",x"351d0d",x"341d0c",x"3d220f",x"3c230f",x"3f2410",x"3d230f",x"3b220f",x"2f1b0c",x"27170a",x"150e07",x"150e07",x"150e07",x"443226",x"3b210f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"54463a",x"442711",x"442511",x"442510",x"512e16",x"6e4b30",x"68452b",x"67452b",x"6f4d32",x"6e4c30",x"614129",x"634229",x"66442a",x"624128",x"63422a",x"62432a",x"704e32",x"614229",x"614229",x"6e4d32",x"6e4d32",x"63432a",x"67452b",x"6d4c30",x"6d4b30",x"64442b",x"66452c",x"745337",x"745236",x"65452d",x"64442c",x"77563a",x"76553a",x"6a4a30",x"68482e",x"7a593c",x"6c4c32",x"6d4e35",x"6b4c32",x"78573b",x"66462d",x"6b4b30",x"7a583b",x"7c5a3d",x"6a4b32",x"6a4a31",x"7b583b",x"7c593c",x"694a31",x"6a492f",x"78563a",x"775437",x"68482e",x"65452d",x"725035",x"6d4c32",x"614128",x"5e3f27",x"69482f",x"67482e",x"604129",x"5f4028",x"6b4b31",x"5c3e26",x"5f4128",x"604028",x"63422a",x"5f4027",x"634329",x"725035",x"69492f",x"614128",x"614229",x"6a492f",x"6f4d32",x"614128",x"66442a",x"6e4c30",x"6f4c30",x"69472d",x"6c492e",x"775538",x"775437",x"6c4a2f",x"6c492e",x"7d5a3c",x"7c583b",x"6e4d31",x"6c4a2f",x"7d5a3d",x"704e33",x"704f34",x"6f4e33",x"7c593b",x"5d4129",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1408",x"1f1408",x"1e1209",x"1f1309",x"1d1108",x"1e1108",x"201309",x"241409",x"231409",x"221308",x"251509",x"2a190a",x"2f1c0a",x"34200c",x"321e0b",x"331f0c",x"2e1b0b",x"28180a",x"29180a",x"28160a",x"331d0c",x"332318",x"35291f",x"3b250d",x"34210b",x"37230b",x"3d270c",x"3b250c",x"36220b",x"2e1d0a",x"2a1b09",x"281909",x"211508",x"1b1108",x"160f07",x"181007",x"231509",x"231409",x"25150a",x"27170a",x"27170a",x"2c1a0b",x"311d0b",x"301c0c",x"331f0c",x"341f0c",x"341f0c",x"341f0c",x"35200d",x"39200d",x"41250f",x"41250f",x"443428",x"201812",x"191008",x"3d2411",x"2f1c0d",x"221409",x"211409",x"211409",x"201209",x"351f0d",x"331d0c",x"28170b",x"301c0b",x"331d0c",x"38210d",x"36200c",x"38210b",x"38220c",x"36220b",x"36220b",x"38220d",x"3a210d",x"432711",x"381d0c",x"1d1208",x"150e07",x"3a200f",x"4b2c14",x"38200e",x"3b210e",x"3e230f",x"3c230f",x"422510",x"422610",x"3d240f",x"3c2210",x"37200e",x"361f0e",x"351f0e",x"2c1a0c",x"36200f",x"371f0f",x"3f230f",x"170f07",x"170f07",x"191007",x"180f07",x"1a1107",x"1d1208",x"170f07",x"1a1107",x"191007",x"190f08",x"251509",x"27180a",x"251609",x"261709",x"311d0b",x"2d1c0a",x"3d220f",x"371f0d",x"27160a",x"180f07",x"150e07",x"150e07",x"3f2510",x"3d230f",x"3d240f",x"38200e",x"251609",x"2d1b0a",x"2c1a0a",x"150e07",x"150e07",x"160e07",x"191007",x"181007",x"1a1107",x"1d1308",x"170f07",x"150e07",x"150e07",x"150e07",x"170e07",x"1f1209",x"1f1209",x"1e1209",x"1e1308",x"1d1208",x"2a190b",x"3d2311",x"211309",x"201309",x"28170a",x"301b0c",x"2b180b",x"1d130a",x"20140b",x"1f140b",x"28180c",x"2f1c0d",x"351e0f",x"341e0f",x"402512",x"402613",x"432712",x"3b2311",x"432611",x"492c13",x"502f17",x"3b220e",x"1d1208",x"1f1209",x"2f1b0c",x"452b19",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"190f07",x"241409",x"27160a",x"29170a",x"29160a",x"29170a",x"29170a",x"251509",x"231408",x"1e1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"27160a",x"25150a",x"2a180b",x"29180a",x"211309",x"1e1208",x"27160a",x"2a180a",x"3b200e",x"331d0c",x"28170a",x"301b0c",x"221409",x"25150a",x"1e1209",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"170f07",x"150e07",x"150e07",x"2d190b",x"241509",x"24150a",x"231509",x"221309",x"201308",x"211309",x"231409",x"201309",x"28160a",x"27160a",x"221308",x"241509",x"29160a",x"29170a",x"27160a",x"371f0d",x"39200e",x"3a200e",x"371e0d",x"2e1a0b",x"2d190b",x"170f08",x"160f07",x"38200e",x"1a1008",x"443226",x"3b210f",x"3b210f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"54463a",x"54463a",x"442711",x"442511",x"442510",x"512e16",x"6e4b30",x"68452b",x"67452b",x"6f4d32",x"6e4c30",x"614129",x"634229",x"66442a",x"624128",x"63422a",x"62432a",x"704e32",x"614229",x"614229",x"6e4d32",x"6e4d32",x"63432a",x"67452b",x"6d4c30",x"6d4b30",x"64442b",x"66452c",x"745337",x"745236",x"65452d",x"64442c",x"77563a",x"76553a",x"6a4a30",x"68482e",x"7a593c",x"6c4c32",x"6d4e35",x"6b4c32",x"78573b",x"66462d",x"6b4b30",x"7a583b",x"7c5a3d",x"6a4b32",x"6a4a31",x"7b583b",x"7c593c",x"694a31",x"6a492f",x"78563a",x"775437",x"68482e",x"65452d",x"725035",x"6d4c32",x"614128",x"5e3f27",x"69482f",x"67482e",x"604129",x"5f4028",x"6b4b31",x"5c3e26",x"5f4128",x"604028",x"63422a",x"5f4027",x"634329",x"725035",x"69492f",x"614128",x"614229",x"6a492f",x"6f4d32",x"614128",x"66442a",x"6e4c30",x"6f4c30",x"69472d",x"6c492e",x"775538",x"775437",x"6c4a2f",x"6c492e",x"7d5a3c",x"7c583b",x"6e4d31",x"6c4a2f",x"7d5a3d",x"704e33",x"704f34",x"6f4e33",x"7c593b",x"5d4129",x"5d4129",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"221409",x"331c0c",x"361f0e",x"301a0b",x"2e1a0b",x"2e190a",x"2b180a",x"331c0c",x"321c0b",x"361e0c",x"39210c",x"3d230d",x"3e250f",x"3b230d",x"41250e",x"3b210e",x"3d220e",x"432610",x"442510",x"3c200d",x"3e281b",x"4b3a2d",x"3f270e",x"38240b",x"3d270c",x"3e270c",x"37230b",x"35220b",x"2e1d0a",x"251708",x"1c1208",x"1f1408",x"1b1108",x"160f07",x"211409",x"25150a",x"221409",x"241509",x"251509",x"221309",x"271609",x"2e1b0b",x"28180b",x"2c1a0b",x"2c1a0b",x"35200d",x"341e0c",x"39220e",x"3f240f",x"462911",x"472913",x"452e20",x"1b120b",x"1a1008",x"1b1108",x"201309",x"28180a",x"28180a",x"251609",x"27170a",x"231409",x"251509",x"231509",x"24160a",x"2c1b0a",x"311e0b",x"311e0a",x"321e0a",x"34200b",x"2f1d0b",x"311e0b",x"2d1c0a",x"2c1a0a",x"241509",x"2e1a0b",x"39200e",x"351e0d",x"3f220d",x"40220e",x"3d210d",x"3c210e",x"3e210e",x"41240f",x"3d220e",x"371f0d",x"311c0b",x"321d0c",x"2d1a0b",x"241509",x"29170a",x"2a180b",x"301c0c",x"221409",x"1d1108",x"170f07",x"170f07",x"181007",x"1b1108",x"1b1108",x"1b1108",x"1e1408",x"1c1107",x"1f1309",x"25160a",x"231509",x"221509",x"251609",x"422511",x"412411",x"3d2310",x"1a1107",x"160f07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"1d1108",x"1d1108",x"1e1208",x"2c1b0b",x"2d1b0b",x"2d1b0a",x"1d1108",x"150e07",x"150e07",x"150e07",x"191007",x"170f07",x"191007",x"160f07",x"150e07",x"150e07",x"1d1108",x"160e07",x"160e07",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"26160a",x"3b2211",x"211309",x"221409",x"221409",x"211409",x"211409",x"28170a",x"371d0b",x"1a120a",x"1b110b",x"26170c",x"351e0f",x"412613",x"422713",x"392210",x"422812",x"4d2e15",x"462b14",x"442913",x"462913",x"3f2510",x"1f1309",x"311c0c",x"3d3229",x"3d3229",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"2d190b",x"28160a",x"311b0c",x"2d190b",x"2b170a",x"2d190a",x"2b180a",x"2b180a",x"28160a",x"261509",x"2b170a",x"2a1609",x"2a1609",x"2c180a",x"2b180a",x"291609",x"271509",x"271509",x"261509",x"2c180b",x"2a180a",x"281509",x"251408",x"2d180a",x"2e190b",x"321c0c",x"301a0b",x"341d0d",x"2d190b",x"301b0b",x"341d0d",x"311b0c",x"351e0d",x"351d0d",x"2f1b0c",x"341d0d",x"321c0d",x"2d1a0b",x"2e1a0b",x"291709",x"2e1a0b",x"281609",x"2f1a0b",x"311c0c",x"2f1b0c",x"2b180b",x"271509",x"2a180a",x"2e1a0b",x"27160a",x"261509",x"2d190b",x"2c180b",x"2f1a0b",x"301a0b",x"321c0c",x"2d190b",x"2b180a",x"2b180b",x"2c190b",x"2e1a0b",x"321c0c",x"351e0d",x"361e0d",x"351d0d",x"301b0c",x"2f1a0b",x"2a170a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c4d41",x"5c4d41",x"462711",x"432511",x"452711",x"432510",x"462611",x"492812",x"422410",x"472711",x"452711",x"41230f",x"3d210e",x"432410",x"42240f",x"3f220f",x"3d210e",x"3d210e",x"381d0c",x"371d0b",x"3d200e",x"3c200d",x"3c200d",x"3e200d",x"3a1e0c",x"381d0b",x"3c210e",x"41230f",x"3b1f0d",x"361a0b",x"371d0c",x"3f210e",x"3f220f",x"432510",x"452611",x"472711",x"462711",x"452610",x"432511",x"482812",x"452711",x"432611",x"462712",x"462812",x"442511",x"3a1f0c",x"40230e",x"472610",x"472710",x"3d210d",x"3c210d",x"472812",x"41240f",x"40230f",x"432510",x"4a2913",x"412410",x"452510",x"4a2912",x"452611",x"452610",x"452610",x"442510",x"452610",x"43240f",x"43240f",x"432510",x"432410",x"462711",x"492912",x"492812",x"452611",x"472811",x"402310",x"442510",x"42240f",x"432410",x"3f220e",x"422511",x"442711",x"4a2911",x"472610",x"44250f",x"4a2911",x"4d2b14",x"4e2c14",x"4f2e16",x"492813",x"4e2d16",x"492812",x"462711",x"462611",x"3f230f",x"462711",x"4a2912",x"27160a",x"27160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a180b",x"2a180b",x"2c1a0b",x"29170a",x"29180a",x"221409",x"211408",x"241608",x"2f1b0b",x"311c0b",x"331d0b",x"341f0c",x"3b240d",x"39220d",x"341f0c",x"361f0c",x"36200c",x"321d0c",x"351d0c",x"39200e",x"351c0c",x"332014",x"342a21",x"3f270f",x"37230b",x"38240b",x"37230b",x"301e0a",x"2b1b09",x"261809",x"1f1408",x"160f07",x"1c1208",x"170f07",x"181007",x"221409",x"201309",x"301c0c",x"301b0c",x"2d190b",x"2f1a0b",x"361f0d",x"371f0d",x"351f0c",x"38200e",x"38200e",x"432811",x"402611",x"482b13",x"4e2e15",x"4f2d15",x"472812",x"412612",x"3e2410",x"221409",x"201309",x"27170a",x"241509",x"26170a",x"27170a",x"27170a",x"28180a",x"251609",x"2a190a",x"2d1b0b",x"301d0b",x"321d0b",x"341f0c",x"3a240d",x"3c240d",x"39220c",x"35200b",x"301d0b",x"2a190a",x"251609",x"221309",x"3d2413",x"2c190c",x"221409",x"2a190b",x"45260f",x"41220d",x"371e0c",x"371e0c",x"3c200c",x"3c210d",x"381e0c",x"311b0b",x"331c0b",x"2b170a",x"29160a",x"261509",x"271409",x"271509",x"221308",x"241509",x"221408",x"27170a",x"3b210e",x"28170a",x"1b1108",x"1b1208",x"1c1107",x"1f1309",x"39200e",x"412611",x"412510",x"432510",x"361f0d",x"160e07",x"1b1108",x"170f07",x"1c1208",x"181007",x"191007",x"160f07",x"150e07",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"312820",x"24160a",x"3d2310",x"3f2512",x"221409",x"1f1208",x"221409",x"150e07",x"150e07",x"150e07",x"1c1108",x"170f07",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"221309",x"3b2311",x"231409",x"211308",x"201308",x"201309",x"211409",x"201309",x"391f0c",x"1a110a",x"1b120a",x"18110a",x"181009",x"311c0d",x"3a210f",x"3d2311",x"402511",x"422712",x"422611",x"492a13",x"4a2c13",x"3e2510",x"1d1208",x"1e1208",x"1e1208",x"1e1208",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1d1208",x"311c0c",x"351e0e",x"38200e",x"2a180b",x"2f1a0b",x"311b0c",x"321c0c",x"2c180a",x"2f180b",x"2e190b",x"38200e",x"331d0d",x"3b2210",x"341e0e",x"3c2210",x"351e0e",x"361f0e",x"311b0c",x"361f0e",x"351d0d",x"321b0c",x"341d0d",x"371f0e",x"39200f",x"39200f",x"39200f",x"3e2310",x"3d2310",x"412612",x"402512",x"402511",x"3d2411",x"3e2411",x"3c2310",x"38200f",x"361e0d",x"331c0d",x"341d0d",x"371f0e",x"301a0b",x"361e0c",x"371e0d",x"341c0b",x"39200f",x"331c0c",x"341d0c",x"331d0d",x"2a170a",x"2f1a0c",x"301b0b",x"311b0b",x"2c180a",x"311b0c",x"311b0c",x"301a0b",x"341d0d",x"301a0b",x"311b0b",x"301b0b",x"321c0c",x"331d0c",x"2e190a",x"331c0c",x"361e0d",x"391f0e",x"39200e",x"391f0e",x"381f0e",x"341d0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"655243",x"655243",x"492812",x"3f2310",x"3b200e",x"442711",x"422511",x"452812",x"472812",x"3e220f",x"3e220f",x"3b200e",x"3f230f",x"3b200e",x"361c0c",x"371c0c",x"3e230f",x"422611",x"432712",x"452913",x"432612",x"412511",x"432712",x"3f2310",x"432612",x"3e230f",x"3b200e",x"402310",x"412511",x"402511",x"422611",x"412511",x"422611",x"442712",x"452813",x"442813",x"482a14",x"472913",x"482a14",x"452813",x"442712",x"3f2310",x"3a200e",x"3f2410",x"462813",x"361d0b",x"3e220e",x"3c210e",x"42240f",x"40230e",x"381f0e",x"351d0c",x"3f2411",x"3d220f",x"3c210f",x"3f230f",x"3a200d",x"3b200e",x"3c210e",x"3d220f",x"3a1f0d",x"3e210e",x"3d210e",x"391f0d",x"3a200e",x"3b200e",x"3d220e",x"391f0d",x"3a1f0d",x"3b200d",x"3b200e",x"3e220f",x"402410",x"3f230f",x"422510",x"3e230f",x"3d210e",x"3f2410",x"3f2310",x"3c210d",x"3b210e",x"381e0c",x"3b200c",x"361d0b",x"3c210e",x"321b0b",x"452712",x"402310",x"412511",x"402410",x"442712",x"452712",x"412611",x"402511",x"432711",x"1b1108",x"1b1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b1a0a",x"2b1a0a",x"29180a",x"2a180a",x"2a180b",x"2c1a0c",x"221408",x"29180a",x"2f1b0b",x"311c0b",x"341f0b",x"38220c",x"37210c",x"3c240e",x"331f0b",x"36200d",x"321e0b",x"321d0b",x"301b0b",x"341c0c",x"381f0d",x"301c0f",x"211710",x"1b1108",x"311f0a",x"2d1c0a",x"2e1d0a",x"33200a",x"301e0a",x"2c1c09",x"1f1408",x"170f07",x"191107",x"191007",x"1a1107",x"251609",x"241509",x"301c0c",x"301b0c",x"2d190b",x"2f1a0b",x"361f0d",x"211309",x"201308",x"221409",x"1e1208",x"1e1208",x"221509",x"201309",x"170f07",x"170f07",x"1f1209",x"412612",x"311b0c",x"1f1208",x"1f1209",x"28170a",x"28170a",x"241509",x"251509",x"29180a",x"26160a",x"2d1b0b",x"29180a",x"28180a",x"2d1a0b",x"301d0b",x"2f1c0b",x"331e0b",x"38220c",x"38220d",x"36210d",x"341f0c",x"2d1b0a",x"2b180a",x"29180a",x"2a180b",x"372112",x"28170a",x"2d1a0b",x"2f1c0b",x"341f0c",x"3a230d",x"543217",x"4c2c14",x"442711",x"482912",x"472a12",x"462811",x"3b220e",x"321c0c",x"321c0c",x"28170b",x"361f0e",x"462711",x"1c1208",x"211408",x"211409",x"452915",x"462b17",x"000000",x"2a190a",x"361f0d",x"321d0d",x"321d0c",x"351e0d",x"1c1208",x"180f07",x"191007",x"160e07",x"191007",x"1d1208",x"1a1107",x"1a1107",x"170f07",x"160f07",x"221409",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"3c342c",x"201309",x"1e1208",x"1f1208",x"2a180a",x"1f1208",x"24150a",x"201309",x"21150b",x"150e07",x"221409",x"221409",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"25150a",x"341e10",x"221409",x"1f1208",x"1f1208",x"1d1108",x"1f1208",x"211408",x"3f230f",x"3f230f",x"181109",x"1b110a",x"19110a",x"29190c",x"3d2311",x"422713",x"442913",x"442812",x"452912",x"462913",x"492b14",x"3f2510",x"331d0d",x"1d1208",x"1d1208",x"1d1208",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"2d190b",x"2f1a0c",x"381f0e",x"311c0c",x"2f1b0c",x"2a180b",x"28170a",x"301b0c",x"2a180b",x"2f1b0c",x"2d1a0b",x"311b0c",x"29170a",x"311b0b",x"351e0d",x"3a210f",x"311c0c",x"3e2411",x"39200e",x"432612",x"422612",x"3b210f",x"3c230f",x"3e2311",x"3f2411",x"402411",x"422611",x"3e220f",x"3f2410",x"3f2310",x"3d2310",x"422612",x"452914",x"442813",x"452914",x"3a2210",x"3d2411",x"321c0c",x"381f0d",x"2e1a0b",x"311b0b",x"311c0c",x"2e1a0b",x"311c0c",x"311c0d",x"331d0d",x"29170a",x"2a180b",x"29170a",x"321c0d",x"321c0d",x"311c0c",x"351d0d",x"3d220f",x"3c2310",x"3e2411",x"3d2411",x"3b2210",x"39210f",x"3d2310",x"3f2410",x"3f2410",x"3e230f",x"442611",x"402410",x"3b210e",x"341d0d",x"2d190b",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"604e40",x"604e40",x"4c2c15",x"4b2a13",x"482711",x"4d2c14",x"4a2a13",x"4a2913",x"472711",x"4b2a13",x"492a12",x"4f2d15",x"4c2b13",x"4a2a12",x"4d2b14",x"4e2c14",x"4a2913",x"492912",x"4c2b14",x"482812",x"472611",x"40230f",x"4f2d15",x"442611",x"492913",x"502e16",x"4f2c15",x"533118",x"4f2f16",x"4a2a13",x"4a2a14",x"502e16",x"4f2d15",x"4c2b14",x"4c2b14",x"502e16",x"4c2b14",x"502d15",x"523017",x"553219",x"533118",x"513017",x"512f17",x"523218",x"4e2d15",x"4a2913",x"45260f",x"4a2811",x"42240f",x"462711",x"482c15",x"452610",x"4f2d15",x"4a2912",x"452711",x"472812",x"482811",x"4f2d15",x"533016",x"452510",x"4f2e15",x"4d2b14",x"533016",x"543118",x"512f17",x"512e16",x"502e16",x"4e2c14",x"482913",x"4c2b13",x"4d2b14",x"4d2c15",x"4b2b14",x"4b2a13",x"4c2a13",x"4a2912",x"4a2912",x"4d2b13",x"472812",x"371d0b",x"41230e",x"4b2912",x"43250f",x"43250f",x"4b2911",x"3a1f0c",x"472710",x"4d3017",x"4d2c14",x"492812",x"4b2b14",x"543118",x"523017",x"4d2b14",x"4e2d14",x"331d0d",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1b0b",x"2d1b0b",x"3a230f",x"3b230f",x"35210e",x"321d0c",x"2f1b0b",x"291809",x"361f0c",x"331d0c",x"36200d",x"3c240e",x"3b240e",x"442911",x"43280f",x"43280f",x"42260e",x"40250f",x"3e240f",x"422711",x"361e0d",x"3b2211",x"221409",x"201309",x"2c1c0b",x"36220b",x"301e0a",x"35210b",x"2e1d0a",x"1f1408",x"271909",x"1c1208",x"231608",x"191007",x"221608",x"341e0c",x"311c0b",x"211409",x"211409",x"221409",x"201308",x"1f1208",x"221409",x"1f1208",x"201208",x"221409",x"1e1208",x"1d1108",x"211409",x"201309",x"1f1209",x"26170a",x"26160a",x"25160a",x"241509",x"241509",x"231409",x"26160a",x"25160a",x"241409",x"231509",x"241509",x"24150a",x"27180a",x"2a180a",x"2b190b",x"2d1a0a",x"2e1b0a",x"311d0b",x"35200c",x"341f0c",x"37210c",x"311d0b",x"301d0b",x"231508",x"1f1308",x"1f1308",x"1e1209",x"211409",x"1d1208",x"2e1b0b",x"341f0c",x"39220d",x"341e0c",x"39200c",x"523116",x"492a12",x"42250f",x"472913",x"422611",x"412612",x"3b2110",x"351d0d",x"321d0d",x"331d0c",x"241609",x"231509",x"1c1108",x"27170a",x"462c1a",x"361e0d",x"2d190b",x"361f0d",x"2f1c0b",x"191007",x"181007",x"1a1107",x"191007",x"160f07",x"180f07",x"1a1107",x"1a1107",x"191008",x"201309",x"211409",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"211409",x"1d1108",x"201309",x"21170e",x"34281e",x"2f2015",x"21150a",x"211409",x"211409",x"201309",x"211409",x"201309",x"21150b",x"22150c",x"20150b",x"20150b",x"1e1208",x"1d1108",x"1c1108",x"1c1108",x"231509",x"3c2311",x"1f1208",x"221409",x"231409",x"1e1208",x"221308",x"271709",x"3a1f0d",x"412310",x"17100a",x"181009",x"19110a",x"1c1309",x"3d2512",x"3e2411",x"402510",x"492b13",x"3f2511",x"462a13",x"4e3015",x"432812",x"422510",x"23150a",x"1e1209",x"1e1209",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"311c0d",x"211309",x"1f1308",x"29180a",x"150e07",x"150e07",x"150e07",x"2d190b",x"381f0e",x"2b180b",x"3b220f",x"2d1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2410",x"1f1209",x"150e07",x"150e07",x"221409",x"3c220f",x"341f0e",x"211409",x"3c210f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"422510",x"371f0d",x"331c0c",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"514339",x"514339",x"4b2912",x"482811",x"4d2b13",x"4c2b14",x"462913",x"512f16",x"4d2b14",x"492812",x"4d2b13",x"502e15",x"522f16",x"482711",x"4d2b13",x"4e2c14",x"482711",x"4f2d15",x"523017",x"503117",x"4a2e15",x"4f2f15",x"502e15",x"472812",x"4e2f16",x"573319",x"4e2c14",x"58351b",x"4e2d15",x"56351a",x"54351a",x"5a381d",x"5c381c",x"55341a",x"59351a",x"5c381d",x"59351b",x"563419",x"543319",x"563419",x"5a381c",x"5b381c",x"5a361b",x"502f16",x"533118",x"56341a",x"482812",x"4a2913",x"472711",x"4f2d15",x"543118",x"573319",x"533017",x"512d15",x"4f2c14",x"482812",x"4a2912",x"4d2b14",x"522f16",x"5a361a",x"563218",x"512e16",x"512e16",x"553116",x"4f2c15",x"4c2b14",x"512d15",x"512e15",x"522e16",x"4e2b14",x"4e2b14",x"4f2b14",x"4a2813",x"4d2b13",x"492712",x"452610",x"4c2a14",x"482812",x"4f2d15",x"4a2911",x"432510",x"4a2911",x"482810",x"3f220d",x"45250f",x"4b2a11",x"3f220e",x"42240f",x"4d2d16",x"502e15",x"4c2a13",x"4c2c15",x"4a2912",x"4f2c14",x"4a2912",x"251509",x"251509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1a0b",x"2a1a0b",x"2b1a0b",x"2a190b",x"2c190b",x"2f1c0c",x"2c190b",x"29170a",x"311d0c",x"2f1a0b",x"2c190b",x"29180b",x"38200f",x"28170a",x"3b230c",x"3f250d",x"40260e",x"3e240e",x"3d230f",x"3f2410",x"361e0d",x"301a0b",x"281609",x"28180a",x"28180a",x"37220c",x"2f1d0a",x"2d1c0a",x"251708",x"1e1308",x"221608",x"211508",x"1f1408",x"1f1408",x"1a1107",x"231608",x"221608",x"211409",x"211409",x"221409",x"201308",x"201308",x"211309",x"1f1208",x"1d1108",x"1f1208",x"201208",x"201308",x"1f1208",x"211409",x"493528",x"241509",x"26160a",x"25160a",x"241509",x"241509",x"231409",x"251509",x"25160a",x"241509",x"241509",x"231509",x"2b180b",x"1e1309",x"301b0c",x"341e0c",x"311c0b",x"211508",x"201408",x"271809",x"261709",x"271809",x"2d1b0b",x"291909",x"221509",x"211408",x"201309",x"1e1209",x"211409",x"1d1208",x"1d1208",x"1f1309",x"1f1309",x"221409",x"1d1108",x"1d1208",x"40250e",x"432611",x"4f2f15",x"412610",x"472b14",x"39210f",x"36200f",x"4c2f17",x"3d220f",x"2d1a0b",x"1b1108",x"1b1108",x"2f1b0c",x"2f1b0c",x"331d0c",x"261609",x"1f1408",x"231608",x"231608",x"1a1107",x"170f07",x"181007",x"170f07",x"1b1108",x"1b1108",x"211409",x"201309",x"211409",x"221509",x"23150a",x"211409",x"211309",x"211309",x"201309",x"38200f",x"3a210f",x"371f0e",x"211409",x"241911",x"2d241d",x"24170c",x"1a1008",x"201309",x"211309",x"211409",x"221409",x"201309",x"22150b",x"20140b",x"20140b",x"20140a",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"3a2311",x"221409",x"201308",x"211308",x"1d1108",x"201308",x"271709",x"432812",x"160e07",x"150e07",x"171009",x"1b1209",x"2a1a0c",x"36200e",x"37200f",x"422711",x"3c2210",x"422711",x"412711",x"4c2c15",x"341c0c",x"412613",x"231509",x"201309",x"24150a",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"341e0d",x"27170b",x"180f07",x"150e07",x"150e07",x"2d1a0c",x"221409",x"1a1008",x"2b190b",x"150e07",x"170f07",x"150e07",x"1d1108",x"28180b",x"27160a",x"2e1a0c",x"341e0e",x"37200f",x"351e0e",x"3f2512",x"331f0e",x"382311",x"34200f",x"32200f",x"29190b",x"36200f",x"3f2612",x"382110",x"37200f",x"321d0e",x"3c2310",x"36200f",x"37200f",x"37200f",x"331e0e",x"150e07",x"231409",x"37200f",x"150e07",x"150e07",x"2c1a0c",x"2c190b",x"29180b",x"1e1208",x"462913",x"26160a",x"150e07",x"150e07",x"23150a",x"27170a",x"28170b",x"2c190b",x"2b190b",x"311c0c",x"311b0c",x"311b0c",x"311b0c",x"321c0c",x"341e0d",x"321d0d",x"3a200f",x"2c1a0c",x"361f0e",x"2f1c0d",x"2c1a0c",x"4d2d16",x"381f0e",x"351e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c4536",x"5c4536",x"472912",x"402410",x"412511",x"432612",x"412511",x"422611",x"472913",x"442712",x"482a14",x"482a14",x"482914",x"3d220f",x"3a1f0e",x"432611",x"402410",x"3f240f",x"412511",x"412511",x"402510",x"412410",x"442711",x"462913",x"402511",x"412611",x"412612",x"3f2611",x"452b15",x"412813",x"392411",x"432914",x"452913",x"462c15",x"4a2c16",x"4e2f16",x"4c2d16",x"482a14",x"492b15",x"4a2c15",x"492b15",x"472a14",x"442813",x"3e220f",x"3a200e",x"462a14",x"482a15",x"472a15",x"452813",x"412410",x"412511",x"422612",x"4d2d16",x"482a14",x"442813",x"462914",x"442712",x"3d2411",x"402410",x"432712",x"3f2310",x"3d220f",x"3d210e",x"3f230f",x"3e230f",x"452712",x"452812",x"432711",x"412511",x"462813",x"472913",x"482a14",x"4a2b15",x"462914",x"442713",x"482a14",x"432712",x"452812",x"442711",x"452812",x"41240f",x"41230f",x"351d0b",x"3f220e",x"42240f",x"371e0c",x"371e0d",x"3a200d",x"452813",x"3f2410",x"3e230f",x"3f2410",x"432611",x"422511",x"3f240f",x"231509",x"231509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1a0b",x"2b1a0b",x"2a190b",x"2c190b",x"2f1c0c",x"2c190b",x"3b3027",x"43372d",x"32271e",x"28170a",x"341d0d",x"402511",x"2c1a0c",x"24150a",x"24150a",x"24150a",x"221409",x"24150a",x"231409",x"24150a",x"271509",x"2c1a0b",x"271709",x"28180a",x"34200b",x"281909",x"271809",x"221508",x"211509",x"271809",x"291a09",x"231608",x"251709",x"251709",x"251809",x"231608",x"201409",x"201309",x"201309",x"201309",x"1e1208",x"1f1208",x"1b1108",x"1d1208",x"1d1108",x"1a1008",x"1c1108",x"1c1108",x"1b1108",x"402410",x"241509",x"25150a",x"26150a",x"251609",x"261609",x"2b1a0b",x"27160a",x"28170a",x"27170a",x"27170a",x"271709",x"231409",x"2c1f15",x"341e0d",x"221508",x"231608",x"231608",x"271909",x"271909",x"2b1b09",x"251708",x"221508",x"221608",x"1d1308",x"1d1208",x"190f08",x"180f07",x"191008",x"1a1108",x"1b1107",x"1e1209",x"1e1209",x"422611",x"25160a",x"221409",x"24160a",x"24160a",x"28180b",x"3a210e",x"482b14",x"432914",x"492c14",x"452811",x"4e2c13",x"39220c",x"371f0e",x"251509",x"361e0d",x"331f0b",x"251708",x"1d1208",x"1f1408",x"211508",x"251709",x"221508",x"170f07",x"170f07",x"160f07",x"22150a",x"23150a",x"23150a",x"201309",x"221409",x"221409",x"23150a",x"331c0d",x"39220f",x"341e0e",x"38200f",x"3c2310",x"402511",x"3a200e",x"452611",x"432611",x"3f2614",x"180f07",x"1e1208",x"211409",x"221409",x"211409",x"221409",x"221409",x"23160b",x"23160c",x"23160b",x"21150b",x"1e1209",x"1f1309",x"1e1209",x"1c1108",x"1c1108",x"24150a",x"24150a",x"211308",x"1e1208",x"201308",x"211408",x"271709",x"4b2d15",x"160e07",x"150e07",x"150e07",x"1b1108",x"2f1c0b",x"361f0d",x"3b2110",x"3c220f",x"432812",x"432811",x"432811",x"442811",x"432811",x"412411",x"28170a",x"221409",x"221409",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"37200f",x"150e07",x"150e07",x"201309",x"2c1a0c",x"311c0d",x"311b0c",x"2e1a0b",x"221409",x"432511",x"150e07",x"1c1108",x"27160a",x"2f1b0c",x"29160a",x"311b0c",x"351d0d",x"2f1a0b",x"311b0c",x"371f0e",x"39210f",x"3a210f",x"351e0e",x"301a0b",x"311c0c",x"311b0b",x"331c0d",x"361f0e",x"351e0d",x"321c0c",x"2e190b",x"321b0c",x"301b0c",x"341e0d",x"241509",x"2b190b",x"180f07",x"150e07",x"150e07",x"231409",x"27170b",x"311d0d",x"2b1b0c",x"22150a",x"392311",x"432713",x"150e07",x"23150a",x"341e0e",x"341f0e",x"331d0d",x"2d1a0b",x"301c0c",x"37200f",x"361f0e",x"39200f",x"361f0e",x"371f0e",x"3a210f",x"38200e",x"3c2210",x"3d2411",x"3c2310",x"3e2410",x"3a220f",x"4d2d15",x"341d0d",x"321c0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5d4a3d",x"5d4a3d",x"4a2912",x"442611",x"452712",x"492a14",x"402410",x"462812",x"452712",x"462812",x"442712",x"442712",x"462813",x"3f2310",x"3c210e",x"391f0e",x"3f220f",x"3f230f",x"402510",x"3e2310",x"422510",x"3e220f",x"3c200e",x"412410",x"3d210e",x"3c200e",x"3f2410",x"422511",x"442712",x"432612",x"3d220f",x"3c200e",x"422511",x"3c200e",x"442812",x"452812",x"412410",x"3c200e",x"3b200e",x"3d210e",x"402410",x"422611",x"462813",x"452813",x"381f0d",x"32190b",x"391f0d",x"442712",x"422914",x"452a15",x"422813",x"442b15",x"462914",x"4c2d16",x"4e2e17",x"4a2b15",x"422913",x"452812",x"422611",x"442711",x"472813",x"462813",x"452812",x"462813",x"452813",x"482a14",x"462812",x"452712",x"442713",x"492b15",x"462813",x"492a14",x"462813",x"462813",x"4a2c15",x"472812",x"432611",x"492a13",x"482914",x"452712",x"3f2310",x"472912",x"462710",x"371e0b",x"3b200d",x"371e0c",x"3f230e",x"472a14",x"462812",x"452812",x"422510",x"41240f",x"40230f",x"452611",x"3d210e",x"211309",x"211309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291b10",x"332418",x"31261f",x"40362d",x"382210",x"3a2311",x"412913",x"2f1c0d",x"2b1a0b",x"27170a",x"24160a",x"22150a",x"25160a",x"25160a",x"24150a",x"231509",x"221409",x"23150a",x"28180a",x"2e1d0a",x"382e25",x"311c0d",x"24160a",x"29190b",x"2e1b0d",x"39210f",x"211409",x"201309",x"1e1208",x"201309",x"201409",x"211409",x"221409",x"231409",x"221409",x"231409",x"221409",x"24160a",x"23150a",x"1b1008",x"180f07",x"191008",x"191008",x"1d1208",x"361e0d",x"231409",x"221409",x"221409",x"261609",x"241509",x"281709",x"271709",x"2c1a0a",x"2d1b0a",x"29180a",x"29180a",x"231509",x"432510",x"2b190b",x"211508",x"271809",x"291a0a",x"291a0a",x"291a0a",x"2a1a0a",x"251609",x"241609",x"241709",x"1e1309",x"1c1208",x"1c1107",x"170f07",x"170f07",x"170f07",x"180f07",x"191007",x"1c1107",x"402311",x"2b180b",x"28170a",x"2b180b",x"2b180b",x"261509",x"26150a",x"251509",x"4d2c14",x"351f0c",x"38200d",x"3b230d",x"39220c",x"43280f",x"3e240d",x"351f0b",x"43270f",x"2a1909",x"321d0c",x"301c0b",x"2b180a",x"231608",x"1f1408",x"27170a",x"24160a",x"27190e",x"3a3027",x"211309",x"1f1208",x"2b190b",x"1e1208",x"2b190b",x"211409",x"22150a",x"201208",x"231409",x"3e2411",x"2c1c0f",x"342111",x"382212",x"351f11",x"341e0f",x"351e0f",x"321c0c",x"2c1a0b",x"221409",x"221409",x"211409",x"231509",x"23150a",x"23160b",x"23160b",x"22160b",x"21150b",x"21150b",x"1e1209",x"1d1108",x"1c1108",x"1c1108",x"3e2414",x"221409",x"201308",x"28170a",x"271609",x"180f08",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"1b1108",x"2a180a",x"321c0b",x"371f0d",x"37200c",x"3f250e",x"3d220e",x"3f250e",x"492a10",x"442711",x"412411",x"28170a",x"221409",x"221409",x"000000"),
(x"150e07",x"150e07",x"150e07",x"180f07",x"29180a",x"351d0d",x"150e07",x"150e07",x"1c1108",x"2b180b",x"2b180b",x"241409",x"2d190b",x"221309",x"150e07",x"150e07",x"201309",x"2c190b",x"371f0e",x"38200e",x"351d0d",x"361f0e",x"351e0e",x"3b220f",x"3a210f",x"371f0e",x"371f0e",x"38200e",x"361f0e",x"37200f",x"39200f",x"361f0e",x"341e0e",x"331d0d",x"321c0d",x"2f1b0c",x"38200f",x"301c0d",x"1e1208",x"341d0d",x"3d220f",x"150e07",x"150e07",x"1c1108",x"2f1c0d",x"2d1b0d",x"2e1b0d",x"2f1c0d",x"2b1a0c",x"311e0e",x"150e07",x"150e07",x"1b1108",x"2f1b0c",x"2f1b0c",x"2c190b",x"2f1a0b",x"2c190b",x"2e1a0b",x"361f0e",x"361e0d",x"3a210f",x"361f0e",x"361e0d",x"321b0b",x"301a0b",x"2f1a0b",x"331c0c",x"2e190b",x"2e190a",x"452510",x"39200e",x"351e0d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"321c0c",x"321c0c",x"38200d",x"39200e",x"3b2110",x"3a2110",x"3b2110",x"402411",x"3f2311",x"3d2210",x"412412",x"412511",x"3c2110",x"381f0f",x"371f0f",x"361e0f",x"351e0f",x"341e0f",x"321d0e",x"301c0d",x"311c0e",x"311c0e",x"311c0e",x"5c4638",x"4c2b14",x"482812",x"4b2b14",x"4b2a13",x"482812",x"492812",x"462711",x"462711",x"462711",x"462711",x"452711",x"432611",x"472812",x"4a2912",x"4a2a13",x"492913",x"482913",x"4a2a13",x"4b2a14",x"472812",x"482912",x"482913",x"482812",x"42240f",x"432510",x"472812",x"472811",x"422511",x"4a2a14",x"4d2c15",x"4b2b14",x"492a13",x"4e2d15",x"4e2d15",x"4e2d15",x"4b2a14",x"4a2913",x"4a2a14",x"4f2e16",x"4c2c15",x"4a2913",x"4e2d16",x"4f2e16",x"523118",x"513118",x"4f2f17",x"4e2f17",x"4d2e16",x"462812",x"452711",x"492913",x"4f2d16",x"513017",x"523117",x"523117",x"4c2c15",x"4c2c15",x"523017",x"502f16",x"4e2d15",x"4a2a13",x"492913",x"462711",x"4c2b14",x"4b2b14",x"4c2c15",x"4d2d15",x"4d2d16",x"4a2a14",x"4d2c14",x"4c2b14",x"492a13",x"4c2c14",x"4d2d15",x"4c2c14",x"4d2c14",x"4e2d15",x"4c2c14",x"462712",x"482912",x"4b2b14",x"4a2b14",x"4e2d15",x"4d2d15",x"492a14",x"4b2b14",x"4d2d15",x"432510",x"41240f",x"442510",x"482711",x"492811",x"4a2912",x"2b180b",x"361e0e",x"351d0d",x"361e0d",x"38200e",x"39200f",x"3a200e",x"3b210f",x"3e2310",x"3c210f",x"3a200e",x"3e2310",x"3b210f",x"3c2210",x"381f0e",x"371e0e",x"3a210f",x"351d0d",x"331d0c",x"321c0c",x"301b0c",x"2f1a0c",x"2d1a0b",x"2b190b",x"2c190b",x"2d190b",x"2e1a0c",x"2f1a0c",x"311c0c",x"351e0e",x"36200e",x"341e0d",x"321c0c",x"331d0d",x"311c0d",x"2e1a0c",x"2b190b",x"26160a",x"221409",x"211309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e130b",x"22180f",x"302115",x"3a2f26",x"452914",x"4b2e17",x"432b14",x"3c2411",x"3c2410",x"331e0d",x"2a180a",x"231409",x"221409",x"211309",x"201308",x"23150a",x"221409",x"24150a",x"24150a",x"32261d",x"3c2f26",x"271c13",x"2a170a",x"2e190b",x"301b0b",x"311a0b",x"211308",x"1e1208",x"221509",x"201309",x"24150a",x"201309",x"221409",x"231409",x"231509",x"231409",x"221409",x"24160a",x"211309",x"201208",x"1f1208",x"221409",x"261609",x"371f0e",x"211309",x"3d2311",x"301c0d",x"2f1c0c",x"2d1a0b",x"2f1a0b",x"2a180b",x"28180a",x"28170a",x"2b190a",x"2c1b0a",x"271709",x"201408",x"412813",x"2a180a",x"271709",x"251609",x"261709",x"2a1a0a",x"2b1b0a",x"2b1a0a",x"281809",x"2a1909",x"221509",x"261709",x"261709",x"1d1208",x"1b1008",x"1b1008",x"1a1008",x"190f08",x"190f08",x"1a1007",x"1c1108",x"1d1208",x"1f1308",x"1c1108",x"1c1108",x"180f07",x"28180a",x"221509",x"341e0c",x"251609",x"2a1a0a",x"311e0b",x"321f0b",x"321f0b",x"2d1c0b",x"301e0b",x"321e0b",x"321f0b",x"2c1b0a",x"3d2410",x"2b190b",x"3f230f",x"3f230f",x"3a200f",x"2e1c10",x"382f26",x"43372c",x"442712",x"39200e",x"28180b",x"271b11",x"30261e",x"23150a",x"211409",x"201409",x"38200e",x"4a2912",x"21160d",x"21160c",x"21160d",x"25170b",x"25170b",x"25170c",x"27160a",x"27170a",x"211409",x"211309",x"1f1208",x"1f1208",x"1e1208",x"20140b",x"1f130a",x"1f130b",x"20140b",x"20140b",x"1d1209",x"1e1209",x"1c1108",x"2f1a0c",x"492a16",x"492a16",x"1a1008",x"1b1108",x"1a1108",x"180f07",x"190f07",x"191007",x"181007",x"160e07",x"1f1208",x"221409",x"2e1b0b",x"2b190a",x"2e190a",x"371f0c",x"3b220e",x"3d230e",x"3a210e",x"48290f",x"492c12",x"492c12",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1a0f07",x"2c190b",x"2b180b",x"2e1b0c",x"150e07",x"150e07",x"221409",x"28170a",x"28170a",x"2b190b",x"28170a",x"462711",x"150e07",x"150e07",x"1f1208",x"2b190b",x"2c190b",x"351e0e",x"2e1a0b",x"321d0d",x"2a190b",x"2c1a0c",x"311c0d",x"2c190b",x"351e0d",x"2e1a0c",x"301b0c",x"311c0d",x"311d0d",x"3b2310",x"331d0d",x"29160a",x"2f1b0c",x"23150a",x"150e07",x"482a14",x"201409",x"29180b",x"492b15",x"150e07",x"150e07",x"1c1108",x"29180a",x"23150a",x"27180b",x"150e07",x"3c2310",x"28190b",x"150e07",x"150e07",x"231409",x"321d0d",x"2c190b",x"3d2311",x"361f0e",x"2a180b",x"2f1b0c",x"361f0e",x"341d0d",x"351e0d",x"331d0d",x"37200f",x"37200f",x"3b2310",x"3b2411",x"2d1a0c",x"341d0d",x"482812",x"351d0d",x"341d0d",x"150e07",x"150e07",x"150e07",x"000000",x"2f1a0b",x"301b0c",x"321c0c",x"38200d",x"39200e",x"3b2110",x"3a2110",x"3b2110",x"402411",x"3f2311",x"3d2210",x"412412",x"412511",x"3c2110",x"381f0f",x"371f0f",x"361e0f",x"351e0f",x"341e0f",x"321d0e",x"301c0d",x"311c0e",x"311c0e",x"311c0e",x"321d0e",x"331d0f",x"2d190b",x"341e0e",x"321d0d",x"331d0d",x"311c0c",x"331d0d",x"311c0c",x"2e1a0b",x"321c0c",x"311b0c",x"301b0c",x"301b0c",x"2d190b",x"2e1a0b",x"301b0c",x"2e1a0c",x"2f1b0c",x"301b0c",x"301b0c",x"331d0d",x"351f0e",x"351f0e",x"321c0c",x"341d0d",x"341d0d",x"331c0c",x"321c0c",x"341d0d",x"38210f",x"39210f",x"3d2311",x"3d2310",x"341c0c",x"3c2210",x"3c2310",x"39210f",x"38200f",x"3d2411",x"3e2411",x"3b210f",x"3a200e",x"3d2310",x"402713",x"3f2813",x"3f2813",x"3c2612",x"37200e",x"371f0e",x"371f0e",x"39200f",x"402511",x"3f2410",x"3e2511",x"3e2410",x"3c220f",x"3e230f",x"422612",x"432712",x"452812",x"492b14",x"482a14",x"442712",x"432712",x"412511",x"402511",x"3d2310",x"3c2310",x"392310",x"3b210f",x"3b210f",x"3a220f",x"39210f",x"38200f",x"37200f",x"361f0e",x"371f0e",x"381f0e",x"3a210f",x"3b210f",x"3a200e",x"3c230f",x"3c220f",x"3b220f",x"381f0e",x"351d0d",x"361e0d",x"341d0d",x"341d0c",x"351d0d",x"361f0d",x"361e0d",x"371f0e",x"371f0e",x"361e0e",x"351d0d",x"361e0d",x"38200e",x"39200f",x"3a200e",x"3b210f",x"3e2310",x"3c210f",x"3a200e",x"3e2310",x"3b210f",x"3c2210",x"381f0e",x"371e0e",x"3a210f",x"351d0d",x"331d0c",x"321c0c",x"301b0c",x"2f1a0c",x"2d1a0b",x"2b190b",x"2c190b",x"2d190b",x"2e1a0c",x"2f1a0c",x"311c0c",x"351e0e",x"36200e",x"341e0d",x"321c0c",x"331d0d",x"311c0d",x"2e1a0c",x"2b190b",x"26160a",x"211309",x"1e1208",x"1b1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"24150a",x"221409",x"1d1309",x"1f150d",x"413226",x"3c220e",x"37200d",x"3a200d",x"331e0c",x"341f0d",x"311c0b",x"301d0b",x"3e230f",x"351e0d",x"25160a",x"24150a",x"231409",x"23150a",x"23150a",x"231509",x"231509",x"38261a",x"382d24",x"3f2511",x"422712",x"412812",x"402511",x"311b0c",x"28180a",x"29180a",x"211409",x"1f1309",x"1f1209",x"1f1209",x"27170a",x"2a190b",x"1e1209",x"1e1208",x"1e1208",x"2c1a0c",x"201208",x"1f1208",x"221409",x"261609",x"1f1208",x"26170a",x"3f2411",x"432712",x"3e2411",x"3f2511",x"37200e",x"39210e",x"412812",x"3f2914",x"3e2711",x"36200d",x"412510",x"4f3017",x"4e3017",x"221508",x"211508",x"2f1d0a",x"34200b",x"2e1c0b",x"2b1a0a",x"2e1c0a",x"28190a",x"231509",x"271809",x"271809",x"201308",x"1d1208",x"1f1308",x"1c1108",x"1b1008",x"211309",x"211309",x"1c1109",x"27180b",x"1f1408",x"1d1208",x"1c1108",x"1a1108",x"1a1008",x"211508",x"211409",x"23150a",x"26170a",x"2d1b0a",x"2f1d0b",x"2f1c0b",x"36210b",x"38220c",x"3a230d",x"36210c",x"301d0a",x"301d0b",x"29190a",x"321f0e",x"271a0e",x"311c0d",x"4a2f1d",x"48362a",x"443a30",x"463c33",x"3e2310",x"392414",x"493b2e",x"524134",x"4c4137",x"2f251d",x"322820",x"322920",x"33251a",x"39200e",x"22160d",x"23170e",x"24180d",x"25170c",x"26180c",x"27170c",x"27160a",x"211309",x"221509",x"261609",x"2a190a",x"28190b",x"2b1a0b",x"27180c",x"26180c",x"23160b",x"20150b",x"20150b",x"23150a",x"1d1208",x"1e1208",x"3f2411",x"482b16",x"1c1108",x"1b1108",x"1a1008",x"1c1208",x"180f08",x"180f07",x"1b1107",x"160f07",x"1d1108",x"26160a",x"27160a",x"2e1a0b",x"301c0c",x"341e0d",x"351d0c",x"42270f",x"351f0d",x"3c230e",x"442710",x"3d230e",x"3d230e",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"170e07",x"211409",x"331d0e",x"150e07",x"231409",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"26160a",x"442611",x"231409",x"371f0e",x"190f08",x"150e07",x"2e1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"2b190b",x"150e07",x"150e07",x"150e07",x"27170a",x"311c0d",x"4a2c15",x"150e07",x"150e07",x"150e07",x"150e07",x"402914",x"150e07",x"25160a",x"452913",x"150e07",x"28180b",x"38200f",x"351f0e",x"37200f",x"39210f",x"38210f",x"321d0e",x"331e0e",x"3d2411",x"341e0d",x"311b0c",x"331d0d",x"341d0d",x"321c0c",x"341d0d",x"27170b",x"351f0e",x"4e2d15",x"311c0d",x"361f0e",x"472813",x"442612",x"442612",x"2c1a0a",x"2f1c0b",x"2f1a0b",x"39210e",x"3c230f",x"3c2310",x"3d2412",x"3f2412",x"422713",x"442814",x"472a16",x"472a15",x"452814",x"452915",x"412612",x"3d2311",x"3a2111",x"382110",x"362010",x"341e10",x"321e0f",x"321d0f",x"311d0f",x"311d0e",x"311c0e",x"301c0e",x"301c0e",x"2f1a0d",x"301b0c",x"321c0d",x"331e0e",x"341e0e",x"321d0d",x"2f1b0c",x"2d190b",x"2b170a",x"2a160a",x"2e190b",x"301b0c",x"2f1b0c",x"2b180b",x"2c180b",x"2d1a0c",x"2e1a0b",x"301b0c",x"331d0d",x"331d0d",x"341e0e",x"341d0e",x"351e0e",x"361e0e",x"361f0e",x"38210f",x"371f0e",x"351f0e",x"321c0c",x"331d0d",x"39200f",x"39200e",x"3b210f",x"3d2310",x"3c2310",x"361f0e",x"38210f",x"37200f",x"38210f",x"39210f",x"39200f",x"3a210f",x"3a2210",x"3c2411",x"351e0d",x"39210f",x"3c2512",x"3d2613",x"392512",x"3f2511",x"3e2511",x"412612",x"412612",x"422612",x"432713",x"422612",x"432712",x"472a14",x"482a15",x"472914",x"472a15",x"442713",x"3e2310",x"3b210f",x"38200e",x"371f0e",x"361e0e",x"39210f",x"3b2311",x"392110",x"361f0e",x"351f0e",x"341e0e",x"321d0d",x"321c0d",x"36200f",x"38210f",x"39210f",x"3a2210",x"3a210f",x"3c2310",x"3c2310",x"3c2310",x"3c2210",x"3b2210",x"3a2210",x"39210f",x"37200f",x"361f0e",x"361f0e",x"351f0e",x"341d0e",x"351e0e",x"351e0e",x"341e0e",x"351f0e",x"36200f",x"39210f",x"38200e",x"3d2411",x"3b220f",x"3c210f",x"371e0d",x"38200e",x"3c2310",x"3b220f",x"3b2210",x"3a2210",x"39200e",x"371f0e",x"301a0b",x"2c180a",x"2c180a",x"2d190b",x"2b190b",x"29170a",x"27160a",x"2a180b",x"2c190b",x"2d1a0b",x"301c0c",x"301c0c",x"311c0d",x"321d0d",x"311c0d",x"301b0c",x"2d1a0c",x"2c190b",x"28170a",x"24150a",x"1f1309",x"1b1108",x"170f07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25160a",x"25160a",x"23150a",x"3d2310",x"432611",x"412511",x"3b220f",x"221409",x"27180d",x"3c2e23",x"453529",x"2a190a",x"2a180a",x"2d1a0a",x"311c0b",x"27160a",x"241509",x"432713",x"2e1b0d",x"23150a",x"1f130b",x"2a1a0e",x"382d23",x"3d230f",x"492912",x"462811",x"432811",x"462913",x"442811",x"36200e",x"2b1a0b",x"221509",x"1f1209",x"1e1208",x"1f1309",x"22140a",x"1e1209",x"1e1208",x"201309",x"25160a",x"26160a",x"2d190b",x"000000",x"33261c",x"1f1208",x"201309",x"2b190b",x"422612",x"3f2511",x"402511",x"2c1a0b",x"251509",x"2b1a0a",x"301d0b",x"3a210e",x"3d2510",x"432914",x"402712",x"4f3017",x"231608",x"29190a",x"2f1d0a",x"2d1c0a",x"2c1b0b",x"2c1b0b",x"271809",x"281809",x"271809",x"201309",x"2d1a0c",x"201309",x"371f0e",x"221409",x"1f1208",x"211409",x"1f1208",x"201309",x"201309",x"341d0d",x"1b1107",x"1b1108",x"1b1108",x"1c1108",x"1d1208",x"201308",x"24160a",x"25170a",x"2b1a0a",x"2f1d0b",x"311e0b",x"331f0b",x"36210c",x"38220d",x"35200c",x"36210c",x"37210c",x"331f0b",x"321e0c",x"26180d",x"1f1208",x"3f2411",x"422816",x"41342a",x"483d33",x"4f443a",x"4c2b15",x"462f20",x"554538",x"554537",x"55483c",x"4a3f36",x"483d34",x"40372d",x"382f27",x"2c1c0f",x"26190e",x"23170e",x"25180d",x"28190d",x"2b1b0d",x"2d1b0e",x"2b1a0c",x"28180b",x"231509",x"28180a",x"29190a",x"2b1a0a",x"2d1c0b",x"29190c",x"2d1c0c",x"26190c",x"22160b",x"221409",x"23150a",x"24160a",x"201308",x"1c1108",x"1b1108",x"1c1108",x"1e1308",x"1a1008",x"1e1208",x"1a1008",x"191008",x"1d1208",x"1d1208",x"1d1208",x"26160a",x"2c1a0c",x"2d1b0c",x"2e1b0c",x"331e0d",x"321d0d",x"3b230f",x"3b220f",x"3b2410",x"432812",x"39200d",x"39200d",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"170f07",x"231409",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"482913",x"3e2411",x"442813",x"331d0d",x"2b180b",x"2a180b",x"2b190b",x"28170a",x"25160a",x"2a180b",x"150e07",x"150e07",x"26160a",x"402512",x"452813",x"513017",x"402512",x"38200f",x"3f2411",x"452611",x"412511",x"3a2110",x"492a15",x"442611",x"412511",x"452712",x"442712",x"462813",x"3d2310",x"3e2411",x"4a2c16",x"533118",x"4b2b15",x"3c2210",x"502f17",x"4e2e16",x"412511",x"4a2b15",x"4d2d16",x"4c2c15",x"432712",x"2a180b",x"26160a",x"27170a",x"29170b",x"251509",x"2d190b",x"2e1a0c",x"2d1a0c",x"341e0e",x"351e0e",x"512f17",x"39200e",x"341d0d",x"462712",x"462712",x"462712",x"2f1b0b",x"2c1a0a",x"321e0d",x"341e0d",x"341e0d",x"36200f",x"382110",x"3b2311",x"3d2412",x"3e2412",x"3e2412",x"3e2511",x"3c2311",x"3a2110",x"361e0f",x"321d0e",x"2e1b0d",x"2c1a0d",x"29190d",x"27180c",x"27180c",x"27180d",x"25170b",x"25170b",x"26170b",x"26170c",x"27180c",x"29190c",x"2b1a0d",x"2c1a0d",x"2c1a0d",x"2a180b",x"29170a",x"2c1a0c",x"2d1a0c",x"2e1b0c",x"2e1b0c",x"2d1a0b",x"2a170a",x"2a170b",x"2c190b",x"2b180b",x"28160a",x"29170a",x"2a170a",x"2c190b",x"311c0d",x"321d0e",x"321d0d",x"321c0d",x"311b0c",x"341e0d",x"341d0d",x"341e0e",x"351f0e",x"331d0d",x"361f0f",x"37200f",x"3a210f",x"3d2411",x"3a2110",x"392110",x"36200f",x"331e0e",x"2d190b",x"311c0c",x"321d0d",x"331d0e",x"331d0d",x"321d0d",x"321d0d",x"321d0d",x"341e0e",x"321c0d",x"351f0e",x"3b2311",x"3d2411",x"3d2411",x"3b210f",x"3d2310",x"402612",x"3c2210",x"3f2411",x"3f2411",x"412612",x"412611",x"3f2411",x"3f2411",x"3b220f",x"3b220f",x"321b0c",x"311b0c",x"321d0d",x"321c0d",x"331d0d",x"331d0d",x"331d0e",x"321d0d",x"311c0d",x"2e1b0c",x"2d1a0c",x"2e1b0c",x"2f1c0d",x"311d0e",x"311d0d",x"321d0d",x"321d0d",x"321c0d",x"331d0d",x"331e0e",x"331e0d",x"331d0d",x"311c0d",x"2f1b0c",x"2d1a0c",x"2b190b",x"29180b",x"29170a",x"28160a",x"27160a",x"26160a",x"26160a",x"26160a",x"27170a",x"29180b",x"2c190b",x"2d1a0b",x"2f1a0b",x"301b0c",x"321c0c",x"331d0d",x"331d0d",x"321d0d",x"311c0d",x"301b0c",x"331d0d",x"351e0d",x"351f0e",x"321d0d",x"2e1a0c",x"28160a",x"251509",x"26150a",x"26160a",x"241509",x"251509",x"251509",x"26160a",x"2a180b",x"2c1a0c",x"2c1a0c",x"2b190b",x"28170a",x"28170a",x"26160a",x"221409",x"1f1309",x"1a1008",x"170f07",x"150e07",x"2a190b",x"2a190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201309",x"201309",x"1f1209",x"24150a",x"311c0c",x"442712",x"442712",x"402511",x"311d0d",x"31251c",x"4c392c",x"4a382c",x"4a382c",x"2a180a",x"2d1a0a",x"311b0b",x"27160a",x"241509",x"211309",x"3d2411",x"201309",x"1c1108",x"1d1208",x"3f220f",x"42240f",x"361e0c",x"341c0b",x"38200c",x"311c0a",x"321d0b",x"281709",x"241509",x"311c0c",x"3a210f",x"2c1a0c",x"201409",x"201309",x"201309",x"201309",x"201309",x"211309",x"28170b",x"2d190b",x"261a11",x"2c2017",x"36271d",x"25160a",x"301c0c",x"331d0d",x"361f0d",x"3a200e",x"331e0c",x"2e1c0b",x"2d1b0b",x"321e0b",x"331e0c",x"2f1c0b",x"2e1c0c",x"301c0c",x"2f1c0c",x"301c0c",x"29190a",x"2f1d0a",x"201309",x"201309",x"221509",x"3f2310",x"23150a",x"432511",x"2a180b",x"25160a",x"201409",x"24150a",x"211309",x"201208",x"211309",x"221409",x"251509",x"2b180b",x"3b210f",x"1b1108",x"1c1108",x"1d1208",x"1e1209",x"1f1309",x"211309",x"251609",x"29180a",x"2c1a0b",x"2d1c0b",x"2d1b0b",x"321e0c",x"35200c",x"321d0b",x"37220d",x"38220c",x"36210d",x"301d0c",x"28180a",x"24160a",x"3e2410",x"201309",x"412613",x"403328",x"4a4036",x"594b3f",x"1d1108",x"4b3323",x"57473b",x"5d4e42",x"58493d",x"4c4138",x"40362d",x"3b3128",x"3c332a",x"26180d",x"21160d",x"22160d",x"2c1c0d",x"2a1b0c",x"2d1b0e",x"2e1b0c",x"2a190b",x"29180b",x"402511",x"422611",x"482a12",x"472911",x"482a12",x"462913",x"452913",x"3c2310",x"24150a",x"23150a",x"2d1a0c",x"3c2311",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"201409",x"1e1208",x"1a1008",x"1b1108",x"231609",x"231509",x"201309",x"2a190b",x"2e1b0b",x"2a180b",x"301b0c",x"2d190b",x"351e0c",x"351f0c",x"361f0d",x"37200d",x"452812",x"3f250f",x"3f250f",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"190f08",x"231409",x"150e07",x"4a2a14",x"321c0d",x"341e0e",x"422612",x"482913",x"3f230f",x"482812",x"4d2c14",x"27170a",x"2b190b",x"3a200e",x"1a1008",x"150e07",x"150e07",x"1a1008",x"1e1208",x"1e1108",x"27170a",x"2b190b",x"27170b",x"221409",x"150e07",x"1a1008",x"492913",x"150e07",x"38200e",x"2d190b",x"341d0d",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"3d2310",x"301c0c",x"150e07",x"150e07",x"1b1108",x"1e1208",x"2c1a0c",x"2e1b0d",x"3c2311",x"502e17",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"28180b",x"361f0e",x"29170b",x"150e07",x"150e07",x"150e07",x"1b1108",x"27160a",x"2a180b",x"24150a",x"2e1a0b",x"2d190b",x"26160a",x"29180b",x"2e1a0c",x"2b190b",x"4b2b14",x"38200e",x"351e0e",x"422510",x"432510",x"3e2511",x"331d0c",x"2e1c0b",x"2d1a0b",x"2e1b0c",x"301c0f",x"311d0f",x"311d0e",x"341e0f",x"372010",x"361f10",x"341e0f",x"351e0f",x"321c0e",x"2f1c0f",x"2c1a0e",x"2a190e",x"27180d",x"24170e",x"22160d",x"1f150c",x"1f150c",x"20150c",x"20160c",x"21160d",x"22170e",x"22150c",x"23150b",x"24160c",x"26180c",x"27170c",x"29180d",x"28190c",x"28180c",x"27180c",x"2a1a0d",x"2b1b0d",x"29180b",x"2a180b",x"29170a",x"2e1a0c",x"2d1a0b",x"2e1b0c",x"2b180b",x"27160a",x"27160a",x"27160a",x"28170a",x"28170a",x"27160a",x"2c190b",x"2e1a0c",x"321d0d",x"331e0e",x"321d0e",x"2f1b0c",x"301b0c",x"321c0c",x"351e0e",x"331c0c",x"321c0c",x"351f0e",x"321d0d",x"301c0d",x"2d1a0b",x"241409",x"2b190b",x"2e1a0c",x"2f1b0c",x"301c0d",x"311d0e",x"301c0d",x"311c0d",x"331e0e",x"341e0e",x"351e0e",x"341e0e",x"341e0d",x"361f0f",x"371f0e",x"3a2210",x"39210f",x"39210f",x"361e0d",x"3b220f",x"39200f",x"3d2310",x"3d2310",x"371f0e",x"38200e",x"351e0e",x"331d0d",x"2f1b0c",x"2d1a0b",x"2c190b",x"2e1a0c",x"2e1a0c",x"2f1b0c",x"2f1b0c",x"2f1c0d",x"2f1b0c",x"2d1a0c",x"2c190b",x"2a180b",x"2a180b",x"2b190b",x"2c1a0c",x"2c190b",x"2c190b",x"2b190b",x"2b190b",x"2c190b",x"2b190b",x"27170a",x"25150a",x"231509",x"211309",x"1f1208",x"1f1208",x"1e1208",x"1c1108",x"1c1108",x"1b1108",x"1c1108",x"1d1108",x"201309",x"231409",x"26160a",x"29180b",x"28170b",x"29170a",x"2c190b",x"2c1a0c",x"2d1a0c",x"2e1b0c",x"2e1b0c",x"2e1a0c",x"301b0c",x"321e0e",x"2d1a0b",x"2a180b",x"241509",x"231509",x"231409",x"231509",x"23150a",x"201308",x"211309",x"211309",x"221409",x"221409",x"211309",x"221309",x"241509",x"231509",x"221409",x"1f1309",x"1a1008",x"170f07",x"150e07",x"150e07",x"301b0c",x"341d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201309",x"1f1309",x"201309",x"201309",x"392110",x"392110",x"231509",x"231509",x"472d1b",x"453528",x"42372e",x"453a30",x"463b31",x"463b31",x"000000",x"000000",x"000000",x"000000",x"000000",x"211309",x"221409",x"221409",x"211409",x"2c180a",x"3a200d",x"41240f",x"3a200d",x"341c0b",x"38200c",x"432612",x"432612",x"2e1a0c",x"211409",x"211308",x"241509",x"2e1a0b",x"351e0d",x"351e0d",x"321c0c",x"341e0e",x"351f0e",x"28170b",x"201309",x"2d190b",x"1f140a",x"1f140a",x"352316",x"2d190b",x"341d0d",x"371f0d",x"321c0c",x"3a200d",x"3a210d",x"351f0c",x"38220d",x"331e0b",x"331f0c",x"2f1c0b",x"2b190b",x"2a190b",x"2f1c0c",x"301c0c",x"241509",x"271709",x"1f1309",x"1f1309",x"2d190b",x"211409",x"2f1b0b",x"221409",x"211409",x"211409",x"211409",x"211409",x"221409",x"211409",x"231509",x"25160a",x"26160a",x"351f0c",x"35200d",x"3a210e",x"402610",x"3c230f",x"3b220f",x"402510",x"452811",x"231509",x"28170a",x"2c1b0b",x"2a1a0a",x"2d1b0b",x"2d1b0b",x"311d0b",x"301d0b",x"321d0b",x"35200c",x"331e0c",x"2d1b0a",x"2b1a0a",x"27180a",x"381f0d",x"381f0d",x"392110",x"3c3026",x"473b32",x"55453a",x"412512",x"4c3220",x"514032",x"5d4d41",x"5e5044",x"5e5044",x"3f362d",x"372d25",x"31281f",x"2f1c0d",x"28190e",x"291a0e",x"321f0e",x"35200f",x"38220f",x"36200e",x"361f0c",x"2d1b0b",x"321d0c",x"422611",x"482a12",x"472911",x"28170a",x"251609",x"2b1a0b",x"24150a",x"24150a",x"2b190b",x"3c2310",x"4c2c15",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"221509",x"1e1308",x"1c1108",x"1d1108",x"221509",x"221509",x"201309",x"241509",x"301c0b",x"241509",x"331e0b",x"2f1a0b",x"2b180a",x"341e0c",x"39210e",x"361f0d",x"452811",x"3b220f",x"3b220f",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"2e1b0c",x"150e07",x"412510",x"311c0d",x"452712",x"150e07",x"3a210f",x"361e0d",x"371e0d",x"150e07",x"412511",x"150e07",x"150e07",x"1f1208",x"201308",x"29170a",x"2c190b",x"301c0c",x"2f1b0c",x"29180a",x"28160a",x"1b1008",x"1f1208",x"452611",x"150e07",x"150e07",x"311c0d",x"351e0d",x"402410",x"150e07",x"1f1309",x"2a180b",x"2e1a0c",x"29170a",x"2d190b",x"28170a",x"361f0e",x"452814",x"231509",x"201308",x"321c0c",x"3c220f",x"482a13",x"150e07",x"150e07",x"1b1108",x"29180b",x"361f0f",x"37200f",x"301c0d",x"29180b",x"462913",x"4c2b14",x"150e07",x"28170b",x"2f1b0c",x"29180b",x"341d0d",x"37200f",x"331d0d",x"331c0c",x"331c0c",x"341d0c",x"321c0c",x"331c0c",x"311b0c",x"482812",x"3b220f",x"331c0c",x"412410",x"422410",x"4e2f15",x"3d2310",x"321d0b",x"2f1b0b",x"321d0f",x"372010",x"341e0f",x"361f0f",x"3b2212",x"3b2311",x"3b2312",x"382010",x"362112",x"342012",x"2d1c10",x"291a0f",x"27190f",x"24180f",x"241a11",x"211710",x"221810",x"211811",x"221810",x"221810",x"21170f",x"22170f",x"24180f",x"25180f",x"24180f",x"25170d",x"26190e",x"26190e",x"26180e",x"26180d",x"25170b",x"27180c",x"28180c",x"29180c",x"27160a",x"27160a",x"271609",x"2d190b",x"2b190b",x"29170a",x"27160a",x"251509",x"27160a",x"28170a",x"2a180b",x"2b190b",x"2b190b",x"2c190b",x"2a170a",x"2b180a",x"2c190b",x"2f1b0c",x"311c0c",x"341d0d",x"351e0d",x"331d0d",x"321c0c",x"311c0c",x"301b0c",x"2d190b",x"28160a",x"2a170a",x"29170a",x"2e1b0c",x"2f1c0d",x"2f1b0c",x"29170a",x"29170a",x"2d1a0b",x"311c0d",x"321c0d",x"331d0d",x"361f0e",x"361f0e",x"38210f",x"392210",x"38200f",x"38200f",x"37200f",x"38200f",x"361f0e",x"38200f",x"3b2310",x"381f0e",x"371f0e",x"361f0e",x"351f0e",x"2f1b0b",x"2a180a",x"29170a",x"2a170a",x"28160a",x"29170a",x"2c190b",x"2f1b0c",x"2e1b0c",x"2f1b0c",x"331d0d",x"311c0d",x"2a170a",x"261509",x"261609",x"29180b",x"29180b",x"29180b",x"29180b",x"29180b",x"2a180b",x"2a180b",x"26160a",x"25150a",x"231509",x"201309",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"191008",x"190f08",x"180f07",x"191008",x"1b1008",x"1d1108",x"1f1208",x"211309",x"241509",x"231409",x"251509",x"26160a",x"28170a",x"28170a",x"28170a",x"2a180b",x"301c0c",x"2e1b0c",x"2d1a0b",x"29170a",x"231409",x"1f1208",x"1f1208",x"211309",x"201309",x"201309",x"201309",x"1f1208",x"201309",x"231409",x"221409",x"221409",x"211409",x"1f1208",x"1e1208",x"1c1108",x"1a1008",x"170f07",x"160e07",x"1b1008",x"341d0e",x"3b210f",x"462712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1208",x"1e1208",x"201309",x"201309",x"1d1108",x"2e1b0c",x"2e1b0c",x"2a180b",x"3f2410",x"412613",x"443429",x"473c32",x"4a3f35",x"4b4036",x"4b4036",x"000000",x"000000",x"000000",x"26170a",x"261709",x"241609",x"221409",x"211409",x"211409",x"201309",x"1f1309",x"1f1309",x"1e1208",x"3a3129",x"000000",x"3a210f",x"361f0e",x"211409",x"1f1208",x"211309",x"221409",x"2e1a0b",x"351e0d",x"361e0d",x"2f1b0c",x"2b180b",x"211409",x"3b2210",x"221509",x"2d190b",x"1d1208",x"1d1208",x"2f1c0f",x"341e0d",x"3b220f",x"3a210e",x"40240f",x"442710",x"361f0c",x"38200c",x"3e240e",x"3a230d",x"37200c",x"341f0c",x"301c0a",x"2a180a",x"241609",x"2a190a",x"241509",x"2a190a",x"2a180a",x"251509",x"231409",x"24160a",x"231509",x"221409",x"211409",x"211409",x"211409",x"311c0d",x"28170a",x"29180b",x"2a180b",x"2e1b0b",x"38200d",x"351f0c",x"271809",x"201408",x"251708",x"231509",x"221509",x"2b180a",x"472913",x"432510",x"1f1309",x"211408",x"231509",x"27170a",x"28180a",x"331e0c",x"2d1b0b",x"34200c",x"2f1c0b",x"35200c",x"331f0c",x"341f0c",x"2e1c0b",x"29190b",x"361f0e",x"331e0e",x"402d20",x"46372b",x"432711",x"4b2b15",x"492f1e",x"524033",x"54463a",x"54493e",x"1e1209",x"1f1309",x"1f1309",x"21160d",x"3b2210",x"25180d",x"2c1c0d",x"301d0e",x"3e2510",x"3f2610",x"3b230d",x"36200d",x"331e0c",x"351f0d",x"351f0d",x"000000",x"26160a",x"26160a",x"2c1a0b",x"301d0d",x"2a180b",x"201409",x"201309",x"1c1108",x"211409",x"2d1a0c",x"29170b",x"2b170a",x"2a170a",x"331d0d",x"351f0e",x"321d0d",x"37200d",x"371f0e",x"37200e",x"3d230f",x"361f0e",x"371f0e",x"39200f",x"351e0d",x"3d230d",x"2e190b",x"2e1a0b",x"351e0c",x"37200d",x"331d0c",x"3f240f",x"371d0c",x"371d0c",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1d1208",x"2a190b",x"180f08",x"412410",x"311c0d",x"301c0d",x"3a2110",x"462913",x"150e07",x"3b210f",x"482812",x"150e07",x"1f1209",x"2b190b",x"321c0c",x"2f1b0c",x"311c0c",x"2e1a0b",x"331d0d",x"2d1a0b",x"241509",x"150e07",x"391f0e",x"211309",x"150e07",x"150e07",x"3b200e",x"150e07",x"150e07",x"150e07",x"211409",x"2e1a0b",x"2a170a",x"351e0d",x"301b0c",x"341d0d",x"351f0e",x"25160a",x"402411",x"2f1b0c",x"231509",x"331d0d",x"482812",x"3d2310",x"150e07",x"150e07",x"28160a",x"29170a",x"2e190b",x"2f1a0b",x"351d0d",x"2f1a0b",x"28160a",x"150e07",x"150e07",x"27160a",x"2e1a0c",x"2a180b",x"361e0e",x"351e0d",x"331e0e",x"3a210f",x"2f1b0c",x"331d0d",x"39200e",x"361f0e",x"311c0d",x"4d2d15",x"3a210f",x"321c0c",x"442610",x"432610",x"4a2b14",x"432711",x"3a220e",x"3c2311",x"3f2512",x"3a2110",x"3a2110",x"381f0f",x"371f0f",x"361f0f",x"382010",x"372011",x"362011",x"362011",x"331e11",x"2e1d10",x"321f12",x"301e12",x"2e1e12",x"2a1b11",x"2b1b11",x"2a1b10",x"2a1b11",x"291b11",x"2d1c12",x"322013",x"311e10",x"2f1d11",x"301e11",x"342012",x"362011",x"382212",x"382212",x"341f10",x"361f0f",x"362010",x"382111",x"372011",x"38200f",x"331c0d",x"351d0d",x"361f0e",x"331d0d",x"361f0e",x"341d0d",x"331c0d",x"351d0d",x"361f0e",x"351e0d",x"361f0e",x"371e0d",x"361e0d",x"361e0d",x"351e0d",x"371f0e",x"3b220f",x"341c0d",x"381f0d",x"391f0d",x"381f0e",x"381f0e",x"39200e",x"361d0d",x"331c0d",x"341d0d",x"371f0e",x"38200f",x"3b220f",x"3b220f",x"371f0e",x"371f0e",x"361f0e",x"361e0d",x"39210f",x"3c2310",x"381f0e",x"361e0d",x"361e0d",x"381f0d",x"341d0c",x"3a200e",x"351e0d",x"361e0d",x"3a200e",x"3e2310",x"3c210e",x"3c210f",x"3e2310",x"3e2310",x"3e2310",x"402511",x"3b220f",x"37200e",x"321d0d",x"361f0e",x"351e0e",x"361f0e",x"38200f",x"321d0d",x"38200f",x"39210f",x"38200e",x"39200e",x"39210e",x"3c220f",x"39200e",x"39210f",x"39200f",x"321c0d",x"2e1a0b",x"2e190b",x"29160a",x"2d190a",x"2c180a",x"2a170a",x"2e1a0b",x"2a170a",x"271609",x"221309",x"251509",x"27160a",x"221309",x"241409",x"211308",x"261509",x"241409",x"251409",x"27160a",x"29170a",x"2d190b",x"2d1a0b",x"311c0c",x"341e0d",x"311c0d",x"341e0e",x"331d0d",x"321c0c",x"37200f",x"341e0e",x"361f0f",x"341e0e",x"2e1a0c",x"2a180b",x"2b180b",x"311c0c",x"2e1a0c",x"2d1a0b",x"2b190b",x"2b190b",x"2e1b0c",x"2d1a0b",x"2e1a0c",x"2c190b",x"2d190b",x"2c180b",x"2c190b",x"2c190b",x"2d1a0c",x"2a180b",x"251509",x"26160a",x"2c190b",x"462712",x"462712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201409",x"201409",x"201309",x"201309",x"201309",x"28180b",x"221409",x"2f1c0d",x"1b1108",x"371f0f",x"3b2e23",x"483c33",x"59493e",x"56473c",x"56473c",x"221509",x"28180a",x"251509",x"26170a",x"251609",x"251609",x"231509",x"221409",x"211409",x"211409",x"221509",x"221509",x"3a3129",x"3a322a",x"30261d",x"4a2b15",x"4a2b15",x"211409",x"221409",x"221409",x"211409",x"211409",x"000000",x"452912",x"3a220e",x"28190a",x"2c1a0a",x"291c11",x"352b22",x"342a22",x"201409",x"1e1308",x"20140b",x"3c210f",x"1f1208",x"201309",x"1d120b",x"2e251e",x"331d0d",x"361f0e",x"3f260f",x"3d250e",x"3c240e",x"3a220e",x"321d0b",x"311c0b",x"2f1b0b",x"28170a",x"2a190b",x"25160a",x"28180b",x"28180b",x"26170a",x"231509",x"231509",x"27170a",x"2a1a0a",x"26170a",x"1f1309",x"201309",x"1d1208",x"1c1108",x"1c1108",x"201409",x"261809",x"241609",x"221509",x"251709",x"271809",x"251709",x"231609",x"1c1108",x"3c210e",x"1f1208",x"27160a",x"211408",x"27170a",x"27170a",x"28180a",x"331e0c",x"2f1c0b",x"34200c",x"35200c",x"3d230d",x"3a220d",x"412710",x"402510",x"2d1c0b",x"29190a",x"28170a",x"2d1a0c",x"331d0c",x"301c0b",x"452711",x"432812",x"2c2016",x"21170f",x"3f362d",x"27160a",x"1f1208",x"1f1208",x"1e1208",x"211409",x"341e0e",x"412411",x"492b14",x"492a13",x"4a2a12",x"472a12",x"482a12",x"432611",x"452812",x"452812",x"231509",x"000000",x"26160a",x"2c1a0b",x"211409",x"201409",x"201309",x"27170a",x"38200e",x"38200e",x"221409",x"231409",x"231509",x"231509",x"25160a",x"25150a",x"221409",x"201309",x"1f1208",x"1d1208",x"1c1208",x"1c1108",x"1d1208",x"1f1308",x"1f1209",x"20130a",x"170f07",x"1c120a",x"201309",x"211409",x"1d120a",x"231911",x"41240f",x"41240f",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"311c0c",x"1d1208",x"492a14",x"321d0d",x"3b2210",x"4c2c15",x"150e07",x"3e2411",x"29180b",x"2b190b",x"150e07",x"2d1a0c",x"37200f",x"361f0e",x"331d0d",x"331d0d",x"301c0d",x"321d0d",x"201309",x"2b190c",x"492a13",x"150e07",x"150e07",x"1c1108",x"482a14",x"150e07",x"150e07",x"2b190b",x"2e1b0c",x"331d0d",x"3a2110",x"3c2310",x"3b2310",x"3d2411",x"3a200f",x"3b2210",x"2d1a0c",x"3d2411",x"512f17",x"301c0d",x"512f18",x"150e07",x"150e07",x"513017",x"150e07",x"150e07",x"29180b",x"2d1a0c",x"2d1a0c",x"331d0e",x"29180b",x"402511",x"502d15",x"150e07",x"1f1208",x"2d1a0b",x"2f1c0d",x"321e0e",x"301c0d",x"2e1b0c",x"361f0e",x"351f0d",x"2b190b",x"39200f",x"321c0d",x"2e1b0c",x"4d2c14",x"38200e",x"341d0d",x"422410",x"422410",x"523117",x"482811",x"432611",x"3f2311",x"412510",x"402310",x"402311",x"412512",x"3e2211",x"452713",x"452815",x"442715",x"3f2513",x"382011",x"3a2112",x"422715",x"412716",x"452a16",x"402616",x"3a2314",x"402615",x"3f2616",x"422716",x"452a17",x"452917",x"432817",x"422714",x"462a17",x"452816",x"442916",x"442815",x"452915",x"422714",x"422714",x"432713",x"432713",x"452913",x"432713",x"492c15",x"462812",x"462813",x"432511",x"442712",x"442712",x"412511",x"412511",x"432712",x"432611",x"472913",x"482a14",x"4a2b15",x"422410",x"482914",x"472712",x"462914",x"492a14",x"4b2c15",x"462813",x"442714",x"472814",x"492a15",x"4a2b16",x"492b15",x"4b2d16",x"492d17",x"472a16",x"492c17",x"4b2d17",x"492c17",x"492c17",x"472b16",x"482b16",x"4a2d18",x"4c2d19",x"4c2f19",x"4d2f1a",x"4d2f19",x"4c2e19",x"452916",x"492b17",x"4a2d18",x"50311b",x"4b2d18",x"432814",x"482a15",x"482a16",x"432613",x"4f3019",x"523219",x"4c2e18",x"4a2c16",x"482b16",x"432715",x"422814",x"432814",x"432814",x"412714",x"452915",x"402613",x"402512",x"442814",x"422613",x"3f2413",x"3c2312",x"402412",x"3e2412",x"3f2312",x"3e2210",x"391e0e",x"3b200f",x"351c0d",x"381f0f",x"3b2110",x"3b2110",x"371e0f",x"331b0d",x"331c0d",x"371e0e",x"3a2010",x"392110",x"3b2110",x"371f0f",x"381f0f",x"391f0f",x"3a2110",x"3b2211",x"3d2411",x"3d2311",x"3b2110",x"3c2211",x"3f2412",x"3e2312",x"442712",x"422612",x"412511",x"402511",x"422611",x"412410",x"452812",x"432712",x"412511",x"3d2310",x"412612",x"39200e",x"3f2411",x"432612",x"3f2411",x"3d230f",x"412511",x"412511",x"402511",x"3b2110",x"3e2310",x"3e2310",x"402511",x"3f2210",x"442712",x"432713",x"432713",x"412511",x"3e2410",x"3f2310",x"452611",x"452611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221408",x"221509",x"24160a",x"221509",x"221409",x"22150a",x"402511",x"472813",x"472813",x"402612",x"423125",x"493c31",x"5a483a",x"59493e",x"221409",x"221509",x"241509",x"29190a",x"28180b",x"27180a",x"27170a",x"29190b",x"28170b",x"251609",x"251609",x"221509",x"211309",x"332a23",x"32241b",x"271a0f",x"3b210f",x"25160a",x"26160a",x"201309",x"201309",x"201309",x"221409",x"221409",x"452912",x"452912",x"402411",x"3a271a",x"3b2f25",x"3a3027",x"26170a",x"251609",x"201308",x"341e0c",x"361e0e",x"2f190b",x"291e16",x"2a211a",x"332a22",x"361f0e",x"1f1209",x"1d1108",x"1d1108",x"1e1208",x"3a220e",x"361f0d",x"321c0c",x"351f0d",x"3d230f",x"3a210e",x"39200e",x"3b230f",x"24150a",x"251609",x"26170a",x"28180a",x"27180a",x"27190a",x"1e1208",x"211409",x"211409",x"201309",x"201409",x"1f1309",x"201309",x"211409",x"221409",x"211409",x"211409",x"201309",x"201309",x"201309",x"211409",x"39200e",x"3f2d20",x"22140a",x"23160a",x"27170a",x"2c1b0b",x"29190b",x"321f0c",x"321f0b",x"2f1d0b",x"37220c",x"35200c",x"38220d",x"36210c",x"301d0b",x"2d1c0a",x"4d2e15",x"27170a",x"39200d",x"331d0c",x"301c0b",x"29180b",x"28170a",x"24150a",x"231509",x"482a15",x"311c0d",x"29180b",x"2d1a0c",x"2e1a0c",x"27170b",x"22150a",x"221409",x"1a120b",x"1d1108",x"231409",x"24160a",x"25160a",x"25160a",x"24160a",x"24150a",x"1f1208",x"231509",x"241509",x"231509",x"271c13",x"281d14",x"281e15",x"33241a",x"2e1c0d",x"201409",x"221409",x"211409",x"211309",x"211309",x"241509",x"261709",x"241609",x"211308",x"1f1108",x"1e1208",x"27160a",x"321c0c",x"371e0d",x"301a0b",x"3b3026",x"1e160f",x"1c130b",x"321c0d",x"381f0e",x"291d15",x"2c231c",x"352c23",x"3c332a",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"201309",x"2f1b0c",x"1f1208",x"3f2310",x"351e0e",x"2f1a0c",x"150e07",x"2a180b",x"1b1108",x"150e07",x"392110",x"150e07",x"311c0d",x"2e1a0c",x"2b190b",x"301b0c",x"311c0c",x"29180b",x"27160a",x"472912",x"26160a",x"150e07",x"1f1309",x"27170b",x"26160a",x"513016",x"150e07",x"1d1208",x"2b190b",x"2f1b0c",x"311d0d",x"351e0e",x"39210f",x"37200f",x"3c2311",x"3a210f",x"341d0d",x"231409",x"341c0c",x"311b0c",x"3b220f",x"150e07",x"150e07",x"221409",x"150e07",x"412612",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1a0c",x"492912",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"221409",x"1c1108",x"25150a",x"26160a",x"1d1108",x"170f07",x"1f1208",x"28170a",x"4c2b14",x"311b0c",x"341d0d",x"452711",x"452711",x"492a14",x"4a2b14",x"492a15",x"4a2b17",x"4b2c16",x"4f2e19",x"502e19",x"512f18",x"4e2d17",x"492a16",x"4b2c18",x"462816",x"492b17",x"432715",x"432817",x"412515",x"3c2315",x"382013",x"2f1b11",x"351d11",x"432815",x"482b17",x"482c17",x"462a17",x"492b17",x"452917",x"472916",x"462915",x"502f19",x"4e2f18",x"4d2d17",x"4d2c16",x"4a2a15",x"482914",x"492a15",x"462713",x"4a2b15",x"492a14",x"4e2d16",x"543117",x"533018",x"523017",x"4d2c15",x"4d2c14",x"4c2b14",x"482812",x"4a2a13",x"4e2d14",x"4d2d14",x"4d2c14",x"4c2b14",x"512e15",x"4d2c14",x"512f17",x"4f2f16",x"533218",x"513017",x"533119",x"512f18",x"502f18",x"513019",x"53321a",x"53321b",x"54321c",x"55341c",x"55351e",x"502f19",x"482b19",x"472b18",x"4a2d1a",x"4e301b",x"4e2e1b",x"51311c",x"53331d",x"54341e",x"55351d",x"54341d",x"55331d",x"52321c",x"54341d",x"4b2d19",x"52311c",x"51311c",x"51301c",x"51321c",x"54331c",x"51311c",x"52311b",x"53321b",x"482b17",x"4e2e19",x"51301b",x"4e2f1a",x"4b2c18",x"452816",x"422514",x"4b2c18",x"4f2f19",x"4f2f19",x"4d2d19",x"492a17",x"492b17",x"4b2b17",x"4c2c15",x"452815",x"4c2c16",x"4b2c16",x"4f2e17",x"4c2c16",x"4c2d16",x"4d2d17",x"472915",x"4a2b16",x"442612",x"412413",x"432612",x"3f2211",x"3f2211",x"3e2211",x"3b1f0f",x"29150a",x"2e170b",x"422512",x"472914",x"492a14",x"472914",x"452714",x"462814",x"432613",x"432511",x"4b2a14",x"4e2e17",x"4c2b15",x"4b2b14",x"4a2912",x"4a2912",x"4a2913",x"4c2b14",x"482812",x"4d2c14",x"4a2a13",x"4c2b15",x"502e16",x"502f16",x"482913",x"4f2e15",x"4c2c14",x"4c2b14",x"4a2913",x"4b2a14",x"4b2b14",x"432611",x"492a13",x"482812",x"4a2a14",x"4d2c15",x"4f2e16",x"4e2d15",x"502e16",x"502e16",x"512e16",x"543117",x"4e2d15",x"4e2d15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25160a",x"251609",x"211409",x"1f1208",x"201309",x"211409",x"201309",x"39200e",x"39200e",x"422611",x"341e0e",x"442d1f",x"46362b",x"1f1208",x"231509",x"221409",x"211409",x"28190a",x"28180a",x"2c1b0a",x"2a190a",x"2e1c0b",x"301d0b",x"2a1a0a",x"271709",x"25160a",x"231509",x"221408",x"30271f",x"29190d",x"170f07",x"3b220f",x"3b220f",x"211409",x"201309",x"201209",x"201208",x"221409",x"211409",x"2a180b",x"432410",x"442a18",x"453529",x"41362c",x"473b31",x"28180a",x"26170a",x"2a180b",x"27160a",x"2c190b",x"3a291d",x"483c32",x"4d3f34",x"453b33",x"462812",x"180e07",x"190f07",x"1e1108",x"201308",x"201308",x"361f0d",x"231509",x"231509",x"231509",x"1f1308",x"29170a",x"2c190b",x"361e0d",x"2c1a0b",x"36200d",x"2f1c0b",x"2c1a0a",x"1e1208",x"1f1309",x"341d0d",x"211409",x"201309",x"201309",x"201309",x"201309",x"201309",x"211409",x"201309",x"201309",x"211409",x"211409",x"201309",x"2a180b",x"191008",x"1a1109",x"24150a",x"251609",x"251609",x"27170b",x"28180b",x"2a1a0b",x"2c1b0b",x"2f1d0b",x"34200c",x"311e0c",x"34200c",x"34200c",x"321e0c",x"2e1c0b",x"38200e",x"302013",x"2a180a",x"231609",x"251709",x"2a1a0a",x"281909",x"251609",x"231509",x"211409",x"211409",x"221509",x"221309",x"201309",x"201309",x"201309",x"1f1208",x"2e251d",x"221409",x"211309",x"211409",x"23150a",x"211309",x"221409",x"231409",x"231409",x"231509",x"241509",x"24150a",x"221409",x"3f362c",x"3f362d",x"352b22",x"2f251c",x"381f0d",x"211309",x"211309",x"211408",x"251509",x"26170a",x"27170a",x"2b1a0a",x"26170a",x"27170a",x"261609",x"201308",x"201308",x"2a170a",x"321c0b",x"453b32",x"2f2720",x"241c15",x"27170a",x"2d2018",x"41362d",x"494037",x"41382f",x"41372e",x"41372e",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"2e1b0c",x"1d1208",x"4a2a14",x"3f240f",x"150e07",x"432510",x"27160a",x"150e07",x"2c190b",x"442612",x"150e07",x"1d1208",x"2f1b0c",x"26160a",x"24150a",x"150e07",x"351f0e",x"4e2d14",x"150e07",x"150e07",x"24150a",x"2a180b",x"2d1a0b",x"301b0c",x"3b210e",x"150e07",x"28170a",x"311c0d",x"361f0e",x"2f1b0c",x"2f1a0c",x"38200e",x"39210f",x"39200f",x"3a210f",x"37200f",x"39200f",x"472913",x"3a210f",x"412612",x"150e07",x"150e07",x"2c190c",x"2b190b",x"191008",x"221409",x"3f230f",x"3f220f",x"3b200d",x"3a1f0d",x"3e220f",x"2b180b",x"311c0c",x"3e230f",x"442712",x"3e2411",x"3e2411",x"37200f",x"361f0e",x"341d0d",x"3d2310",x"3a220f",x"361f0e",x"361f0e",x"351d0d",x"341d0d",x"462812",x"341d0d",x"321c0c",x"452711",x"452711",x"492b14",x"482a16",x"573519",x"57321a",x"58351b",x"59361c",x"56341c",x"52311a",x"472a18",x"4a2b19",x"4a2b18",x"4b2c19",x"51311c",x"482b17",x"4d2d19",x"4e2d1a",x"4c2d1a",x"50301b",x"4d2f1a",x"4c2e1a",x"4d2d17",x"4d2d18",x"502e19",x"55331a",x"56331b",x"4c2c18",x"4d2d18",x"4f2f18",x"54331c",x"502f1a",x"4f2f19",x"4a2814",x"4a2a16",x"523119",x"4e2d15",x"492913",x"452713",x"4b2b14",x"502e15",x"502d15",x"4e2c15",x"4e2d16",x"4b2b15",x"512f15",x"4d2c15",x"4f2d16",x"543016",x"563217",x"502e15",x"532e15",x"4e2d14",x"512f15",x"4f2d15",x"532f15",x"4b2c15",x"512e15",x"492913",x"512e18",x"4c2d17",x"543019",x"533119",x"4f2d18",x"52301a",x"57351c",x"56341c",x"52321b",x"58341d",x"5a371f",x"51311c",x"56341d",x"54331d",x"57351f",x"593820",x"57361d",x"56341d",x"55331d",x"51311b",x"4d2d1a",x"4b2d1a",x"4b2c19",x"482a18",x"4b2d1a",x"4b2d1a",x"52321c",x"53321d",x"50301c",x"5a361e",x"59361f",x"58371f",x"58341d",x"53311a",x"55341c",x"56331c",x"52311c",x"51321c",x"4f2e19",x"442816",x"4b2c17",x"4e2e1a",x"4e2e19",x"4c2d19",x"522f18",x"4f2e18",x"55311b",x"543119",x"512f19",x"56331a",x"5a361c",x"54321a",x"4d2e17",x"502e18",x"432613",x"412514",x"4a2c16",x"472a15",x"452914",x"422613",x"492916",x"492b15",x"4d2d17",x"4a2c16",x"4c2c16",x"502f17",x"4d2c15",x"502f17",x"512f18",x"533219",x"4c2c16",x"4a2a16",x"4f2d16",x"5a361b",x"5a361c",x"543118",x"4d2b14",x"462510",x"4b2b14",x"492a13",x"4d2b13",x"482711",x"442511",x"492913",x"472813",x"4c2b14",x"4e2d14",x"4d2d15",x"4e2e16",x"4c2b14",x"4a2b14",x"502d15",x"4f2d15",x"4a2b14",x"4c2b14",x"4c2a14",x"4d2c14",x"4d2c15",x"4a2913",x"4a2a13",x"492a13",x"472711",x"4a2912",x"4a2913",x"432611",x"472913",x"472913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231509",x"241609",x"231509",x"231509",x"221409",x"221509",x"221409",x"221409",x"462711",x"462711",x"1d1108",x"38200e",x"1f1209",x"1e1209",x"1d1108",x"211408",x"271709",x"251609",x"291909",x"2e1c0b",x"2d1c0b",x"2f1c0b",x"3a210d",x"3a220d",x"3f250e",x"3c230e",x"412711",x"492b13",x"462812",x"2c221b",x"1b1108",x"170f07",x"462a14",x"462a14",x"221409",x"221409",x"201309",x"201309",x"201309",x"211309",x"27170a",x"2f1b0c",x"442915",x"3e3127",x"43382e",x"483e34",x"4a4036",x"26170a",x"261609",x"321c0d",x"472811",x"422f22",x"4e4035",x"4c3e33",x"514236",x"3a200e",x"201309",x"201309",x"201309",x"201309",x"231509",x"211409",x"28180a",x"28180a",x"2a190a",x"251509",x"27170a",x"23150a",x"221409",x"3f2814",x"3f2814",x"211409",x"1f1309",x"1e1208",x"1d1208",x"26160a",x"3f2410",x"4a2c15",x"1e1209",x"211409",x"201309",x"201309",x"201409",x"211409",x"221409",x"1f1208",x"1f1208",x"1f1208",x"1f1209",x"2d190b",x"3a200d",x"221409",x"221409",x"251609",x"251609",x"2d1b0a",x"29180a",x"29180a",x"2d1c0a",x"321e0b",x"2e1c0a",x"2b1a0b",x"2e1c0a",x"28180a",x"28180a",x"402511",x"351d0e",x"231509",x"231409",x"27180a",x"29190a",x"29190a",x"29190a",x"27170a",x"28180a",x"251609",x"241509",x"231509",x"221409",x"201308",x"1e1208",x"1e1209",x"442611",x"201309",x"221409",x"23150a",x"24150a",x"24150a",x"231409",x"231509",x"24150a",x"231509",x"231509",x"221409",x"221409",x"3e342c",x"41372e",x"463c33",x"423930",x"26150a",x"211309",x"231409",x"251509",x"261609",x"2a1a0a",x"2b1a0b",x"2b1a0a",x"2b1a0a",x"2b1a0a",x"2c1a0a",x"321d0b",x"301b0c",x"381f0e",x"311d0e",x"4a3f35",x"3a322a",x"322a22",x"402510",x"4a3423",x"473d34",x"4d3f34",x"4f4338",x"4f4338",x"4f4338",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1a1008",x"241509",x"150e07",x"4b2b14",x"311c0c",x"4e2d15",x"150e07",x"150e07",x"28180b",x"24150a",x"150e07",x"3a210f",x"2a190b",x"150e07",x"150e07",x"150e07",x"462711",x"1f1309",x"150e07",x"150e07",x"25160a",x"211409",x"2c190b",x"28170a",x"2a180b",x"4f2d15",x"150e07",x"221409",x"311c0d",x"29180b",x"2d190b",x"2b180b",x"331c0c",x"2d180b",x"301a0b",x"311a0b",x"301a0b",x"241509",x"422510",x"381f0e",x"3d220f",x"150e07",x"150e07",x"24150a",x"24150a",x"180f07",x"4a2b14",x"361e0d",x"150e07",x"150e07",x"180f08",x"3a210f",x"1c1108",x"190f08",x"412411",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"412410",x"341e0d",x"351e0d",x"452711",x"452711",x"462a15",x"462a16",x"4b2d16",x"4f2f17",x"4c2d18",x"492b18",x"512f1a",x"502f1a",x"55341c",x"5c361e",x"56331c",x"4d2f1b",x"54331c",x"54331c",x"4e301b",x"55341d",x"4b2e1a",x"4b2d18",x"492d18",x"482b18",x"4f2f1b",x"4e2f18",x"492b17",x"54321a",x"4b2d18",x"4d2e19",x"50301b",x"52311a",x"4d2f1a",x"50311a",x"452a16",x"432714",x"4b2c17",x"4b2d18",x"492c17",x"4c2d16",x"513018",x"533218",x"523218",x"4f2f17",x"4b2b14",x"4f2e16",x"4b2c15",x"4f2f16",x"502f17",x"472913",x"462712",x"402410",x"4d2c15",x"502e16",x"4c2c14",x"4f2d14",x"472712",x"4b2b14",x"472912",x"4c2d15",x"4b2c15",x"59351a",x"4b2c16",x"4d2e16",x"4a2b17",x"452815",x"492a16",x"422715",x"432715",x"452815",x"452916",x"462a18",x"4b2d1a",x"50301b",x"4c2d1a",x"52321c",x"4f301c",x"55341d",x"52331d",x"50311d",x"56341e",x"52331e",x"4b2e1b",x"4d2f1b",x"50301c",x"4d2f1b",x"51311b",x"4c2e1a",x"4b2e1b",x"472c19",x"492c1a",x"4b2d1a",x"51301c",x"58341c",x"4e301b",x"51301a",x"53331d",x"53321c",x"462b19",x"482c19",x"4b2d19",x"4a2b17",x"492c18",x"4a2c18",x"462a17",x"51311b",x"52311a",x"51311a",x"53321b",x"4e2e19",x"4b2c16",x"452814",x"533018",x"482916",x"472a16",x"442816",x"492a17",x"553219",x"4b2d16",x"492c17",x"4a2c17",x"503119",x"492c18",x"492b17",x"472a15",x"482a16",x"523018",x"503018",x"4c2c15",x"482914",x"502f18",x"512f17",x"543319",x"553219",x"543219",x"513118",x"4e2f17",x"4a2b14",x"492812",x"523018",x"543117",x"583217",x"553218",x"4b2c14",x"533117",x"533118",x"442712",x"4d2d15",x"442712",x"4d2d16",x"4c2d16",x"4a2b14",x"472812",x"482812",x"492913",x"502e16",x"4a2a14",x"482912",x"462711",x"482a13",x"472812",x"432611",x"3f2410",x"412511",x"412511",x"2d1a0c",x"4a2913",x"4c2b14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"241509",x"241509",x"221408",x"221409",x"201309",x"241509",x"241509",x"29180b",x"3c220f",x"1d1108",x"1d1108",x"1d1208",x"1f1309",x"1f1309",x"231509",x"231509",x"26160a",x"2b190b",x"37200d",x"3d240e",x"3f260f",x"3f250e",x"3d240e",x"3b220d",x"3f250e",x"3c230e",x"472912",x"482914",x"432611",x"402511",x"191008",x"1e1208",x"1d1208",x"412511",x"2f1b0c",x"241509",x"301c0c",x"351e0e",x"25150a",x"221409",x"201309",x"25150a",x"422510",x"3d3127",x"463c33",x"554538",x"59493d",x"000000",x"351d0d",x"351d0d",x"211409",x"463122",x"504134",x"56483c",x"574b40",x"2f1b0c",x"201309",x"211409",x"211409",x"221409",x"231509",x"211409",x"24150a",x"27170a",x"29180a",x"27170a",x"26170a",x"24160a",x"221409",x"442712",x"4d2e16",x"211409",x"201309",x"201309",x"201409",x"191008",x"3d2310",x"3b2210",x"1e1208",x"201309",x"27170a",x"24150a",x"201409",x"211409",x"221409",x"211409",x"231409",x"23150a",x"231409",x"221409",x"3d200d",x"432510",x"221409",x"251609",x"1c1108",x"2b190b",x"201309",x"2e1c0b",x"2c1b0b",x"2d1c0b",x"28190a",x"281809",x"261609",x"211408",x"241409",x"191007",x"422d1e",x"201309",x"201309",x"261609",x"27170a",x"28180a",x"2a1a0b",x"27170a",x"2c1b0a",x"29190a",x"27180a",x"241609",x"25160a",x"25160a",x"201409",x"1f1209",x"24150a",x"201309",x"1f1208",x"1f1208",x"211309",x"211409",x"231509",x"221409",x"23150a",x"24150a",x"221409",x"201309",x"23150a",x"433931",x"3d332a",x"372e25",x"2b2119",x"381f0e",x"2c190b",x"331e0e",x"321d0d",x"341e0c",x"351f0d",x"321c0b",x"321c0c",x"331d0c",x"321d0b",x"3d240f",x"412610",x"472912",x"492a11",x"422613",x"4d4035",x"372e26",x"2f271f",x"29170a",x"452d1f",x"554539",x"4f4135",x"574b40",x"55493f",x"55493f",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"150e07",x"4b2b14",x"3b2210",x"150e07",x"1f1309",x"321c0d",x"321d0d",x"2a190b",x"231409",x"311b0c",x"3f2411",x"3e2411",x"442712",x"3a210f",x"150e07",x"150e07",x"1b1108",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a200e",x"150e07",x"150e07",x"25150a",x"26160a",x"2d1a0b",x"331d0d",x"311b0c",x"311b0b",x"341d0c",x"341d0d",x"361f0e",x"2b190b",x"412611",x"412511",x"150e07",x"4b2c15",x"150e07",x"150e07",x"351e0d",x"351e0d",x"150e07",x"150e07",x"28170a",x"28170a",x"231509",x"1c1108",x"482a13",x"180f08",x"150e07",x"150e07",x"28180b",x"28180b",x"2e1a0c",x"2b190c",x"2f1b0d",x"321d0d",x"2e1a0b",x"29180b",x"27170a",x"301c0d",x"2f1c0d",x"4b2b15",x"371e0e",x"331c0d",x"442712",x"442712",x"472a16",x"472b16",x"3a2313",x"4e2f18",x"4d2d17",x"4d2e1a",x"4f2e18",x"57321b",x"51311b",x"5c371d",x"5c381e",x"57351c",x"4f311b",x"4f301a",x"402817",x"4d301b",x"4f311b",x"57361d",x"472d1a",x"432a18",x"56341c",x"51321c",x"50301b",x"51301a",x"472c18",x"4d2f1b",x"4f301b",x"53321c",x"492d19",x"4b2e19",x"4d2f19",x"51301a",x"4b2d17",x"4e2d17",x"452915",x"4b2c16",x"4a2b16",x"4c2d16",x"432714",x"452915",x"422611",x"40220f",x"422511",x"492a14",x"4a2b14",x"482913",x"482813",x"482913",x"4a2b13",x"4c2b14",x"4f2c15",x"492a13",x"4b2a14",x"452812",x"432712",x"472814",x"422512",x"482813",x"4b2c15",x"402513",x"412615",x"422714",x"492c18",x"472a17",x"422615",x"452918",x"492c19",x"4d2e1b",x"492d1a",x"4a2e1b",x"4d301c",x"50321c",x"4b2f1a",x"50311d",x"51311d",x"492e1c",x"4d2f1c",x"482d1a",x"432a19",x"4a2d1b",x"4b2d1b",x"4b2e1b",x"472c1a",x"4d301c",x"5c3921",x"52331d",x"5e3a20",x"53341e",x"5a371f",x"4f311c",x"50321c",x"55331d",x"452918",x"442918",x"56341c",x"4a2d1a",x"4e301c",x"4f311c",x"452b17",x"4b2d18",x"432816",x"3d2515",x"432816",x"472a17",x"53301a",x"4b2d18",x"4e2e19",x"4d2e17",x"5a341a",x"4d2d17",x"442815",x"462a17",x"4c2d18",x"492b17",x"4e2e18",x"472a16",x"4e2f18",x"4f2f19",x"492c17",x"4f2f19",x"472b17",x"492c17",x"4c2e18",x"54311a",x"4d2d17",x"472b16",x"503118",x"58341a",x"4c2e18",x"513019",x"523017",x"56351a",x"503018",x"533219",x"513017",x"563118",x"512f16",x"593419",x"583318",x"522e16",x"482a13",x"472913",x"402612",x"3f210f",x"442511",x"512e16",x"462913",x"432611",x"4e2d15",x"472912",x"4a2a13",x"4d2c15",x"402511",x"412511",x"462812",x"4d2c14",x"3d230f",x"3d220f",x"3f230f",x"40240f",x"311b0c",x"3b220f",x"472812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26170a",x"211409",x"221409",x"221409",x"231509",x"221409",x"23150a",x"22150a",x"221509",x"221509",x"1d1108",x"1d1108",x"1f1309",x"251509",x"2d1a0c",x"311c0c",x"341f0d",x"301c0c",x"37200d",x"3d240e",x"3f260f",x"3f250e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462913",x"3c2310",x"2f1c0c",x"241609",x"1d1208",x"3b220f",x"37200e",x"2a190b",x"251609",x"231509",x"221409",x"211409",x"201309",x"261408",x"371f0e",x"3b2c22",x"483a2f",x"4f4237",x"554538",x"000000",x"361d0d",x"361d0d",x"432713",x"4c3221",x"57493d",x"5c4e42",x"584a3e",x"402410",x"231509",x"221509",x"231409",x"24150a",x"25160a",x"24150a",x"25160a",x"28180a",x"27170a",x"28180a",x"25160a",x"25160a",x"23150a",x"1f1208",x"3d2311",x"221509",x"211409",x"211409",x"211309",x"201309",x"311b0c",x"2f1b0c",x"201309",x"1e1108",x"201309",x"1f1208",x"221409",x"231509",x"221509",x"231509",x"231509",x"231509",x"221409",x"221409",x"2a190b",x"3b200d",x"1a1008",x"1c1108",x"1c1108",x"1c1108",x"331c0c",x"331c0c",x"2c1b0b",x"2a190b",x"281809",x"29190a",x"241609",x"26170a",x"251609",x"191008",x"27170b",x"190f07",x"23150a",x"26160a",x"261709",x"2a190a",x"2f1c0b",x"2d1b0a",x"2c1a0a",x"26170a",x"2b1a0a",x"24160a",x"241509",x"211409",x"221509",x"1f1309",x"201409",x"26160a",x"432712",x"422712",x"361f0f",x"351f0e",x"2d1b0c",x"27170b",x"23150a",x"221409",x"28170b",x"25160a",x"25160a",x"25160a",x"3a3128",x"2c221a",x"1d1108",x"201409",x"27160a",x"27160a",x"231509",x"25150a",x"26160a",x"24150a",x"241509",x"231509",x"29180a",x"2f1c0b",x"311d0b",x"351f0d",x"442811",x"3c2210",x"4b3c30",x"2c241c",x"211811",x"4b2d16",x"4e3321",x"4c4036",x"55473b",x"55473c",x"53463b",x"53463b",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"28170b",x"150e07",x"321d0d",x"341e0e",x"311c0d",x"2c1a0c",x"231409",x"241409",x"211308",x"301a0b",x"39200e",x"402410",x"422411",x"3a1f0e",x"321c0c",x"301a0b",x"341c0c",x"3c200e",x"3e210f",x"2d190b",x"150e07",x"150e07",x"432510",x"150e07",x"150e07",x"150e07",x"29180b",x"351f0f",x"371f0e",x"321c0d",x"3d2310",x"3e2411",x"3c2311",x"2e1b0d",x"472a14",x"150e07",x"150e07",x"2c1a0c",x"150e07",x"37200f",x"150e07",x"150e07",x"201309",x"29170b",x"27160a",x"211309",x"28170a",x"211309",x"2d190b",x"150e07",x"150e07",x"241509",x"241509",x"2d190b",x"2c190b",x"2d1a0b",x"2b180b",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"281609",x"2e1a0b",x"2c190b",x"482812",x"351d0d",x"361f0e",x"422511",x"422511",x"422511",x"3a2313",x"392314",x"392413",x"3e2716",x"452a17",x"422717",x"482d1a",x"56341d",x"55341d",x"58361d",x"58361f",x"51311b",x"4f301b",x"492d1a",x"4d2f1b",x"442a17",x"442a18",x"51311c",x"4e301a",x"59361d",x"492d1a",x"54331c",x"58351d",x"4e2f1a",x"4f2f1a",x"4e2f1a",x"50301b",x"472b18",x"442916",x"432715",x"422614",x"3d2313",x"442814",x"4e2e18",x"4a2c16",x"472a15",x"503017",x"4c2d17",x"472a16",x"452813",x"412411",x"391e0d",x"3c200d",x"3e220f",x"3f2410",x"40230f",x"432511",x"3b200e",x"3b200d",x"391e0d",x"422410",x"422410",x"402311",x"442612",x"4d2b15",x"492914",x"422513",x"402513",x"472916",x"492c17",x"4e2f19",x"4b2d1a",x"452a17",x"4a2d1a",x"4b2e1b",x"4c2f1c",x"50311d",x"54351e",x"53341e",x"53341f",x"50321e",x"58371e",x"58361f",x"4e301c",x"50311c",x"52321d",x"492e1c",x"472c1a",x"4c2e1b",x"4c2e1a",x"4d2e1b",x"472c1b",x"492d1a",x"53321d",x"51311b",x"472b1a",x"52301c",x"462b19",x"492c1a",x"4b2d1b",x"492d1a",x"472c1a",x"472b19",x"482b18",x"402616",x"472b18",x"462b18",x"482b18",x"4d2d19",x"432917",x"412817",x"452918",x"4a2d1a",x"52321b",x"5b361d",x"4d2e1a",x"4e2f1a",x"482c18",x"452a18",x"482b18",x"52301a",x"4a2d19",x"462b18",x"55331d",x"472b18",x"51311b",x"4e2e19",x"4b2d19",x"4d2e19",x"513019",x"50301a",x"492a16",x"523019",x"4e2e19",x"51311a",x"4c2e18",x"4c2e19",x"4b2d18",x"4b2d17",x"54321a",x"482a14",x"402512",x"402311",x"3e220f",x"422411",x"523017",x"502f17",x"4e2d15",x"4b2c15",x"4f2e16",x"492a14",x"422611",x"3d220e",x"361c0c",x"331c0b",x"3f230f",x"482912",x"4e2b13",x"422411",x"472711",x"442510",x"3d210f",x"3c200d",x"412411",x"3f2311",x"3d2111",x"381f0f",x"371f0f",x"311c0e",x"27170b",x"432713",x"402511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"211409",x"211309",x"201309",x"1f1208",x"1f1208",x"1f1208",x"23150a",x"23150a",x"000000",x"1d1108",x"1f1309",x"251509",x"2d1a0c",x"311c0c",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231509",x"241609",x"1e1208",x"3b220f",x"37200e",x"2a190b",x"251609",x"231509",x"221409",x"211409",x"1d1007",x"2c1609",x"311c0c",x"3b271a",x"413126",x"483a2f",x"000000",x"000000",x"351d0c",x"402612",x"442813",x"503523",x"534336",x"52463c",x"564c42",x"432610",x"3a220f",x"27180a",x"2c190b",x"351e0e",x"301b0d",x"25160a",x"25150a",x"25160a",x"27170a",x"27170b",x"25150a",x"221409",x"201309",x"412411",x"211409",x"201409",x"211409",x"211409",x"201309",x"201409",x"381f0d",x"1d1208",x"1e1209",x"1e1208",x"1e1108",x"221409",x"221408",x"241609",x"231509",x"221409",x"201308",x"1f1208",x"1e1108",x"1f1208",x"26150a",x"3d220f",x"1d1108",x"1b1008",x"1b1108",x"1c1108",x"2f1a0b",x"2f1a0b",x"000000",x"000000",x"000000",x"26170a",x"25160a",x"26170a",x"251609",x"000000",x"190f07",x"1e1208",x"24160a",x"28170a",x"27170a",x"2c1a0b",x"2c1a0b",x"2c1b0a",x"2f1c0b",x"28180a",x"2a190a",x"25160a",x"241509",x"211409",x"221509",x"000000",x"201309",x"201309",x"24150a",x"29180b",x"201309",x"27170a",x"24160a",x"27170b",x"23150a",x"221409",x"211409",x"201309",x"1f1208",x"1f1208",x"2d231b",x"271d15",x"311c0c",x"2c190b",x"29180b",x"2b180b",x"25160a",x"27170a",x"27170a",x"27170a",x"24150a",x"24150a",x"231509",x"29180b",x"2c190b",x"37200f",x"442813",x"422611",x"473327",x"231b14",x"1a1008",x"3d220e",x"51341f",x"544032",x"4e443a",x"53483e",x"53483e",x"53483e",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"1d1208",x"412511",x"150e07",x"26160a",x"2f1a0c",x"2f1a0b",x"28170a",x"27160a",x"150e07",x"412410",x"3a200e",x"1b1108",x"150e07",x"150e07",x"170f07",x"351c0c",x"28160a",x"2d190b",x"371e0c",x"1a1008",x"150e07",x"150e07",x"221309",x"41240f",x"2b180b",x"27160a",x"321c0c",x"3d220f",x"150e07",x"25150a",x"361e0d",x"321c0c",x"331d0d",x"341d0d",x"301b0c",x"2b180b",x"432410",x"150e07",x"231409",x"211309",x"28160a",x"371f0e",x"150e07",x"150e07",x"27170b",x"29180b",x"311c0d",x"2d1a0c",x"321c0d",x"29180b",x"37200f",x"150e07",x"150e07",x"231509",x"2b180b",x"2d190b",x"321d0e",x"301c0d",x"311d0d",x"361f0e",x"36200f",x"331e0e",x"321d0d",x"321c0d",x"311b0c",x"492912",x"321c0c",x"361f0e",x"150e07",x"150e07",x"150e07",x"000000",x"392413",x"352114",x"322013",x"492d19",x"4d2e19",x"51331c",x"52331c",x"53341d",x"56341d",x"5d3920",x"54351d",x"5a371f",x"56361f",x"55331c",x"472b19",x"4c2d1a",x"4f301c",x"50311c",x"53331c",x"5c371e",x"5f3a20",x"52331c",x"5b381f",x"51311b",x"56341c",x"58361d",x"4f2d19",x"57351b",x"4f2f19",x"523019",x"4a2c17",x"512f19",x"4f2e17",x"4a2c15",x"4e2d16",x"472915",x"4b2b15",x"4b2b15",x"462813",x"4d2c16",x"452713",x"422410",x"3e210e",x"3b200d",x"3e220e",x"43240f",x"3b200d",x"40220f",x"3c200d",x"41230f",x"412310",x"40220f",x"422411",x"4c2a13",x"452713",x"492a15",x"4f2d17",x"492a15",x"4a2b17",x"4a2b17",x"482c18",x"482a16",x"412717",x"4b2d19",x"492c19",x"442a18",x"472b19",x"482c1a",x"4b2d1a",x"492e1b",x"4a2d1b",x"53331d",x"54341e",x"54341e",x"57361f",x"52311d",x"52331d",x"5c3920",x"50321c",x"5d3a20",x"593620",x"55351f",x"53341f",x"4e301d",x"50301c",x"492d1c",x"50321e",x"50321d",x"50311d",x"56351e",x"56351d",x"5c3820",x"56361f",x"59371f",x"452a18",x"472a19",x"56351d",x"52341d",x"58361e",x"55331c",x"4e2f1a",x"4b2e19",x"4f2f1a",x"51311a",x"5c371d",x"54331c",x"4f301a",x"4d2f1b",x"4e311b",x"51321c",x"4d2f1a",x"50301b",x"53321d",x"54331c",x"53321b",x"51311a",x"4d2d18",x"56321a",x"53301a",x"59341d",x"5c371d",x"57331c",x"513119",x"52321b",x"55331c",x"4f301a",x"57341b",x"55331b",x"55331a",x"482a15",x"4b2c14",x"4d2e16",x"462713",x"4c2b15",x"4a2913",x"462812",x"492812",x"4f2d15",x"442611",x"452712",x"452612",x"4e2c15",x"412410",x"3e220f",x"3c200e",x"3c200e",x"3f220f",x"482711",x"462610",x"3c200d",x"42230f",x"3d200d",x"3f220e",x"3c1f0d",x"3c200d",x"442510",x"3b210e",x"321d0e",x"2c1a0c",x"27170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211409",x"211309",x"201309",x"1f1208",x"1f1208",x"1f1208",x"23150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39200e",x"29180b",x"29180b",x"453022",x"000000",x"000000",x"000000",x"000000",x"38200f",x"482a14",x"4a2b15",x"1f1309",x"1f130b",x"3c322b",x"482a13",x"3b220e",x"2e1b0b",x"231509",x"25160a",x"24150a",x"25160a",x"25160a",x"2a1a0b",x"28180b",x"27170b",x"231509",x"211409",x"221409",x"412512",x"211409",x"211409",x"211409",x"201309",x"201309",x"231509",x"452712",x"221409",x"1f1209",x"211409",x"211409",x"231409",x"241609",x"29180a",x"221509",x"201309",x"1f1208",x"1e1108",x"1f1208",x"1e1208",x"2a180a",x"3b210f",x"1d1208",x"1c1108",x"1b1108",x"1d1108",x"241509",x"361e0d",x"361e0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1208",x"24160a",x"28170a",x"27170a",x"29190a",x"2c1a0b",x"2c1b0a",x"2f1d0b",x"28180a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201309",x"24150a",x"211409",x"201309",x"27170a",x"24160a",x"000000",x"000000",x"000000",x"211409",x"1f1209",x"1f1208",x"000000",x"000000",x"1f1309",x"2f1a0c",x"2c190b",x"28170a",x"29170b",x"28170b",x"29170a",x"26160a",x"2e1b0c",x"341e0d",x"341e0e",x"321d0e",x"311b0c",x"361e0d",x"3c2310",x"442711",x"4b2b14",x"422511",x"3b200e",x"1a1008",x"24160b",x"482912",x"241609",x"20150b",x"352b22",x"53483e",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"24150a",x"180f08",x"24150a",x"150e07",x"231409",x"2a180b",x"221409",x"150e07",x"221409",x"432611",x"1a1008",x"150e07",x"180f08",x"26160a",x"25160a",x"28170a",x"150e07",x"442612",x"351e0e",x"150e07",x"150e07",x"231409",x"251408",x"221208",x"201208",x"1b1008",x"341c0c",x"341d0c",x"2c180b",x"2d190b",x"150e07",x"221409",x"2c190b",x"2b180b",x"25150a",x"231509",x"4b2a13",x"150e07",x"201309",x"311c0d",x"361f0e",x"301c0c",x"150e07",x"492813",x"150e07",x"150e07",x"180f07",x"2b190b",x"2b190b",x"2a190b",x"150e07",x"452813",x"3a2210",x"150e07",x"150e07",x"2d1a0c",x"24150a",x"26160a",x"2e1a0c",x"2b190b",x"2a180b",x"2c190b",x"2b180a",x"311b0c",x"2e1a0b",x"2d1a0b",x"4b2b14",x"351f0e",x"361f0e",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"322013",x"3a2415",x"402715",x"59371c",x"53331c",x"55341c",x"55351e",x"58381f",x"56361e",x"5b3720",x"4c2f1c",x"5a381f",x"50321d",x"53321c",x"4f2f1c",x"4f301b",x"4e2f1b",x"4b2e1a",x"4e2e1a",x"4e2e1b",x"56341c",x"5c371f",x"50301a",x"4f2f1a",x"4c2d18",x"50301a",x"4d2d17",x"502f18",x"4d2c16",x"4a2b17",x"502e17",x"543219",x"4c2c16",x"4b2c16",x"462813",x"4e2d16",x"4f2e16",x"4d2c16",x"4a2912",x"452712",x"3f2310",x"452712",x"472812",x"4c2c15",x"4a2a13",x"4b2b14",x"4f2d15",x"4c2c15",x"4f2d14",x"4b2a13",x"3d200c",x"3a1c0c",x"40230f",x"422511",x"422612",x"442713",x"4a2a15",x"452715",x"482915",x"4c2d18",x"462916",x"482c19",x"4b2e19",x"4d2e1a",x"482d19",x"4f311d",x"52331d",x"55341e",x"56351d",x"54321d",x"50311c",x"52321d",x"4b2e1b",x"4f321e",x"51331e",x"593720",x"573620",x"5c3920",x"593620",x"58361f",x"53331f",x"57361f",x"593720",x"5e3b21",x"553520",x"50331e",x"54321e",x"4f311d",x"54331d",x"4c2f1c",x"472b19",x"482b19",x"4e301c",x"4a2d1a",x"4c2e1c",x"56351d",x"50311d",x"52321d",x"4f2f1b",x"4d2f1b",x"54331c",x"54331d",x"54321c",x"4e2e1b",x"4f2f1b",x"53331c",x"51311c",x"4d2f1b",x"4c2f1a",x"53341c",x"5a3720",x"54331d",x"502f1a",x"53331c",x"52321c",x"4d2e1a",x"57331d",x"4f2e19",x"4a2b18",x"4d2d18",x"533019",x"452917",x"4f2d18",x"55331b",x"513019",x"4c2d18",x"4e2d17",x"4d2d18",x"4a2b16",x"4d2c15",x"4d2c16",x"4f2d15",x"4c2c15",x"522f15",x"4b2a13",x"4d2b14",x"472813",x"4f2d15",x"442712",x"4a2913",x"452711",x"492912",x"452713",x"422511",x"442611",x"4a2c14",x"4b2b14",x"4e2d15",x"543116",x"573318",x"4e2c14",x"4b2a13",x"3b1e0c",x"331a0a",x"34190a",x"1b1108",x"1d1108",x"321d0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2310",x"29180b",x"29180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"482a14",x"422612",x"2f1b0c",x"211409",x"1c1108",x"231a11",x"482a13",x"3b220e",x"2e1b0b",x"231509",x"25160a",x"24150a",x"29180a",x"29180a",x"26160a",x"261509",x"2c190b",x"2b180b",x"28160a",x"29170a",x"472812",x"211409",x"211409",x"211409",x"26160a",x"201309",x"211309",x"38200f",x"27170a",x"201309",x"211409",x"221409",x"241609",x"271709",x"2c1a0b",x"24160a",x"231509",x"231509",x"231509",x"231509",x"221409",x"2b180b",x"3e2411",x"1f1308",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"2d190b",x"2d190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201209",x"180e07",x"1e1108",x"1f1007",x"2d190a",x"2e1a0b",x"2f1b0c",x"2f1b0c",x"2c190b",x"311b0c",x"311b0c",x"361e0d",x"3c210f",x"442711",x"4b2b14",x"452813",x"341d0c",x"211309",x"23160b",x"37200e",x"261709",x"291a09",x"261b11",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"3d2210",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1a0b",x"492912",x"27160a",x"150e07",x"1c1108",x"241509",x"2d190b",x"2c180b",x"2e1a0b",x"301b0c",x"2b190b",x"3b210f",x"3c220f",x"150e07",x"2a180b",x"311c0d",x"351f0e",x"392110",x"37200f",x"2c1a0b",x"26160a",x"2b190c",x"3e2411",x"402511",x"412511",x"150e07",x"150e07",x"1d1208",x"3b210f",x"502d15",x"150e07",x"170f07",x"2b180b",x"2f1a0c",x"341d0d",x"311d0d",x"341e0e",x"1c1108",x"22150a",x"5b371b",x"1f1309",x"150e07",x"150e07",x"150e07",x"422712",x"191008",x"2c1a0c",x"462913",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"25160a",x"4b2b15",x"39210f",x"39210f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"402715",x"3f2615",x"3f2715",x"56331c",x"52311b",x"51311c",x"55341d",x"56341d",x"57361f",x"502f1b",x"54321c",x"58351d",x"52311d",x"492c1a",x"4c2f1b",x"56351e",x"52341e",x"58371f",x"52321c",x"5b371d",x"53321c",x"53331d",x"55331c",x"55331c",x"52301b",x"54331b",x"543119",x"512f19",x"512f19",x"512f17",x"502f18",x"4b2c16",x"472814",x"452613",x"4d2c15",x"4a2a14",x"442512",x"482811",x"4a2912",x"4b2812",x"492813",x"4d2b14",x"4a2a14",x"583217",x"4d2b14",x"4b2a13",x"4d2b13",x"4c2a13",x"4f2d15",x"573219",x"59361c",x"543319",x"4d2d16",x"513019",x"533019",x"55331c",x"58341d",x"4a2c19",x"482c19",x"4b2d19",x"4f2f1a",x"4f2e1b",x"50301b",x"51311c",x"4d2f1b",x"4b2d1b",x"502f1b",x"54321d",x"51321c",x"553620",x"563720",x"583821",x"5b3b23",x"5c3b22",x"54341f",x"52331e",x"56361f",x"5d3a23",x"583721",x"5e3b23",x"52331c",x"4e301d",x"51331f",x"563621",x"4a2e1b",x"4e2f1c",x"50321e",x"4f301d",x"4e2f1c",x"56361f",x"4f311c",x"53341f",x"56351f",x"52331e",x"56361f",x"56351f",x"51331e",x"52321d",x"593820",x"56361f",x"4e311c",x"54351e",x"59371f",x"58351e",x"57341d",x"53311d",x"4c2f1b",x"54311c",x"4e2f1c",x"52311c",x"54331d",x"53321c",x"4b2c1a",x"4f2f1b",x"4f301a",x"4b2d19",x"4d2f1a",x"4d2f1a",x"5a3720",x"5a371e",x"56331c",x"56341c",x"50301a",x"59361d",x"52311b",x"54331c",x"4b2c16",x"502f19",x"4d2d18",x"492b15",x"4d2c16",x"502e16",x"513016",x"522e16",x"4a2911",x"4b2a13",x"472811",x"492812",x"452611",x"422410",x"492912",x"422410",x"3e220f",x"442611",x"452711",x"4f2c15",x"492a13",x"512e15",x"4b2a14",x"452712",x"4c2c14",x"553219",x"513017",x"3d2411",x"341e0e",x"301c0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1b0c",x"211409",x"1c1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29180a",x"29180a",x"26160a",x"261509",x"2c190b",x"2b180b",x"28160a",x"29170a",x"221409",x"23150a",x"221409",x"221409",x"211309",x"1f1209",x"1f1208",x"1f1309",x"2f1a0c",x"3b210f",x"39200e",x"331d0d",x"241609",x"28180a",x"28180a",x"221409",x"221409",x"221409",x"221409",x"211309",x"211309",x"29180b",x"26160a",x"25170a",x"25160a",x"201309",x"1f1309",x"201309",x"3d210f",x"3d210f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"180e07",x"1e1108",x"1f1007",x"2d190a",x"2e1a0b",x"2f1b0c",x"2f1b0c",x"2c190b",x"311b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211309",x"23160b",x"37200e",x"2e1c0b",x"291a09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1e1208",x"331d0d",x"301a0b",x"361e0d",x"3e220e",x"371d0d",x"3f220e",x"1f1208",x"150e07",x"150e07",x"150e07",x"221409",x"261509",x"231409",x"261509",x"29170a",x"2e190b",x"2c190b",x"321c0c",x"150e07",x"150e07",x"29180b",x"301c0d",x"321c0d",x"331d0d",x"341d0d",x"341d0d",x"2f1b0c",x"24150a",x"361f0f",x"321e0e",x"3c2311",x"4e2c14",x"4b2a13",x"563319",x"321e0e",x"150e07",x"150e07",x"27170a",x"321d0d",x"2e1a0b",x"351e0e",x"321c0c",x"2e1a0b",x"301c0d",x"180f08",x"150e07",x"191008",x"4c2c14",x"4b2b14",x"502f17",x"422713",x"2f1c0d",x"341e0e",x"462914",x"4e2f17",x"533218",x"4e2d16",x"512f18",x"513017",x"472913",x"462711",x"482812",x"432611",x"4a2b14",x"4b2b15",x"3d2310",x"482913",x"351e0e",x"39210f",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"442a18",x"4b2c18",x"472b18",x"52321c",x"4e301b",x"4e301c",x"4e301b",x"52331d",x"50321d",x"4f301c",x"4d2f1d",x"4e2f1c",x"51331e",x"51321c",x"4e301b",x"4f301c",x"4b2d1a",x"472b19",x"4b2c19",x"4c2e19",x"4d2e19",x"4d2e1a",x"50301a",x"432715",x"442815",x"432612",x"432513",x"422513",x"442714",x"442713",x"402412",x"402412",x"402310",x"402310",x"402210",x"402310",x"3f2210",x"3d200e",x"3f210e",x"40220e",x"40220e",x"41230f",x"442510",x"462611",x"452711",x"482812",x"4a2a13",x"4d2c15",x"4c2c15",x"4b2c15",x"4c2c16",x"4b2b16",x"4d2e17",x"4e2d17",x"4f2f1a",x"52311b",x"51311a",x"4f2f1a",x"4a2c18",x"4f311c",x"55341d",x"52331d",x"50311c",x"53331e",x"4c301c",x"4d2f1b",x"4c2f1b",x"4f311d",x"4b2f1c",x"53331f",x"543520",x"53331f",x"50331f",x"52331f",x"50311e",x"553620",x"583721",x"543720",x"4f331f",x"53351f",x"583922",x"553721",x"563520",x"52341f",x"523420",x"52331f",x"4d301d",x"442a1a",x"4d2f1c",x"4e301c",x"4d311d",x"4f311d",x"4d2f1c",x"50311d",x"4f311d",x"4e301d",x"4e311d",x"4f321d",x"52341f",x"563620",x"54351f",x"4e311d",x"4e311d",x"4c311d",x"4f311c",x"4d311c",x"4e301d",x"4e301b",x"4d301c",x"50321c",x"4b2f1c",x"482d1a",x"4e301b",x"4d2e1a",x"4d301b",x"4b2e19",x"51311b",x"4c2e1a",x"4a2c18",x"472b18",x"472b17",x"492c18",x"4c2d19",x"472a16",x"4a2c18",x"3f2312",x"402412",x"3f2412",x"3d2211",x"3f2210",x"3f2210",x"422511",x"3f220f",x"3d200d",x"3d210e",x"3b1f0d",x"381d0c",x"3a1f0d",x"391f0c",x"391f0c",x"371d0c",x"3a1e0d",x"391e0d",x"3c200e",x"40240f",x"422410",x"462712",x"452611",x"462712",x"462812",x"4a2b14",x"4b2b14",x"492b14",x"472813",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"221409",x"221409",x"211309",x"211309",x"1f1208",x"1f1208",x"201309",x"2f1a0c",x"3b210f",x"39200e",x"331d0d",x"241609",x"28180a",x"221409",x"221409",x"22150a",x"24160a",x"27160a",x"28170b",x"23150a",x"2b1b0a",x"2a1a0a",x"2b1a0a",x"231509",x"201309",x"201309",x"231409",x"39200e",x"39200e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"170f07",x"341e0e",x"412511",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"40220e",x"150e07",x"150e07",x"150e07",x"26160a",x"2c190b",x"2d1a0b",x"331d0d",x"27170a",x"4b2b14",x"452712",x"150e07",x"2a180b",x"2a180b",x"2e1a0c",x"2f1b0c",x"2d1a0b",x"2a180b",x"27160a",x"3c210f",x"462711",x"462611",x"170f07",x"150e07",x"180f07",x"221409",x"180f08",x"3f230f",x"1e1208",x"150e07",x"201208",x"2b180a",x"301b0b",x"2c190b",x"2a190b",x"150e07",x"4f2f17",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"2d190b",x"1f1208",x"211309",x"150e07",x"150e07",x"150e07",x"191008",x"1d1108",x"1e1209",x"211409",x"211409",x"22150a",x"29180b",x"28180b",x"25160a",x"24150a",x"523018",x"361f0e",x"3a2210",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"24150a",x"221409",x"26160a",x"4d2f1a",x"462a19",x"53341d",x"54321d",x"57351f",x"57361d",x"54331d",x"59361f",x"5a3820",x"5b3a21",x"533620",x"53351e",x"4f331e",x"563820",x"54341e",x"55341d",x"5b3820",x"5b3920",x"5e3a20",x"593820",x"5b381f",x"59371d",x"57331b",x"513119",x"57331b",x"4f2d18",x"512e19",x"502e18",x"4b2a15",x"4a2a14",x"4b2a14",x"452713",x"422410",x"462812",x"472712",x"472611",x"4c2911",x"482811",x"4a2912",x"4c2a14",x"522f16",x"563118",x"512e15",x"4f2d15",x"522f16",x"512e15",x"4f2d15",x"4c2b14",x"4e2d16",x"4b2a14",x"4b2b15",x"4c2c16",x"4e2d17",x"4c2c17",x"4c2c16",x"492b17",x"4d2d18",x"4b2c18",x"4b2d1a",x"4f2e19",x"4f2f1a",x"4d2e1a",x"492c1a",x"442818",x"472b19",x"4c2e1a",x"50321d",x"54341f",x"573620",x"563620",x"583721",x"543420",x"593720",x"593821",x"583620",x"53331e",x"51311d",x"533320",x"55341e",x"573721",x"593820",x"563520",x"54341f",x"56351f",x"5c3a22",x"563821",x"5c3a22",x"593821",x"543520",x"53341f",x"4e321d",x"4e321f",x"543620",x"5b3922",x"593821",x"563521",x"553721",x"5b3a22",x"5b3a22",x"5d3b23",x"5c3a21",x"5a3920",x"5d3b23",x"55361f",x"56371e",x"52321d",x"53331e",x"56351e",x"563620",x"4f311d",x"563620",x"5c3a21",x"58381f",x"593820",x"4d311c",x"583820",x"58371f",x"53321c",x"57361d",x"5b391f",x"59371e",x"53321b",x"56361d",x"58351d",x"4f3119",x"513019",x"502f18",x"4e2d17",x"4c2d15",x"4e2e16",x"4b2a14",x"492812",x"472710",x"44250f",x"41220e",x"42240f",x"42240f",x"3f220e",x"3f220f",x"40230f",x"3d210f",x"432511",x"492913",x"4c2c15",x"502e16",x"4e2d15",x"512f16",x"502e15",x"4f2d14",x"4b2a14",x"4a2b15",x"523118",x"492b14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b2210",x"442812",x"462913",x"462813",x"452813",x"442711",x"432611",x"402410",x"3f2410",x"492a11",x"472910",x"4f2e13",x"3f2310",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"221409",x"211309",x"211309",x"1f1208",x"1f1208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221409",x"22150a",x"24160a",x"27160a",x"28170b",x"2e1c0b",x"2e1c0b",x"2c1a0a",x"29180a",x"231509",x"221409",x"211309",x"201309",x"211309",x"211309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"341d0d",x"28180b",x"3d2311",x"150e07",x"25150a",x"2d1a0c",x"2d1a0c",x"1b1108",x"150e07",x"2e1b0c",x"3c220f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301c0d",x"361f0e",x"38200f",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"361d0d",x"40230f",x"2b180b",x"3f230f",x"1d1108",x"150e07",x"2d190b",x"371e0d",x"311b0c",x"301b0b",x"27160a",x"3c210f",x"150e07",x"150e07",x"29180b",x"2f1b0c",x"231409",x"3e230f",x"211309",x"150e07",x"1a1008",x"25160a",x"2a180b",x"2a180a",x"2c190b",x"1c1108",x"3a200e",x"452611",x"150e07",x"25150a",x"2e1b0c",x"341e0d",x"321c0d",x"2f1a0b",x"321c0d",x"3a2110",x"351f0e",x"321d0d",x"331d0d",x"39200e",x"311c0d",x"4b2b14",x"2b180b",x"36200f",x"150e07",x"150e07",x"150e07",x"000000",x"201309",x"24150a",x"221409",x"26160a",x"2a180b",x"2e1a0b",x"432a18",x"422919",x"412a19",x"402919",x"432b1b",x"452c1a",x"4c311d",x"5d3b21",x"563620",x"482e1c",x"422a1a",x"462c1a",x"442b19",x"462c1a",x"52341e",x"56351f",x"593820",x"5a3820",x"58361e",x"5b3820",x"54311a",x"54311a",x"482a17",x"4f2d17",x"4b2b17",x"4b2e19",x"4d2f18",x"57331b",x"4f2f18",x"502f18",x"4b2c15",x"492a14",x"4a2914",x"4a2a14",x"492a14",x"502e15",x"4a2a14",x"4e2d16",x"4d2c16",x"4a2b15",x"482a13",x"4d2c15",x"462812",x"472812",x"422510",x"492812",x"492914",x"4f2c15",x"4a2914",x"4d2c15",x"492a15",x"452815",x"462815",x"3d2515",x"472a17",x"4a2d18",x"442917",x"482a18",x"482a18",x"4a2c19",x"4a2c1a",x"492c19",x"492e1c",x"4e301c",x"4e301c",x"492e1c",x"412a1a",x"3c2618",x"4a2e1c",x"4a2f1c",x"4d301d",x"4e301c",x"4b2e1b",x"55351e",x"4d301d",x"51311d",x"4c301c",x"472d1b",x"4b2e1b",x"4e321d",x"50331e",x"4a2e1c",x"492d1c",x"51331e",x"52331f",x"51331e",x"4d301e",x"482d1c",x"59361f",x"553520",x"50321d",x"4e321f",x"4c311d",x"482e1c",x"51321f",x"543520",x"4f321f",x"4e321f",x"4c311e",x"492f1b",x"4d301c",x"462b19",x"442a19",x"52321d",x"4d301c",x"432b19",x"4f321d",x"4e321e",x"593720",x"5b3a21",x"4f321d",x"55351d",x"4e2f1b",x"56341f",x"55351d",x"53321d",x"56351e",x"56361f",x"59381e",x"59381f",x"54341e",x"57361d",x"51311a",x"4f2f18",x"492914",x"4c2b15",x"4d2d16",x"523018",x"5a351b",x"512f17",x"4d2d15",x"492a13",x"412511",x"442712",x"452711",x"512f16",x"432611",x"412511",x"371f0e",x"3b220f",x"3e2411",x"3d2310",x"422612",x"472913",x"4a2a13",x"472812",x"432611",x"351d0d",x"5b361a",x"432612",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b2210",x"3b2210",x"442812",x"462913",x"462813",x"452813",x"442711",x"432611",x"402410",x"3f2410",x"492a11",x"472910",x"4f2e13",x"3f2310",x"3f2310",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e1c0b",x"2e1c0b",x"2b190a",x"251609",x"221409",x"211409",x"211409",x"201409",x"201309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231409",x"26160a",x"27160a",x"2e190b",x"150e07",x"191008",x"331d0d",x"361f0e",x"39200f",x"351e0e",x"211409",x"331d0d",x"3e2310",x"4a2b14",x"341e0d",x"2e1a0c",x"3a2210",x"412612",x"3b2210",x"341e0e",x"432712",x"4a2b15",x"3b2210",x"3c2310",x"4b2c14",x"321d0d",x"150e07",x"422510",x"2b180b",x"27160a",x"150e07",x"2f1b0c",x"38200e",x"39200e",x"3b210f",x"3c220f",x"3c220f",x"2b190b",x"4a2913",x"150e07",x"150e07",x"191008",x"4f2d16",x"402410",x"150e07",x"150e07",x"25160a",x"251509",x"2e1b0c",x"331d0d",x"38200e",x"28170a",x"2c190b",x"150e07",x"150e07",x"27160a",x"2a180b",x"331c0d",x"301a0b",x"361e0d",x"371f0e",x"361e0e",x"381f0e",x"311c0d",x"311c0c",x"361f0e",x"321d0d",x"4a2b14",x"351e0d",x"361f0e",x"150e07",x"150e07",x"150e07",x"170f07",x"1b1108",x"201309",x"221409",x"251509",x"29170a",x"2a170a",x"2d190b",x"2c190a",x"241308",x"2a1709",x"311b0b",x"321c0c",x"331c0c",x"341d0c",x"371e0d",x"39200e",x"3b210f",x"3c2210",x"3c2310",x"3b210f",x"3b210f",x"3c220f",x"3c220f",x"3b210f",x"381f0e",x"341d0d",x"301b0c",x"301b0c",x"2b180a",x"2c190b",x"301b0c",x"2e1a0b",x"2d180b",x"341d0d",x"371f0e",x"371f0e",x"39200e",x"39210f",x"39210f",x"38200f",x"371f0e",x"361f0e",x"361f0e",x"351f0e",x"341e0e",x"341e0e",x"331e0e",x"321d0e",x"321d0d",x"331d0e",x"331d0e",x"331d0d",x"341e0d",x"331d0d",x"321c0d",x"311b0c",x"301b0c",x"2f1b0c",x"2f1b0c",x"2f1a0c",x"2f1a0c",x"2f1b0c",x"301b0c",x"311c0d",x"321d0d",x"331e0d",x"331d0d",x"311c0c",x"301b0c",x"2e1b0c",x"2e1b0c",x"2c190b",x"2b190b",x"2a180b",x"29170b",x"27160a",x"27160a",x"28170a",x"2a190b",x"29170a",x"29180b",x"2c190b",x"2c190b",x"2c190b",x"2e1a0b",x"2f1a0b",x"2e190b",x"301b0c",x"321c0d",x"321d0d",x"331d0d",x"341e0d",x"341e0e",x"331d0d",x"331e0d",x"331d0d",x"331d0d",x"331d0e",x"331e0e",x"321d0d",x"321d0d",x"301c0d",x"2d1a0c",x"2b180b",x"28170a",x"26160a",x"251509",x"231409",x"201208",x"1e1208",x"180f07",x"2f1b0d",x"412e22",x"3c2a1e",x"412f22",x"412e22",x"3f2e21",x"402e22",x"3f2c1f",x"412f23",x"442e20",x"432f22",x"422e20",x"412e21",x"463123",x"453225",x"463224",x"3e2a1d",x"443023",x"453022",x"3f2d21",x"432f22",x"3a271a",x"453123",x"412b1c",x"402b1d",x"372417",x"3f291b",x"3c281c",x"3a271b",x"3b2719",x"37261a",x"39281d",x"38281c",x"35261c",x"38271d",x"372417",x"3a2a1e",x"37281d",x"3b2b20",x"382518",x"402c1f",x"3f2f24",x"54341e",x"4f2e16",x"4d2d16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"351f0f",x"2d1a0c",x"2d1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1b0b",x"2b190a",x"251609",x"221409",x"211409",x"211409",x"201409",x"201409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1c1108",x"361f0e",x"1d1208",x"3b220f",x"331c0c",x"150e07",x"26160a",x"2f1b0c",x"301b0c",x"2f1a0b",x"231509",x"2d1a0b",x"321c0c",x"331d0d",x"3a200e",x"150e07",x"412511",x"442712",x"462712",x"40230f",x"452611",x"462812",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200e",x"150e07",x"150e07",x"28170a",x"331c0d",x"341d0d",x"371f0e",x"39200e",x"38200f",x"341d0d",x"3a200f",x"25160a",x"3b210e",x"381d0c",x"150e07",x"341b0c",x"150e07",x"150e07",x"42240f",x"150e07",x"150e07",x"201208",x"261509",x"2a180a",x"27160a",x"1e1208",x"361e0d",x"43250f",x"150e07",x"1a1008",x"2a170a",x"311b0c",x"2c190b",x"29170a",x"2d190b",x"2e190b",x"2b180a",x"2c180a",x"2e190b",x"2d190b",x"2a180a",x"4b2b14",x"321c0d",x"351e0e",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1b1108",x"201309",x"241509",x"27160a",x"29170a",x"2c190b",x"2f1a0c",x"2f1a0b",x"321c0c",x"341e0d",x"341d0d",x"341d0d",x"341d0d",x"361e0d",x"381f0e",x"39200e",x"3a200f",x"3a210f",x"3c2210",x"3b2210",x"3a210f",x"39200e",x"38200f",x"371f0e",x"351e0e",x"2c180b",x"271609",x"28160a",x"2d190b",x"301b0c",x"331d0d",x"301b0c",x"331d0d",x"341d0d",x"361f0e",x"351d0d",x"341d0d",x"341d0d",x"351d0d",x"351e0d",x"341d0d",x"321c0c",x"321d0d",x"311c0d",x"2f1b0c",x"2f1b0c",x"2d190b",x"2c190b",x"2f1a0c",x"311c0d",x"2e1a0c",x"2d1a0b",x"2c190b",x"2c190b",x"2b180b",x"2c180b",x"2b180b",x"2a180a",x"2b180b",x"2c190b",x"2e1a0c",x"2f1b0c",x"311c0c",x"321c0d",x"311c0c",x"301b0c",x"2c180a",x"281609",x"281509",x"281609",x"28160a",x"271609",x"27160a",x"261509",x"251509",x"261509",x"27160a",x"261509",x"261509",x"26150a",x"27160a",x"27160a",x"29170a",x"2a180b",x"2b180b",x"2b190b",x"2a180a",x"2a170a",x"2a170a",x"2a170a",x"29170a",x"29170a",x"2d190b",x"2e1a0b",x"2f1a0c",x"301c0d",x"311c0d",x"311c0d",x"301c0d",x"301c0d",x"2d1a0c",x"2c190b",x"2b190b",x"2b190b",x"29180b",x"26160a",x"231409",x"211309",x"1e1208",x"1a1008",x"39200f",x"39200f",x"3c2a1e",x"412f22",x"412e22",x"3f2e21",x"402e22",x"3f2c1f",x"412f23",x"442e20",x"432f22",x"422e20",x"412e21",x"463123",x"453225",x"463224",x"3e2a1d",x"443023",x"453022",x"3f2d21",x"432f22",x"3a271a",x"453123",x"412b1c",x"402b1d",x"372417",x"3f291b",x"3c281c",x"3a271b",x"3b2719",x"37261a",x"39281d",x"38281c",x"35261c",x"38271d",x"372417",x"3a2a1e",x"37281d",x"3b2b20",x"382518",x"402c1f",x"3f2f24",x"54341e",x"54341e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f08",x"1a1008",x"1b1008",x"1c1108",x"1d1208",x"1e1208",x"1e1208",x"1f1209",x"201309",x"1f1309",x"1f1209",x"1e1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"201309",x"201309",x"201409",x"201309",x"201309",x"201309",x"1f1309",x"201309",x"201309",x"201309",x"1f1209",x"1d1208",x"1c1208",x"1c1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"190f08",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"180f07",x"191008",x"1a1008",x"191008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1209",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f08",x"191008",x"191008",x"1a1008",x"191008",x"190f08",x"180f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201409",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211309",x"2f1c0d",x"221409",x"492912",x"150e07",x"150e07",x"150e07",x"29170a",x"29170a",x"271609",x"241409",x"391f0e",x"3e220f",x"341d0c",x"371e0d",x"42240f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1e1208",x"27170a",x"1c1108",x"492913",x"150e07",x"1f1309",x"2f1b0c",x"341d0d",x"39210f",x"3b220f",x"3a210f",x"3e2310",x"3a210f",x"3a220f",x"361f0e",x"311c0d",x"482a14",x"3a200e",x"29170a",x"1f1208",x"150e07",x"1f1309",x"150e07",x"462812",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"442711",x"1c1108",x"150e07",x"150e07",x"150e07",x"1f1309",x"150e07",x"25160a",x"211409",x"28180b",x"27180b",x"26160a",x"25160a",x"191008",x"201309",x"4a2b14",x"331e0d",x"311c0c",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"170f07",x"1a1108",x"1f1309",x"23150a",x"27170a",x"2a180b",x"2c190b",x"2c190b",x"2c190b",x"2b190b",x"2d1a0b",x"2e1a0b",x"2e1a0b",x"2f1a0b",x"301b0c",x"321c0c",x"311c0c",x"321c0c",x"321c0c",x"311b0c",x"331c0c",x"2e1a0b",x"2d190b",x"2b180b",x"2b180b",x"2a180b",x"26160a",x"261609",x"251509",x"2a180a",x"2c190b",x"2c190b",x"2b180a",x"301a0c",x"321c0c",x"321c0c",x"2f1a0b",x"2c180a",x"301b0c",x"2f1a0b",x"2f1a0b",x"2d190b",x"2c190b",x"29170a",x"2a170a",x"2b180b",x"2a180b",x"2b180b",x"2b190b",x"2b180b",x"29170a",x"29170a",x"29180b",x"2a180b",x"2a180b",x"2a180b",x"2b190b",x"2b190b",x"2c190b",x"2c190b",x"2d1a0b",x"2e1a0c",x"311c0d",x"321d0d",x"331d0d",x"341e0e",x"341d0d",x"2f1a0b",x"2e1a0b",x"2e1a0c",x"2d190b",x"2f1b0c",x"2d1a0c",x"2b190b",x"2b190b",x"2a180b",x"28160a",x"26150a",x"241509",x"25150a",x"25160a",x"28180b",x"29180b",x"29190c",x"29190b",x"2a190b",x"2b190b",x"2c190c",x"2b1a0c",x"2d1a0c",x"2d1b0c",x"2c1a0c",x"2c1a0c",x"2c1a0b",x"2c1a0c",x"2d1a0c",x"2e1b0d",x"2c1a0c",x"2b190b",x"2b190b",x"2c1a0c",x"29180b",x"2a190b",x"2b190c",x"28180b",x"26160a",x"23150a",x"201309",x"1d1208",x"191008",x"331d0e",x"331d0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f08",x"1a1008",x"1b1008",x"1c1108",x"1d1208",x"1e1208",x"1e1208",x"1f1209",x"201309",x"1f1309",x"1f1209",x"1e1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"201309",x"201309",x"201409",x"201309",x"201309",x"201309",x"1f1309",x"201309",x"201309",x"201309",x"1f1209",x"1d1208",x"1c1208",x"1c1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"190f08",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"180f07",x"191008",x"1a1008",x"191008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1e1209",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f08",x"191008",x"191008",x"1a1008",x"191008",x"190f08",x"180f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"27170b",x"1d1208",x"1d1208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"361f0f",x"241509",x"462712",x"3b200e",x"351d0d",x"1d1208",x"150e07",x"180f07",x"150e07",x"1f1208",x"150e07",x"150e07",x"150e07",x"1c1108",x"1e1208",x"2f1b0b",x"4b2b13",x"150e07",x"150e07",x"1f1208",x"28170a",x"2d1a0b",x"2c190b",x"2f1b0c",x"442611",x"150e07",x"28170a",x"341d0d",x"331d0d",x"381f0e",x"3c2310",x"3c2310",x"39200f",x"351e0e",x"3a2210",x"371f0e",x"331c0d",x"442711",x"381f0e",x"442711",x"150e07",x"150e07",x"29180a",x"2c190b",x"150e07",x"2c190b",x"4c2b14",x"4c2c14",x"38200f",x"38200f",x"3a200e",x"241509",x"2a180a",x"3e230f",x"412310",x"2c190b",x"28170a",x"2b180b",x"2d1a0b",x"2a180b",x"2a180b",x"321d0d",x"341e0e",x"2f1c0d",x"311c0c",x"311c0d",x"412611",x"341d0c",x"2f1a0b",x"150e07",x"150e07",x"38200e",x"2d190b",x"22150a",x"201409",x"201309",x"29180b",x"26160a",x"2d1a0c",x"2a180b",x"2f1a0c",x"2d190b",x"2e1b0c",x"311c0d",x"331e0e",x"351e0e",x"38200f",x"362210",x"3a2210",x"392110",x"3b2311",x"361f0e",x"351e0e",x"341d0d",x"311b0c",x"311b0c",x"351f0e",x"321d0d",x"311c0d",x"28160a",x"2a180a",x"2e1a0c",x"2b180b",x"2d1a0b",x"321d0d",x"301b0c",x"311b0b",x"341d0d",x"371f0e",x"361f0e",x"38200e",x"361e0d",x"331c0d",x"321b0c",x"331c0d",x"331c0c",x"301b0c",x"341d0d",x"2f1a0c",x"301b0c",x"2c190b",x"2a170a",x"29170a",x"2b180b",x"2a170a",x"2c190b",x"2b190b",x"2a180b",x"2e1a0c",x"2d1a0b",x"2d1a0b",x"2c190b",x"311c0d",x"321d0d",x"341e0e",x"311c0c",x"311c0c",x"361f0e",x"351e0d",x"341d0d",x"341d0d",x"351d0d",x"321c0c",x"321c0c",x"341d0d",x"301b0c",x"2f1a0c",x"311c0d",x"2e1a0b",x"311c0d",x"311d0d",x"301c0d",x"2b190b",x"2a180b",x"241509",x"29170b",x"231409",x"27160a",x"27160a",x"26160a",x"28170a",x"29180b",x"2b180b",x"2d1a0b",x"2c190b",x"321d0d",x"2d1a0c",x"2e1b0c",x"301c0d",x"2f1b0c",x"301c0d",x"311c0d",x"2d1a0c",x"2a180b",x"27170b",x"2a1b0c",x"28170b",x"2a190b",x"2d1a0c",x"231509",x"27170a",x"241509",x"201309",x"231409",x"412512",x"412512",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"191008",x"1b1008",x"1b1108",x"1d1108",x"1e1208",x"1e1208",x"1f1309",x"1f1309",x"201409",x"201309",x"1f1208",x"1e1208",x"1e1208",x"1f1309",x"1e1208",x"1e1208",x"1f1208",x"1f1209",x"1f1209",x"1f1209",x"201309",x"211409",x"201409",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1209",x"1d1208",x"1c1208",x"1c1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"191008",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"180f07",x"191008",x"1a1008",x"191008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1f1209",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f08",x"191008",x"191008",x"1a1008",x"191008",x"190f08",x"180f07",x"180f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211309",x"341f0e",x"1e1208",x"3f230f",x"381f0d",x"2e1a0b",x"3b210f",x"3b210e",x"351e0d",x"361d0c",x"42220f",x"150e07",x"221309",x"2d190b",x"341d0d",x"371f0e",x"2a180a",x"180f07",x"3e220f",x"27160a",x"150e07",x"211409",x"2f1b0c",x"2e1b0c",x"2b190b",x"3f2310",x"150e07",x"2b190c",x"351f0e",x"341e0d",x"341d0d",x"361e0d",x"341d0d",x"321b0c",x"2e190b",x"2e1a0b",x"331c0c",x"2c180b",x"472812",x"341e0d",x"432712",x"150e07",x"150e07",x"211309",x"221409",x"150e07",x"3a200f",x"422410",x"150e07",x"150e07",x"201309",x"371f0e",x"150e07",x"1b1008",x"3b200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3c220f",x"351d0c",x"251509",x"150e07",x"150e07",x"3c220f",x"3a220f",x"311c0d",x"351d0d",x"361e0d",x"331c0c",x"351d0d",x"38200e",x"3a210f",x"3b2210",x"3c2210",x"3b2210",x"3f2411",x"3d2411",x"432712",x"432713",x"422713",x"3b210f",x"422612",x"3f2310",x"3b210f",x"3d2310",x"3c210f",x"3d220f",x"3a200e",x"3b210f",x"391f0e",x"391f0e",x"331c0c",x"361e0d",x"381f0e",x"39200e",x"39200e",x"371f0d",x"381f0e",x"381f0d",x"3a200e",x"381f0e",x"371e0d",x"371e0c",x"321a0b",x"351d0c",x"331b0b",x"3b210f",x"3b210f",x"3b200e",x"3a200e",x"3c210f",x"3a200e",x"341d0d",x"371e0d",x"381f0e",x"3b210f",x"3d2310",x"3b2210",x"381f0e",x"371f0e",x"3e2310",x"3d2310",x"3b2210",x"3b210f",x"39200e",x"39200e",x"371e0d",x"351d0c",x"371e0d",x"3a200e",x"3c210f",x"3e2310",x"402511",x"412511",x"3f2411",x"3c210f",x"3b200e",x"3a200e",x"371e0d",x"381f0e",x"3a200e",x"3e2311",x"3d2211",x"3b2211",x"3c2311",x"3f2514",x"361f10",x"331d0f",x"361f11",x"382213",x"3b2314",x"392313",x"3a2413",x"382213",x"382213",x"3e2514",x"3c2514",x"3c2514",x"3d2514",x"3e2614",x"362012",x"3c2414",x"3d2615",x"402715",x"3c2515",x"3a2414",x"382213",x"3b2312",x"3b2312",x"382111",x"372011",x"371f10",x"351e0f",x"372010",x"3a2211",x"37200e",x"4b2a14",x"4b2a14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1f1209",x"201309",x"201309",x"211409",x"1f1209",x"1d1108",x"1e1108",x"1f1208",x"201309",x"1f1209",x"201309",x"1f1209",x"1f1209",x"201309",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1309",x"1f1309",x"201309",x"201309",x"1f1309",x"1f1309",x"1e1209",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1b1008",x"1a1008",x"1a1008",x"191008",x"181008",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f08",x"190f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1008",x"1b1008",x"1b1108",x"1c1108",x"1d1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1e1208",x"1f1208",x"1f1209",x"201309",x"1f1309",x"1f1209",x"1f1209",x"1f1309",x"1f1309",x"1e1209",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"190f08",x"180f08",x"190f08",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"190f07",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"170f07",x"321d0d",x"1d1208",x"472812",x"311b0c",x"3f2410",x"2c1a0b",x"371f0e",x"150e07",x"150e07",x"2c1a0c",x"150e07",x"26160a",x"351e0d",x"351e0d",x"351d0d",x"361e0d",x"2f1b0c",x"26160a",x"2f1c0d",x"4e2e16",x"150e07",x"150e07",x"2a190b",x"2c1a0c",x"513017",x"150e07",x"1f1309",x"2f1c0d",x"321c0c",x"361f0e",x"351e0e",x"321c0c",x"341d0d",x"321c0d",x"331d0d",x"38200e",x"29180b",x"361f0e",x"3c2210",x"2e1a0c",x"301b0c",x"150e07",x"150e07",x"341e0d",x"492a14",x"150e07",x"150e07",x"201309",x"28170a",x"221409",x"150e07",x"422611",x"150e07",x"150e07",x"150e07",x"26160a",x"28170a",x"2e1a0c",x"2c190b",x"2c190b",x"301b0c",x"2d190b",x"301a0b",x"2f1a0b",x"2c190b",x"241509",x"3c210e",x"2a180a",x"301b0b",x"150e07",x"150e07",x"502e15",x"472712",x"442611",x"482913",x"4a2b14",x"4a2b14",x"472913",x"472913",x"472813",x"432511",x"422510",x"452711",x"452612",x"442611",x"452711",x"482913",x"472812",x"492a14",x"4c2c15",x"4b2b14",x"4c2d16",x"4c2c15",x"4b2c15",x"492913",x"432511",x"432510",x"422410",x"442611",x"462712",x"422410",x"4b2b14",x"492913",x"4b2b14",x"492a14",x"422410",x"472812",x"4a2a14",x"4a2a14",x"472813",x"472913",x"492a14",x"4a2b15",x"4d2c15",x"472812",x"432711",x"452611",x"442511",x"482812",x"482913",x"492b15",x"4c2c15",x"4d2d16",x"4a2b15",x"4a2c15",x"4e2e17",x"4f2f17",x"4d2d16",x"4b2c15",x"4b2c15",x"482913",x"462813",x"472813",x"452712",x"432511",x"422511",x"432511",x"482913",x"4b2b14",x"4c2c14",x"4b2b14",x"462712",x"452711",x"472913",x"482913",x"4a2c15",x"4c2d16",x"4b2c15",x"462813",x"4b2d17",x"482a16",x"4a2d17",x"4a2c18",x"4c2e19",x"472b18",x"4c2e19",x"4d2f1b",x"472c19",x"4a2d19",x"472b18",x"4a2d19",x"472b18",x"492d1b",x"432917",x"422818",x"452918",x"452b19",x"432918",x"422818",x"472b19",x"442918",x"442919",x"422716",x"432918",x"452a18",x"482b18",x"492d19",x"4c2d19",x"482c18",x"482d19",x"482b17",x"462b17",x"452815",x"412613",x"4c2c16",x"4c2c16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1108",x"1d1208",x"1e1209",x"1f1309",x"201309",x"201309",x"201409",x"201309",x"211409",x"211409",x"211409",x"221409",x"221409",x"221409",x"211409",x"1f1209",x"201309",x"201309",x"201309",x"201309",x"1e1208",x"1e1208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1208",x"1d1208",x"1d1208",x"1d1208",x"1d1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"180f08",x"180f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1208",x"1e1209",x"1f1309",x"201309",x"1f1309",x"1e1209",x"1f1209",x"1f1208",x"1e1208",x"1f1309",x"201309",x"201409",x"201309",x"201309",x"201409",x"211409",x"211409",x"211409",x"211409",x"201409",x"201309",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1e130b",x"1e130a",x"1c1108",x"1b1108",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"1e1208",x"1e1208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"24150a",x"311c0d",x"201309",x"442611",x"27160a",x"341d0d",x"472913",x"150e07",x"221409",x"28170a",x"361f0e",x"150e07",x"2b190b",x"371f0e",x"371f0e",x"38200e",x"39200f",x"3a2110",x"3a2210",x"2d1b0c",x"211409",x"492c15",x"2d1b0d",x"150e07",x"150e07",x"351e0d",x"3a2110",x"150e07",x"1e1209",x"2d1a0c",x"331d0d",x"341d0d",x"301b0c",x"371f0e",x"321c0c",x"311b0c",x"2b180b",x"211409",x"341d0d",x"452711",x"1e1208",x"3a200e",x"150e07",x"2c190b",x"150e07",x"150e07",x"1e1208",x"2a180b",x"2a180b",x"2f1b0c",x"2e1a0c",x"231509",x"341d0e",x"26160a",x"150e07",x"25150a",x"2c190b",x"2e1a0c",x"341d0d",x"331d0d",x"321c0c",x"321c0d",x"351d0d",x"341d0d",x"361f0e",x"311c0c",x"2a180b",x"3f2310",x"2b180a",x"281609",x"150e07",x"150e07",x"3e2310",x"543118",x"533017",x"523018",x"4e2d15",x"512e15",x"543117",x"543118",x"522f16",x"4e2c15",x"492912",x"4c2b14",x"512f17",x"553218",x"543117",x"4e2d16",x"4d2d15",x"4d2d17",x"513118",x"523219",x"543119",x"4f2f17",x"4f2f17",x"502f17",x"513018",x"533218",x"5a361b",x"543218",x"4b2a13",x"4a2913",x"563217",x"522e15",x"502d15",x"512e15",x"4c2a13",x"4c2a13",x"502e15",x"522f17",x"4d2b14",x"4a2912",x"4d2c14",x"553118",x"4e2d15",x"492a13",x"502d15",x"492913",x"4f2d16",x"523118",x"4f3017",x"513018",x"533219",x"543219",x"553319",x"533118",x"523017",x"4b2a14",x"4e2c15",x"543118",x"543218",x"543118",x"522f17",x"543117",x"512d15",x"533016",x"512d16",x"492812",x"4c2a13",x"502d15",x"512e16",x"4e2c14",x"502e15",x"4a2913",x"502e16",x"523118",x"553218",x"4e2d16",x"4f2f17",x"512f19",x"4f2d18",x"53311a",x"503019",x"53321b",x"52321c",x"4e2f1b",x"4a2c19",x"4b2c1a",x"4a2d1b",x"51321e",x"50301c",x"50301c",x"4c2e1b",x"4d2f1c",x"4a2e1b",x"4d2f1c",x"54321d",x"50311d",x"50311e",x"4e301b",x"4d2f1d",x"4d2f1c",x"4e311d",x"53331e",x"55361e",x"54331d",x"58361e",x"57361e",x"51311b",x"4f301b",x"54321c",x"4e2f1a",x"52311b",x"4e2f1a",x"4b2b17",x"4b2c16",x"4b2c16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1b1108",x"1d1208",x"1e1208",x"1d1108",x"1f1208",x"1f1209",x"201309",x"201309",x"211409",x"211409",x"201309",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1309",x"1f1208",x"201309",x"1f1309",x"201309",x"201309",x"1f1309",x"1f1208",x"1e1208",x"1e1208",x"1f1209",x"1f1309",x"1f1309",x"1f1309",x"1f1309",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"190f08",x"180f08",x"180f08",x"170f07",x"160f07",x"160e07",x"18110a",x"18110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1c1108",x"1d1208",x"1d1108",x"1d1108",x"1f1209",x"201309",x"201309",x"1f1209",x"1f1309",x"201309",x"201309",x"211409",x"201409",x"201409",x"211409",x"21150a",x"21150a",x"211409",x"201409",x"201309",x"201309",x"211409",x"201409",x"201309",x"1e1209",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1b1108",x"1c1108",x"1b1008",x"1b1108",x"1b1108",x"1a1008",x"191008",x"180f08",x"1a1008",x"1b1108",x"1c1108",x"1d1208",x"1f140a",x"1e130a",x"1b1108",x"1a1008",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"24150a",x"311c0d",x"211309",x"4a2b15",x"311c0d",x"422611",x"331d0d",x"412511",x"331d0d",x"150e07",x"492a13",x"150e07",x"150e07",x"2d1a0c",x"38210f",x"38200f",x"3d2411",x"38200f",x"3e2310",x"39200f",x"372110",x"27180b",x"26160a",x"543017",x"150e07",x"150e07",x"412511",x"432713",x"29180b",x"25160a",x"150e07",x"2d1a0c",x"341e0e",x"36200f",x"321d0e",x"2d1a0c",x"28170a",x"24150a",x"432611",x"2a180b",x"1b1108",x"37200f",x"422611",x"2e1b0c",x"150e07",x"150e07",x"1f1309",x"2a190b",x"2d1a0b",x"2c190b",x"2a180b",x"1e1108",x"2d190b",x"150e07",x"150e07",x"27160a",x"2b180b",x"311b0c",x"2d190b",x"2e190b",x"351e0e",x"361f0e",x"331d0d",x"311d0d",x"2d1a0c",x"2f1b0c",x"2d1a0c",x"422511",x"2d190b",x"2e1a0b",x"150e07",x"150e07",x"482812",x"24150a",x"472a14",x"502e16",x"4b2c15",x"4d2d16",x"432612",x"4c2c14",x"4d2c14",x"442611",x"522e16",x"4a2a13",x"4f2d16",x"4a2b14",x"4e2e16",x"533118",x"492b15",x"462914",x"472a14",x"4b2c15",x"4b2d17",x"4b2c15",x"442813",x"482a14",x"4c2c15",x"4f2f17",x"513118",x"59351a",x"4c2d16",x"543118",x"4f2e16",x"543016",x"502e15",x"533117",x"502f16",x"502d15",x"502e15",x"4a2913",x"412511",x"462812",x"482912",x"452812",x"452712",x"4c2c15",x"4e2e16",x"4f2f16",x"4b2c15",x"4e2e16",x"4b2c15",x"462812",x"523118",x"4c2e17",x"4f2f16",x"533016",x"502e16",x"4c2b15",x"4d2c15",x"522f17",x"533118",x"502f17",x"563319",x"5f371b",x"533118",x"663c1f",x"5b361b",x"533017",x"522f17",x"553017",x"533116",x"512f16",x"442712",x"4e2e16",x"4c2d16",x"4c2d16",x"583319",x"4d2e18",x"492a15",x"4b2d17",x"482b16",x"502f19",x"4d2b18",x"4a2c19",x"412716",x"58351d",x"50311d",x"4c2f1b",x"4b2d19",x"482c19",x"472b19",x"432919",x"472c1b",x"4f301d",x"4f301d",x"4f311e",x"482d1a",x"51331e",x"53341f",x"4e301d",x"482d1a",x"472b1a",x"492d1a",x"4c301c",x"472e1b",x"4f321d",x"4a2f1c",x"472c19",x"4e2f1c",x"52321c",x"4a2e1a",x"462b19",x"452a17",x"4b2c18",x"482a16",x"4a2c17",x"4a2c17",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1b1108",x"1c1108",x"1d1208",x"1e1209",x"1e1208",x"201309",x"201309",x"201309",x"1f1309",x"1f1209",x"1e1208",x"1f1208",x"221409",x"211409",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"201309",x"201309",x"201309",x"211409",x"211409",x"201409",x"201409",x"1f1208",x"1e1208",x"1e1208",x"1f1309",x"201309",x"1f1309",x"1f1309",x"1e1209",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"190f08",x"190f08",x"180f07",x"170f07",x"170f07",x"160f07",x"18110a",x"181109",x"1a130c",x"181009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f08",x"191008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1e1208",x"1f1309",x"1f1309",x"201309",x"211409",x"211409",x"211409",x"211409",x"201309",x"201309",x"22150a",x"21150a",x"201309",x"201309",x"211409",x"201309",x"201309",x"201409",x"201409",x"1f1309",x"1e1209",x"1d1209",x"1d1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1108",x"1a1008",x"191008",x"180f07",x"1a1008",x"1c1108",x"1c1108",x"1f130b",x"20150d",x"1e130b",x"1d1208",x"1d1108",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"190f08",x"190f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"25160a",x"311c0d",x"1f1208",x"462712",x"25150a",x"351d0d",x"301b0c",x"39200e",x"3d210e",x"3f220f",x"150e07",x"3b200e",x"2b180b",x"150e07",x"150e07",x"25150a",x"361e0d",x"351e0d",x"311c0c",x"341e0d",x"351f0f",x"37200f",x"2e1b0c",x"1e1209",x"2f1a0b",x"422511",x"150e07",x"25160a",x"3c220f",x"3f2411",x"150e07",x"150e07",x"24150a",x"24150a",x"26160a",x"201309",x"211409",x"371e0d",x"241509",x"150e07",x"180f07",x"201309",x"2a190b",x"371f0e",x"2d190b",x"150e07",x"150e07",x"1f1309",x"26160a",x"27170a",x"26160a",x"150e07",x"402410",x"39200e",x"150e07",x"1e1209",x"2b190b",x"2f1c0d",x"311c0d",x"311c0d",x"311c0d",x"2f1b0c",x"2c1a0c",x"2b190b",x"2b190b",x"28170b",x"25160a",x"4a2b14",x"2d190b",x"341d0c",x"150e07",x"150e07",x"241509",x"2c190b",x"231409",x"442813",x"311c0c",x"2d190b",x"351e0d",x"3b220f",x"4c2d15",x"543219",x"412612",x"4d2e16",x"502f17",x"4b2d16",x"402612",x"432713",x"3f2511",x"341e0e",x"3b2311",x"3e2411",x"422712",x"442814",x"3d2411",x"513118",x"3d2411",x"452612",x"3e220f",x"472712",x"3e2411",x"4a2b13",x"492912",x"4d2b14",x"4f2c14",x"402411",x"3d220f",x"412411",x"3e230f",x"412511",x"39200e",x"3b210e",x"331c0c",x"3f220f",x"341d0d",x"3c220e",x"3b210f",x"3c220f",x"4b2a13",x"4c2a14",x"522f15",x"412512",x"4c2e17",x"513118",x"4d2d16",x"5b371c",x"4e2e15",x"4b2a15",x"402412",x"412612",x"432714",x"4e2d17",x"4e2e16",x"4d2d16",x"523118",x"502e17",x"61391c",x"522f17",x"4a2b15",x"4d2c16",x"412411",x"412511",x"472a15",x"462914",x"503018",x"56341a",x"3e2313",x"533119",x"422615",x"472b18",x"53321a",x"57341d",x"53331b",x"4a2d1b",x"4a2d19",x"492d1b",x"4f301d",x"492e1c",x"482d1b",x"543420",x"4b301d",x"462d1c",x"452d1c",x"4a2f1d",x"4b301d",x"422b1c",x"402a1b",x"422a1a",x"422c1c",x"472e1c",x"482e1d",x"482f1d",x"462e1c",x"462d1c",x"462d1c",x"4c311e",x"472d1a",x"4f321e",x"3e2819",x"492d1a",x"3c2617",x"412918",x"432a18",x"4b2e1b",x"56341c",x"3e2515",x"3e2515",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1f1208",x"1f1208",x"1f1208",x"201208",x"1f1208",x"201308",x"211409",x"231409",x"24150a",x"25150a",x"241509",x"241509",x"25150a",x"231509",x"231509",x"24150a",x"241509",x"231509",x"221509",x"231409",x"221409",x"231509",x"231509",x"231409",x"24150a",x"231409",x"211409",x"221509",x"211309",x"1e1108",x"1f1309",x"1f1208",x"1e1208",x"1e1309",x"1e1208",x"1c1108",x"1c1108",x"1a1108",x"191008",x"191008",x"180f07",x"170f07",x"191109",x"1a130c",x"1a130c",x"1a130c",x"18100a",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"191008",x"1a1008",x"1c1108",x"1c1108",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1f1208",x"201309",x"211309",x"211409",x"211409",x"221409",x"231509",x"231409",x"221409",x"231409",x"231409",x"231509",x"231509",x"23150a",x"231509",x"221409",x"211409",x"201309",x"1f1208",x"201309",x"211409",x"211409",x"211309",x"201309",x"1f1208",x"1e1208",x"1e1208",x"1d1208",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"190f08",x"190f08",x"1a1008",x"1c1108",x"1d1108",x"1e1209",x"20140c",x"1f140b",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"190f07",x"180f07",x"381f0e",x"170f08",x"492812",x"4b2a13",x"472812",x"472812",x"4c2c15",x"492a13",x"492812",x"472711",x"462611",x"492812",x"462711",x"472812",x"502f16",x"533118",x"543319",x"57331a",x"533219",x"553319",x"4f2e16",x"543319",x"513018",x"4f2e16",x"4d2d16",x"4e2d15",x"4f2f17",x"4e2d16",x"4a2913",x"4b2a13",x"4c2c14",x"4a2a14",x"4d2c15",x"4d2c15",x"432511",x"432510",x"4a2a13",x"4e2d16",x"4c2c15",x"482a13",x"482812",x"442611",x"432511",x"482812",x"472812",x"432510",x"412410",x"3d220e",x"442712",x"4d2d16",x"4a2b14",x"492a14",x"442711",x"482913",x"4b2a14",x"4a2a13",x"482812",x"442611",x"452711",x"472811",x"4a2b12",x"492a12",x"3b1f0b",x"42240f",x"492a11",x"472811",x"472811",x"482a12",x"482a12",x"472912",x"482912",x"452711",x"472811",x"472812",x"482912",x"452711",x"442610",x"42240f",x"432510",x"472812",x"4a2b13",x"4b2b14",x"4d2d15",x"4c2c15",x"4e2d16",x"4e2d16",x"472914",x"4b2b15",x"4a2c15",x"4c2c15",x"4e2e16",x"513016",x"4c2d14",x"4f2f14",x"4f2e14",x"4b2b13",x"502f14",x"492b13",x"4c2c13",x"502e15",x"543216",x"523015",x"492b11",x"4c2b12",x"492812",x"512d15",x"3f2411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"201309",x"37200f",x"211409",x"492812",x"3e230f",x"3e220f",x"3e220f",x"3c210e",x"3a200e",x"3b200e",x"432511",x"452712",x"150e07",x"2d1a0c",x"412511",x"2e1b0c",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"381f0e",x"150e07",x"311c0c",x"3d220f",x"241509",x"150e07",x"150e07",x"170f07",x"2a180b",x"412611",x"150e07",x"150e07",x"24150a",x"2f1b0d",x"2f1b0d",x"29180b",x"25160a",x"2b190b",x"351e0d",x"231509",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2411",x"150e07",x"2e1b0d",x"472914",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"462913",x"2a180a",x"311b0b",x"39200c",x"39200c",x"39200c",x"231409",x"1f140b",x"201309",x"3a2210",x"3d2411",x"452913",x"452813",x"4c2d15",x"4d2d15",x"502f16",x"4c2d16",x"523118",x"492a15",x"5a351a",x"4b2b16",x"4e2e17",x"462813",x"4a2d16",x"4c2e16",x"4b2c16",x"58351a",x"492b15",x"513017",x"4e2c14",x"4b2b15",x"502f16",x"4f2e16",x"42230f",x"3f200d",x"46260f",x"522f16",x"512f15",x"4b2a13",x"4a2912",x"3f2310",x"452610",x"482812",x"3e220f",x"452611",x"482812",x"4d2c14",x"482913",x"452712",x"4a2a14",x"482913",x"553116",x"522f16",x"523118",x"432511",x"512d15",x"583318",x"5d361b",x"60381c",x"5b351a",x"512e15",x"4b2a13",x"543016",x"4c2b14",x"512d15",x"553016",x"472812",x"3e1f0d",x"4c2a12",x"4e2b13",x"4f2c14",x"512e15",x"4f2d16",x"4b2c16",x"4b2c16",x"533218",x"513018",x"4d2e17",x"523119",x"503019",x"55311a",x"563219",x"502e19",x"54321b",x"57341d",x"5c371e",x"5f3b21",x"56351f",x"553620",x"5f3b23",x"5b3821",x"50331e",x"543520",x"533520",x"4f321f",x"50321e",x"4b301d",x"492e1c",x"492f1d",x"482e1c",x"4a2f1d",x"553620",x"50321f",x"51341f",x"533520",x"50331f",x"4e331f",x"4e2f1b",x"53321e",x"54351f",x"5e3b23",x"54341d",x"52331d",x"57361e",x"4e301c",x"4c2f1b",x"4e2f1b",x"4d2f1b",x"4d2e18",x"4d2e18",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"1d1208",x"231509",x"2c190b",x"331d0d",x"37200f",x"361f0f",x"351d0e",x"361f0e",x"351f0e",x"341d0d",x"351f0e",x"37200f",x"351f0e",x"331e0e",x"341e0e",x"361f0e",x"361f0e",x"351e0e",x"331c0c",x"321c0c",x"341d0d",x"351e0d",x"351e0d",x"341d0d",x"351e0d",x"341d0d",x"331c0d",x"311b0b",x"321c0d",x"351e0d",x"37200e",x"3a210f",x"3c2210",x"3c2310",x"3d2310",x"3d2310",x"3e2311",x"3b220f",x"3a210f",x"39210f",x"38200f",x"351f0e",x"311c0d",x"2f1c0d",x"2f1b0d",x"2d1b0c",x"29180b",x"221409",x"1d1208",x"1f1208",x"211309",x"211309",x"1f1309",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"211309",x"241509",x"29170b",x"2a180b",x"2d190b",x"2b180a",x"2d190b",x"2f1a0b",x"2f1b0c",x"301b0c",x"2e190b",x"2f1a0b",x"2a170a",x"261509",x"2d1a0a",x"291709",x"271609",x"261509",x"251409",x"251409",x"271509",x"28160a",x"261509",x"261409",x"261509",x"271609",x"28160a",x"27160a",x"231409",x"1e1208",x"180f07",x"150e07",x"150e07",x"160f07",x"180f07",x"211309",x"201309",x"1f1208",x"1e1208",x"1e1208",x"1d1208",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"190f08",x"190f08",x"1a1008",x"1c1108",x"1d1108",x"1e1209",x"20140c",x"1f140b",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"5e493a",x"5e493a",x"4e2d14",x"4c2b14",x"4d2b14",x"4b2b14",x"4c2b14",x"4c2a13",x"502d15",x"4e2d16",x"4c2a14",x"4a2913",x"492912",x"492812",x"4b2a13",x"472812",x"472812",x"4c2c15",x"492a13",x"492812",x"472711",x"462611",x"492812",x"462711",x"472812",x"502f16",x"533118",x"543319",x"57331a",x"533219",x"553319",x"4f2e16",x"543319",x"513018",x"4f2e16",x"4d2d16",x"4e2d15",x"4f2f17",x"4e2d16",x"4a2913",x"4b2a13",x"4c2c14",x"4a2a14",x"4d2c15",x"4d2c15",x"432511",x"432510",x"4a2a13",x"4e2d16",x"4c2c15",x"482a13",x"482812",x"442611",x"432511",x"482812",x"472812",x"432510",x"412410",x"3d220e",x"442712",x"4d2d16",x"4a2b14",x"492a14",x"442711",x"482913",x"4b2a14",x"4a2a13",x"482812",x"442611",x"452711",x"472811",x"4a2b12",x"492a12",x"3b1f0b",x"42240f",x"492a11",x"472811",x"472811",x"482a12",x"482a12",x"472912",x"482912",x"452711",x"472811",x"472812",x"482912",x"452711",x"442610",x"42240f",x"432510",x"472812",x"4a2b13",x"4b2b14",x"4d2d15",x"4c2c15",x"4e2d16",x"4e2d16",x"472914",x"4b2b15",x"4a2c15",x"4c2c15",x"4e2e16",x"513016",x"4c2d14",x"4f2f14",x"4f2e14",x"4b2b13",x"502f14",x"492b13",x"4c2c13",x"502e15",x"543216",x"523015",x"492b11",x"4c2b12",x"492812",x"512d15",x"3f2411",x"3f2411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"211409",x"361f0e",x"3b210f",x"3b220f",x"3b2210",x"311c0d",x"492912",x"2a180b",x"301b0c",x"40230f",x"311b0b",x"331c0c",x"381f0d",x"422510",x"452611",x"41230f",x"472711",x"3f220e",x"442510",x"482711",x"4c2a13",x"4a2912",x"442611",x"492912",x"4a2a13",x"512e15",x"4d2c14",x"452712",x"412410",x"422410",x"452711",x"3e220f",x"3c200d",x"40230f",x"361e0d",x"371f0e",x"331c0c",x"381e0d",x"301b0b",x"29170a",x"2a170a",x"462711",x"351e0d",x"2f1a0b",x"3d210e",x"361e0d",x"2c190b",x"2d190b",x"3c210f",x"40240f",x"432510",x"361d0c",x"391f0d",x"3a200e",x"3a200e",x"422410",x"462711",x"4e2b14",x"4c2b13",x"4c2b14",x"452812",x"4e2c14",x"4b2c15",x"4b2b15",x"513018",x"4a2c16",x"4c2d15",x"452813",x"281709",x"2f1a0b",x"3b200d",x"3b200d",x"3b200d",x"000000",x"201309",x"2d180a",x"2b170a",x"492c15",x"492c15",x"502f17",x"4e2e17",x"573319",x"472812",x"4e2c14",x"492a14",x"4e2d16",x"523118",x"523119",x"4f3017",x"56331a",x"523118",x"4f2f17",x"523119",x"422511",x"4c2c15",x"4d2d16",x"4c2c13",x"4e2d15",x"512f17",x"5c371b",x"573217",x"4a2912",x"4e2c14",x"4f2c14",x"4a2913",x"593318",x"4c2b14",x"553218",x"4e2c14",x"4c2b13",x"4a2913",x"4c2a13",x"482711",x"452711",x"452510",x"4a2912",x"512c14",x"462610",x"4a2a12",x"452610",x"40210e",x"482712",x"4b2912",x"4e2c14",x"4e2b13",x"4f2c14",x"532f16",x"522e15",x"502d15",x"522f16",x"532f15",x"4c2a14",x"4b2912",x"4b2a13",x"472610",x"4c2a13",x"492912",x"4d2b14",x"4e2c14",x"492812",x"452610",x"462711",x"472912",x"482813",x"472914",x"4c2c16",x"472916",x"492a16",x"4c2d18",x"482a16",x"4e2d19",x"502f1b",x"4d2e1a",x"4d2e19",x"472b1a",x"472b18",x"52311d",x"4d2f1d",x"4d2f1c",x"482d1a",x"4c2f1d",x"4f311d",x"4e311e",x"4f301c",x"4f321e",x"4d321e",x"513320",x"523620",x"543620",x"573620",x"51321d",x"573721",x"563620",x"533420",x"5c3a23",x"52331e",x"563720",x"543520",x"593820",x"58371f",x"5c3a21",x"56351d",x"55361e",x"56351c",x"432917",x"4f3019",x"4f3019",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"1d1208",x"231509",x"2c190b",x"331d0d",x"37200f",x"361f0f",x"351d0e",x"361f0e",x"351f0e",x"341d0d",x"351f0e",x"37200f",x"351f0e",x"331e0e",x"341e0e",x"361f0e",x"361f0e",x"351e0e",x"331c0c",x"321c0c",x"341d0d",x"351e0d",x"351e0d",x"341d0d",x"351e0d",x"341d0d",x"331c0d",x"311b0b",x"321c0d",x"351e0d",x"37200e",x"3a210f",x"3c2210",x"3c2310",x"3d2310",x"3d2310",x"3e2311",x"3b220f",x"3a210f",x"39210f",x"38200f",x"351f0e",x"311c0d",x"2f1c0d",x"2f1b0d",x"2d1b0c",x"29180b",x"221409",x"1d1208",x"1f1208",x"211309",x"211309",x"1f1309",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"211309",x"241509",x"29170b",x"2a180b",x"2d190b",x"2b180a",x"2d190b",x"2f1a0b",x"2f1b0c",x"301b0c",x"2e190b",x"2f1a0b",x"2a170a",x"261509",x"2d1a0a",x"291709",x"271609",x"261509",x"251409",x"251409",x"271509",x"28160a",x"261509",x"261409",x"261509",x"271609",x"28160a",x"27160a",x"231409",x"1e1208",x"180f07",x"150e07",x"150e07",x"160f07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594638",x"594638",x"472814",x"482b15",x"4c2d16",x"452913",x"412612",x"422612",x"422612",x"432713",x"452813",x"432713",x"462914",x"432713",x"452813",x"422713",x"422713",x"462a14",x"452914",x"472a15",x"442813",x"3e2310",x"402410",x"3e2310",x"432712",x"472a14",x"422713",x"472a14",x"4b2d16",x"442814",x"432713",x"3f2612",x"3a200f",x"37200f",x"3a2310",x"3a210f",x"3d2310",x"402512",x"3f2512",x"3f2410",x"3a200e",x"3c210f",x"39200f",x"371f0d",x"3d230f",x"3c2210",x"402511",x"3d220f",x"3b210e",x"3b210f",x"39200e",x"361e0d",x"351d0c",x"351d0d",x"371e0d",x"371e0d",x"361e0d",x"3b200e",x"301b0c",x"341c0c",x"371e0d",x"361e0d",x"3b210f",x"311b0c",x"3b210f",x"3c220f",x"3c220f",x"3e2310",x"3f2310",x"3f240f",x"3e240f",x"3d240e",x"3a230d",x"39210d",x"3c220d",x"3e250e",x"3a210e",x"3d230f",x"3a220d",x"361f0c",x"381f0d",x"38200d",x"361f0d",x"351e0c",x"3c230e",x"3b220d",x"3c230d",x"331e0c",x"341d0c",x"321d0b",x"361e0d",x"361e0c",x"341d0c",x"331d0c",x"341c0c",x"331d0c",x"361e0d",x"311c0c",x"351e0d",x"341e0d",x"38200e",x"39200e",x"3e240f",x"39220e",x"3e2510",x"402712",x"3e2510",x"3c2410",x"3d2410",x"3c2410",x"422711",x"482c12",x"442811",x"432811",x"422811",x"39220f",x"462914",x"361f0f",x"361f0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"241509",x"351e0e",x"351d0d",x"231409",x"351c0c",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"341c0b",x"150e07",x"371c0c",x"150e07",x"150e07",x"1b1108",x"211309",x"1c1108",x"211308",x"221308",x"201208",x"211308",x"241509",x"221409",x"1e1208",x"27170b",x"231509",x"25150a",x"25150a",x"231409",x"170f07",x"150e07",x"150e07",x"150e07",x"311c0c",x"180f08",x"150e07",x"150e07",x"331e0e",x"492c15",x"150e07",x"150e07",x"150e07",x"191008",x"170f07",x"27160a",x"422511",x"201309",x"1c1108",x"150e07",x"150e07",x"2d1a0c",x"341e0e",x"37200f",x"3b2311",x"351f0f",x"39200f",x"361f0e",x"301c0c",x"311b0c",x"29170a",x"2f1b0c",x"2f1b0c",x"2b190b",x"2f1b0c",x"27160a",x"2c190b",x"3c210f",x"2b180a",x"2d190b",x"381f0c",x"3a200d",x"3a200d",x"000000",x"000000",x"2b170a",x"3a2110",x"3d2511",x"502f17",x"543319",x"543218",x"5e381c",x"4e2d16",x"4f2f16",x"563318",x"4e2d15",x"4e2d15",x"502e16",x"4f2e16",x"4c2d15",x"502e15",x"482812",x"462710",x"3f230f",x"402410",x"4a2912",x"482812",x"4c2b14",x"4d2b14",x"462711",x"452610",x"482811",x"462711",x"4b2a12",x"432510",x"472610",x"3f220e",x"40230e",x"3d220e",x"462610",x"43230f",x"3f220e",x"41230e",x"41230e",x"41220e",x"3c1f0d",x"3f230e",x"43240f",x"41230f",x"432410",x"43240f",x"44240f",x"45250f",x"46260f",x"482711",x"553116",x"543117",x"543117",x"553117",x"563117",x"522e15",x"532e16",x"502d15",x"4d2a14",x"512d15",x"4f2b14",x"4c2913",x"492912",x"4f2b14",x"593419",x"57341a",x"5b381c",x"5d391d",x"5a361c",x"5a361c",x"56351c",x"57331b",x"4f2e18",x"4e2d18",x"59351d",x"5c3920",x"5a3920",x"5e3b21",x"5d3a21",x"553520",x"5b3a22",x"5c3b23",x"613d24",x"593620",x"55351f",x"57361f",x"513420",x"4d311f",x"4a2f1d",x"4a2f1d",x"492f1d",x"4e311e",x"4c301e",x"462c1c",x"51321f",x"533420",x"53331f",x"56351e",x"5a371f",x"553420",x"54341f",x"5c3922",x"56361f",x"523520",x"52331d",x"50321d",x"53351e",x"5b391f",x"51331d",x"5a381e",x"442b17",x"442b17",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"201309",x"2b190c",x"331e0e",x"39210f",x"3b2311",x"38200f",x"341d0d",x"321c0c",x"351d0d",x"39210f",x"392210",x"38210f",x"38200f",x"37200f",x"38210f",x"3c2311",x"3d2512",x"3a2210",x"38200f",x"38200f",x"37200e",x"361e0e",x"361e0e",x"361e0e",x"361e0e",x"371f0e",x"361e0e",x"331c0c",x"321c0c",x"341d0d",x"381f0e",x"3b220f",x"3c220f",x"3d2310",x"3e2310",x"3f2411",x"412612",x"402512",x"3f2511",x"3d2411",x"3b2210",x"392210",x"36200f",x"321e0e",x"301c0d",x"2d1b0c",x"28180b",x"221409",x"1f1309",x"211409",x"24150a",x"23150a",x"201309",x"1d1208",x"1c1108",x"1b1108",x"1c1108",x"1d1108",x"221409",x"27160a",x"28170a",x"29170a",x"2b180a",x"2d190b",x"2f1a0b",x"2e1a0b",x"2e1a0b",x"2b170a",x"2c180a",x"2c180a",x"2a170a",x"29170a",x"2f1b0a",x"2b1809",x"281609",x"271509",x"271509",x"271509",x"271609",x"28160a",x"29170a",x"28160a",x"271609",x"261509",x"261509",x"261509",x"241409",x"201309",x"191008",x"150e07",x"150e07",x"160f07",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5f4b3e",x"5f4b3e",x"3b210f",x"39200f",x"331d0c",x"341c0d",x"341d0d",x"361f0e",x"3b220f",x"3c220f",x"371f0e",x"39200f",x"38200f",x"392110",x"3a2210",x"37200f",x"3d2411",x"3b2210",x"3e2411",x"3e2511",x"3b2310",x"3f2411",x"3a2310",x"38210f",x"3a210f",x"38200e",x"38200f",x"37200f",x"331d0d",x"381f0e",x"321c0c",x"301b0c",x"2f1a0b",x"26160a",x"311b0c",x"2e1a0b",x"321c0c",x"341d0d",x"2e1a0b",x"2d190b",x"301b0c",x"301a0b",x"251509",x"2f1a0b",x"2e1a0b",x"2d180a",x"28160a",x"2b180a",x"2a170a",x"29170a",x"2a170a",x"2a170a",x"29160a",x"281509",x"281509",x"261509",x"251509",x"2e190b",x"150e07",x"8b7156",x"7f674f",x"897355",x"8f785b",x"8c7157",x"8a7056",x"957a5d",x"8d7558",x"876e54",x"65523e",x"39210d",x"37210d",x"301c0b",x"351f0c",x"321d0c",x"36200c",x"3a220d",x"38210c",x"341d0c",x"3b220e",x"3e2610",x"3a230f",x"3e260f",x"3a230e",x"3d240f",x"412710",x"41270f",x"3c230e",x"331e0b",x"39210e",x"3a210f",x"331e0d",x"341f0e",x"331e0e",x"36200e",x"341f0e",x"341f0f",x"37200e",x"37210e",x"35200d",x"38220e",x"331f0d",x"2d1a0b",x"341f0d",x"39220d",x"37200c",x"36200c",x"321d0b",x"341e0c",x"38210d",x"37210d",x"3d240e",x"3d250e",x"36210c",x"36200c",x"39220e",x"351f0d",x"3f2511",x"201309",x"201309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"241509",x"341e0e",x"321c0c",x"3f220e",x"150e07",x"1c1108",x"261409",x"2a170a",x"2b170a",x"2b180a",x"1f1208",x"3f230f",x"150e07",x"191008",x"2d190b",x"2e190b",x"311c0c",x"321c0c",x"381f0e",x"39200e",x"38200e",x"361e0d",x"341d0c",x"351d0d",x"38200e",x"39210f",x"3b2310",x"3b2210",x"351e0d",x"351d0d",x"301b0c",x"341d0d",x"321d0d",x"2f1b0d",x"191008",x"1f1309",x"3b2210",x"2f1c0d",x"492a14",x"150e07",x"150e07",x"25160a",x"311d0d",x"351f0f",x"321d0e",x"2b190b",x"39210f",x"4f2d15",x"150e07",x"25160a",x"27170b",x"36200f",x"382110",x"3c2411",x"3b2311",x"3c2311",x"3a2210",x"37200f",x"351f0e",x"37200f",x"351f0e",x"331d0e",x"392110",x"351f0f",x"2f1b0c",x"311d0d",x"341f0e",x"4b2c15",x"301b0b",x"321c0b",x"361d0b",x"361d0b",x"361d0b",x"000000",x"000000",x"000000",x"3f2612",x"412712",x"3f2512",x"58351a",x"56341a",x"59361b",x"56341a",x"543119",x"4f2e16",x"58351a",x"57341a",x"59351a",x"58351a",x"563419",x"533117",x"4c2c15",x"4d2d15",x"4e2d16",x"4c2c15",x"422410",x"3b200e",x"472711",x"492912",x"482812",x"4d2c14",x"4c2b14",x"4a2a13",x"492812",x"482711",x"43230f",x"3f220e",x"3c200d",x"391e0c",x"3d1f0d",x"40220e",x"42230e",x"442510",x"462611",x"442510",x"472711",x"43250f",x"43240f",x"492912",x"4a2912",x"462711",x"4d2c14",x"4c2b14",x"4b2b13",x"482811",x"452610",x"4d2b14",x"4d2d14",x"523017",x"512f17",x"4d2c15",x"4a2a13",x"492812",x"4d2b14",x"512f16",x"523017",x"523017",x"513017",x"502f17",x"522f16",x"513017",x"503017",x"513017",x"523119",x"4b2d18",x"503019",x"54331c",x"57341d",x"4e2f1c",x"4b2e1b",x"52321c",x"54341f",x"57361f",x"52331e",x"553620",x"583720",x"583822",x"593821",x"593921",x"5c3a23",x"563620",x"533520",x"533521",x"523420",x"50341f",x"4d311f",x"4f321f",x"503320",x"5a3921",x"563721",x"563621",x"553620",x"53341e",x"55351e",x"52341f",x"57361f",x"53341e",x"53331e",x"4f321d",x"56351e",x"573620",x"58371f",x"58371f",x"58371f",x"57361e",x"52321c",x"52321c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"191008",x"211409",x"2b190b",x"321d0d",x"39210f",x"3a2110",x"3b2210",x"3c2310",x"3b2310",x"3b220f",x"39200f",x"3b2210",x"3c2310",x"37200f",x"37200f",x"3b2311",x"3b2310",x"3d2311",x"3e2411",x"3d2411",x"3b2210",x"3a220f",x"3b2210",x"3c2310",x"3c2310",x"3c2310",x"3c2311",x"371f0e",x"3e2511",x"3e2411",x"3c2310",x"3f2512",x"422712",x"422712",x"432813",x"452914",x"452914",x"422712",x"402511",x"3e2411",x"3e2411",x"3e2411",x"3d2411",x"392210",x"36200f",x"341f0f",x"2e1b0c",x"2a190b",x"27170b",x"24160a",x"27170b",x"2a190c",x"29180b",x"26170b",x"221509",x"221409",x"211409",x"201309",x"1f1208",x"221409",x"27160a",x"2b190b",x"2d190b",x"321d0d",x"341d0d",x"341d0d",x"331c0c",x"311b0c",x"2f1a0b",x"2e190b",x"2c180a",x"291609",x"29160a",x"2d190a",x"2c190a",x"2c180a",x"2b180a",x"2b180a",x"2b180a",x"2c180a",x"2a170a",x"2e1a0b",x"2e1a0b",x"2e1b0b",x"2f1b0c",x"301c0c",x"2d190b",x"27160a",x"201308",x"1a1008",x"160e07",x"150e07",x"170f07",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574132",x"574132",x"3f2411",x"3c220f",x"3d2311",x"3e2511",x"3e2411",x"3d2411",x"37200f",x"3e2411",x"3a2110",x"3d2411",x"3d2411",x"3d2411",x"3a2110",x"361f0e",x"3b2210",x"3c2311",x"3b2310",x"3c2311",x"3b2311",x"422713",x"3d2411",x"361f0e",x"3e2511",x"382210",x"3b2311",x"3d2512",x"3b2311",x"3b2310",x"361e0e",x"38200f",x"2c1a0c",x"331d0e",x"311c0c",x"301b0b",x"2c180b",x"29180a",x"331c0d",x"321d0d",x"341d0d",x"361f0e",x"2e1a0b",x"311b0b",x"2e190b",x"2e190b",x"2d190a",x"2c170a",x"2c170a",x"291609",x"2a170a",x"2a170a",x"29170a",x"211309",x"2c180b",x"29170a",x"2c180a",x"29170a",x"967d5e",x"967d5f",x"987d61",x"957c5d",x"93795c",x"826c50",x"987b60",x"987d60",x"967d5f",x"947a5d",x"876d51",x"37200e",x"311c0b",x"331d0c",x"331e0b",x"35200c",x"37210d",x"3f2610",x"38220e",x"39220e",x"3b220e",x"3f260f",x"40260f",x"3d240f",x"39220e",x"3c240f",x"412710",x"412811",x"432910",x"3b240e",x"3a230e",x"38220d",x"39220f",x"3c2410",x"351f0d",x"39210e",x"3c2410",x"39220e",x"36200e",x"3d2510",x"351f0e",x"38210e",x"37210e",x"331e0d",x"2f1c0c",x"321e0d",x"37220d",x"38210d",x"341f0c",x"39230f",x"37220e",x"36200d",x"3e260f",x"432811",x"36210d",x"3d240f",x"35200e",x"36200e",x"3d2311",x"26170a",x"26170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"231409",x"38200f",x"3a200d",x"150e07",x"150e07",x"241409",x"2a170a",x"2a1609",x"2a1609",x"2c180a",x"28160a",x"150e07",x"150e07",x"29170a",x"321c0c",x"351e0d",x"351e0d",x"371f0e",x"351e0d",x"311b0b",x"301a0b",x"311b0c",x"3a200e",x"381f0e",x"391f0d",x"361d0c",x"381f0d",x"3d230f",x"341e0c",x"3e2410",x"3d230f",x"331e0c",x"38200d",x"39210e",x"38200d",x"2f1c0b",x"1c1208",x"482a14",x"1b1108",x"1d1308",x"2a180b",x"2a190b",x"301c0d",x"3c2311",x"37200f",x"321d0e",x"3c2311",x"150e07",x"150e07",x"2b190b",x"2e1b0c",x"3d2411",x"3b2311",x"3b2310",x"3b2411",x"3d2411",x"402612",x"371f0f",x"351f0e",x"3e2411",x"331e0e",x"37200f",x"371f0e",x"2d1a0b",x"28170a",x"2e1a0c",x"341e0e",x"4a2b14",x"331c0c",x"29170a",x"3b200d",x"3a1f0d",x"3a1f0d",x"000000",x"000000",x"000000",x"000000",x"4a2a14",x"472812",x"57341a",x"553219",x"502f17",x"543018",x"523117",x"533118",x"522f17",x"533118",x"513017",x"5a361a",x"59361b",x"533118",x"512f17",x"533117",x"502f16",x"4d2b14",x"4e2d15",x"4d2c15",x"4f2e16",x"512f16",x"543118",x"4a2912",x"482711",x"492711",x"462611",x"472610",x"452510",x"43240f",x"43230e",x"41230e",x"42230e",x"3d200d",x"41210e",x"452610",x"472711",x"4d2b13",x"472812",x"4e2c14",x"4c2a13",x"4d2b13",x"512d15",x"502d15",x"482811",x"41230e",x"46250f",x"472711",x"4d2b13",x"492812",x"452510",x"432510",x"4f2c14",x"512e16",x"553117",x"543117",x"512f16",x"502d15",x"533016",x"563117",x"522f16",x"543017",x"563218",x"58351a",x"553218",x"56341b",x"58331b",x"513019",x"5a361d",x"5f3c20",x"603c21",x"5a371f",x"5b3920",x"59361e",x"593720",x"5d3a22",x"5f3c22",x"5f3c23",x"5c3922",x"5e3b23",x"633f24",x"643f24",x"5e3c24",x"543521",x"5a3923",x"583821",x"5a3822",x"533420",x"4b301d",x"4e321f",x"4f321f",x"533521",x"53341f",x"53351f",x"54321d",x"52321d",x"4f311d",x"53341f",x"51321e",x"53321d",x"472c1b",x"55341e",x"5a3920",x"5a3920",x"5c3a21",x"57351e",x"59371e",x"53321b",x"3b2515",x"3b2515",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f08",x"1b1108",x"25150a",x"2f1b0d",x"3a2210",x"3d2310",x"3f2411",x"432813",x"452814",x"452914",x"462a14",x"3f2411",x"402511",x"402512",x"422713",x"422713",x"3f2511",x"422713",x"432814",x"412612",x"402612",x"3b210f",x"3e2411",x"3f2411",x"3e2411",x"3e2411",x"3b220f",x"3a210f",x"3a200e",x"3c2310",x"3d2311",x"3e2411",x"3d2310",x"3f2310",x"3f2310",x"402410",x"402410",x"402410",x"3f2310",x"402411",x"442813",x"442914",x"432813",x"3f2512",x"3c2311",x"351f0e",x"331d0e",x"321d0d",x"2d1b0c",x"29180b",x"27170b",x"2c1a0c",x"311d0e",x"311d0e",x"2d1b0c",x"29180b",x"28180b",x"26160a",x"25150a",x"28180b",x"2c190b",x"301c0d",x"341e0e",x"361f0e",x"341d0d",x"341d0d",x"351d0d",x"341d0c",x"331c0c",x"341c0c",x"321b0b",x"301a0b",x"2f190b",x"2d170a",x"301b0a",x"2d190a",x"2f1a0b",x"2f1a0b",x"321c0c",x"311c0c",x"321c0c",x"311c0c",x"321c0c",x"341d0d",x"331c0d",x"2f1a0b",x"2b170a",x"2c180a",x"2a180b",x"241509",x"1b1008",x"160e07",x"150e07",x"160e07",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c4434",x"5c4434",x"3b210f",x"331c0d",x"3a210f",x"3a2210",x"3e2411",x"3d2310",x"3a210f",x"351e0d",x"331d0d",x"3b210f",x"331d0d",x"371f0e",x"341d0d",x"321d0d",x"331e0e",x"402612",x"3b2310",x"3e2511",x"3c2311",x"38210f",x"3a2210",x"3c2310",x"392110",x"3a2110",x"39210f",x"37200f",x"3c2411",x"37200f",x"341e0e",x"39210f",x"321d0d",x"311c0c",x"361f0e",x"361f0f",x"2f1b0c",x"321d0d",x"39210f",x"321c0c",x"311c0c",x"311b0c",x"2f1a0b",x"2e190b",x"2d190b",x"331c0c",x"2e190a",x"2b170a",x"2a170a",x"2a1609",x"271509",x"29170a",x"2d190b",x"2e1a0b",x"301b0c",x"2f1b0c",x"321c0c",x"2c190b",x"987c60",x"977e60",x"987d5f",x"836d53",x"92795c",x"af9274",x"977b60",x"987c60",x"957c5d",x"917a5d",x"897257",x"361f0d",x"3d240f",x"3b230e",x"3d240e",x"351f0c",x"3a230d",x"3d240f",x"37210c",x"38200d",x"38220d",x"3e2610",x"321e0b",x"3b240e",x"3b240e",x"3c250e",x"3b240f",x"422910",x"3c250f",x"3f2710",x"402710",x"35200c",x"38210e",x"3a230f",x"3c2410",x"3d2511",x"3b230f",x"3a220f",x"38220f",x"38220f",x"3d250f",x"331e0c",x"321d0d",x"301c0c",x"351f0d",x"331f0c",x"37200d",x"35200c",x"321e0b",x"3c240e",x"2f1d0b",x"37210e",x"3a220d",x"3a220d",x"37200d",x"331e0b",x"321e0c",x"2f1c0b",x"39200e",x"231509",x"231509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"2a190b",x"402512",x"351c0c",x"281609",x"150e07",x"1f1208",x"251509",x"2a170a",x"331d0c",x"2f1b0b",x"2d1a0b",x"4a2912",x"150e07",x"1d1108",x"341e0d",x"331c0d",x"311b0b",x"361e0d",x"38200e",x"3b2210",x"371f0e",x"381f0e",x"361e0d",x"38200e",x"3b2210",x"3a210f",x"3f2410",x"3b2210",x"361f0e",x"39210f",x"38200e",x"38200e",x"39200d",x"331d0d",x"361f0d",x"321d0c",x"301c0b",x"201409",x"4d2d15",x"1c1208",x"191007",x"26160a",x"2f1b0c",x"2e1b0c",x"2f1b0c",x"1d1208",x"422713",x"523018",x"150e07",x"1c1108",x"2d1b0d",x"36200f",x"301c0d",x"361f0f",x"392210",x"37200f",x"341e0e",x"36200f",x"36200f",x"361f0e",x"331d0d",x"351e0e",x"2d1a0c",x"2f1b0d",x"36200f",x"3b2310",x"361f0e",x"4b2b15",x"2d190a",x"2e1a0a",x"462710",x"462710",x"462710",x"000000",x"000000",x"000000",x"4f301c",x"482c19",x"311f14",x"513727",x"513727",x"513623",x"503827",x"553824",x"4f3422",x"4d3423",x"4b372a",x"433124",x"483224",x"493425",x"4b3222",x"463021",x"432d1e",x"3f2b1e",x"3d2d22",x"422f24",x"473326",x"473123",x"493325",x"4b3324",x"462e20",x"463022",x"453023",x"39291d",x"403025",x"452f21",x"483123",x"4b3426",x"483021",x"493020",x"482e1e",x"4b301f",x"4c3322",x"4a3120",x"4d3220",x"4e3322",x"503423",x"4d3322",x"4e3422",x"4d3423",x"4b3221",x"493222",x"493121",x"493121",x"482f20",x"452d1e",x"483020",x"4c3323",x"4b3223",x"493325",x"513927",x"4f3624",x"4b3221",x"4d3322",x"503524",x"4d3524",x"503726",x"4c3527",x"4f3828",x"553b2b",x"4f3626",x"513829",x"543b2a",x"4f3320",x"523724",x"543928",x"4d3627",x"513725",x"4e3627",x"573b29",x"583d2b",x"583c28",x"563a28",x"503827",x"513726",x"4d3626",x"4e3827",x"423328",x"4c3729",x"523828",x"4d3628",x"4b3525",x"503727",x"503827",x"4e3727",x"4e3929",x"4e392b",x"50392a",x"4c3626",x"513827",x"543a28",x"4e3627",x"4d3626",x"4d382a",x"46362a",x"433429",x"4b382b",x"4e3a2c",x"4e3727",x"4c3424",x"4f3727",x"4c3627",x"543e2f",x"523e30",x"504034",x"3d2a1c",x"3d2a1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"1a1008",x"1d1208",x"29180b",x"321c0d",x"39200e",x"402411",x"442712",x"452813",x"422511",x"422511",x"472914",x"472914",x"482a15",x"462914",x"482a15",x"452914",x"422612",x"422713",x"442814",x"422712",x"3e2411",x"432813",x"412612",x"3c210f",x"3c210f",x"3f2411",x"412612",x"422712",x"422713",x"412511",x"3f2411",x"402511",x"442713",x"452813",x"482a14",x"4a2b15",x"4a2c15",x"472914",x"452713",x"442712",x"432611",x"452813",x"432713",x"432713",x"402612",x"3a2210",x"37200f",x"36200f",x"311d0d",x"2d1a0c",x"2e1b0c",x"331e0e",x"37200f",x"37200f",x"341f0e",x"2e1a0c",x"2d1a0b",x"29170a",x"2b190b",x"2d190b",x"301b0c",x"311b0c",x"341d0d",x"361e0d",x"321b0b",x"321b0b",x"321b0b",x"331c0b",x"341c0b",x"351c0c",x"341c0b",x"361d0c",x"321b0b",x"331c0c",x"3a210e",x"361f0d",x"361e0d",x"341d0d",x"351e0d",x"351d0d",x"351e0d",x"341d0d",x"311b0b",x"351d0d",x"39210f",x"3b220f",x"3a210f",x"351e0d",x"301b0c",x"28170a",x"1f1309",x"170f07",x"150e07",x"160f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b3c31",x"4b3c31",x"3d2411",x"402512",x"3e2511",x"3c2310",x"3f2511",x"39210f",x"3c2310",x"3b2210",x"392110",x"3e2511",x"3e2411",x"3a210f",x"37200f",x"361f0e",x"341e0d",x"3b2310",x"3f2411",x"3b2310",x"3f2512",x"3e2411",x"3f2511",x"3f2411",x"38200f",x"39210f",x"3c2311",x"3b2310",x"3a2210",x"3c2311",x"37200f",x"301b0c",x"331c0c",x"331d0d",x"2e1a0c",x"331c0d",x"301c0c",x"331d0d",x"301b0c",x"2f1a0b",x"2e190a",x"2c170a",x"2b170a",x"2b180a",x"2c180a",x"2e190a",x"2b180a",x"29170a",x"2c180a",x"2d190b",x"341d0d",x"341d0d",x"2e1a0c",x"321c0c",x"2f1b0c",x"301b0c",x"311c0c",x"29170a",x"957b5f",x"987c60",x"977d5f",x"876f54",x"8d7458",x"a98b6b",x"887256",x"91775b",x"8e7758",x"92785b",x"846d52",x"3d2410",x"3c230f",x"38210e",x"3d250f",x"321e0b",x"331e0c",x"36200c",x"37210d",x"3b230d",x"311d0d",x"341f0d",x"38220e",x"37200c",x"36200d",x"36200d",x"39230e",x"3c240e",x"39230d",x"37220d",x"38220e",x"331e0d",x"38220e",x"3a230e",x"3a230f",x"402710",x"38210f",x"39220e",x"3c2410",x"3b230f",x"37200e",x"3a2310",x"331e0d",x"271709",x"341e0c",x"321e0d",x"38210e",x"2d1c0b",x"3c240f",x"39220d",x"36210d",x"3a220e",x"3b230e",x"36200d",x"38210e",x"301d0c",x"341f0e",x"341e0d",x"3d2310",x"221409",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"28170a",x"351e0e",x"391f0e",x"251509",x"472711",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422510",x"150e07",x"4a2912",x"150e07",x"150e07",x"27160a",x"29170a",x"2b180a",x"2a170a",x"2e1a0b",x"321d0d",x"2d190b",x"331d0d",x"321d0d",x"341e0e",x"331d0d",x"2f1b0c",x"2d1a0b",x"2f1b0c",x"2c190b",x"2b180b",x"2a180b",x"27160a",x"2b180b",x"26160a",x"26160a",x"29180b",x"201309",x"150e07",x"442611",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"2f1c0d",x"422611",x"1d1108",x"150e07",x"150e07",x"150e07",x"1e1209",x"24150a",x"211409",x"26170b",x"1f1208",x"27170a",x"321d0e",x"29180b",x"29180b",x"2b190b",x"2b190b",x"1b1108",x"26160a",x"25150a",x"2a180b",x"27160a",x"4a2a13",x"301b0b",x"311b0b",x"361d0b",x"371e0b",x"371e0b",x"000000",x"000000",x"000000",x"58371f",x"58371f",x"4e2f1b",x"502f1a",x"4f301c",x"54321c",x"54331d",x"4d2f1a",x"53341c",x"53331e",x"52321d",x"55351e",x"54351e",x"57361f",x"54341d",x"51311c",x"50311b",x"4e2f1a",x"50311c",x"51321d",x"4f311c",x"4d2f1c",x"492c19",x"52331d",x"4a2d1a",x"50301c",x"492d1a",x"4b2c18",x"4b2d19",x"492b18",x"482b19",x"482b18",x"482b18",x"4b2e19",x"482b17",x"482a18",x"472b18",x"482b17",x"462917",x"492b17",x"482b17",x"422615",x"492b17",x"422716",x"432715",x"422715",x"4e2f1a",x"482b17",x"4a2b16",x"50301a",x"4d2e19",x"4c2d18",x"492b17",x"492c17",x"4a2c17",x"442814",x"432714",x"422613",x"442714",x"432713",x"462814",x"482a15",x"4f2f19",x"4e2f19",x"4c2e17",x"472916",x"4d2e18",x"513119",x"4c2e1a",x"4f301a",x"4e2f1a",x"52331d",x"4c2e1a",x"4c2f1b",x"4c2e1b",x"50321e",x"52331d",x"573720",x"54351f",x"4f3320",x"533520",x"51331d",x"482d1c",x"503220",x"4e321f",x"4f331f",x"50321e",x"4f321e",x"4b2f1c",x"4b301d",x"4a2f1c",x"472d1c",x"4a2f1d",x"4d301c",x"472d1c",x"4c2f1c",x"492d1a",x"452919",x"462c19",x"4b2f1c",x"50321e",x"4e2f1b",x"4c2e1b",x"482b17",x"4a2c18",x"492c18",x"472915",x"452916",x"4d2d18",x"432714",x"432714",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"17100a",x"17100a",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"1b1108",x"1f1309",x"28170a",x"341e0d",x"3d2311",x"412511",x"472a14",x"472a14",x"492b15",x"452813",x"442712",x"432612",x"442711",x"452813",x"452814",x"452813",x"432713",x"412612",x"442813",x"331b0b",x"3e2411",x"3f2511",x"3e2411",x"3e2410",x"3f2411",x"3f2411",x"3d2310",x"3c220f",x"3c210f",x"3d2310",x"3c2310",x"3e2310",x"3e230f",x"3d210e",x"3b200e",x"402310",x"452812",x"472914",x"482a14",x"462813",x"412411",x"412511",x"402411",x"3b210f",x"39200e",x"361f0e",x"341d0d",x"331d0d",x"311c0d",x"2f1b0d",x"311c0d",x"361f0e",x"392110",x"3a2210",x"37200e",x"341e0d",x"321d0d",x"311c0c",x"321d0d",x"341e0d",x"351e0e",x"361e0d",x"39200f",x"3f2411",x"3b200e",x"3c210e",x"3b200e",x"3d210f",x"3d220f",x"3d220f",x"3c220e",x"3b200e",x"3b210e",x"3b220f",x"3c210e",x"39200e",x"371f0e",x"361e0d",x"341d0d",x"331c0c",x"341c0c",x"311b0b",x"39200e",x"351d0d",x"351d0d",x"381f0d",x"3d2310",x"351d0d",x"341e0d",x"2d1a0c",x"211409",x"170f07",x"150e07",x"160e07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503d30",x"503d30",x"38200e",x"3b210f",x"3c210f",x"39200e",x"3a210e",x"351e0d",x"381f0e",x"311b0c",x"331c0c",x"38200e",x"38200f",x"3c2310",x"38200f",x"341e0d",x"341d0d",x"331d0d",x"351e0d",x"2e1a0b",x"2e1a0c",x"321d0d",x"331d0d",x"331d0d",x"39210f",x"37200f",x"3a2210",x"3c2311",x"3c2310",x"38200f",x"36200e",x"39200f",x"331d0d",x"371f0e",x"341e0e",x"351e0d",x"341e0d",x"2e1a0b",x"37200f",x"321c0c",x"341d0d",x"351d0c",x"2e190b",x"2f1a0b",x"321c0c",x"331c0c",x"321c0c",x"2d190b",x"2f1b0c",x"311b0c",x"301b0c",x"2f1a0b",x"321c0c",x"2e1a0b",x"2f1a0b",x"2a180a",x"2c180a",x"2c190b",x"8d745a",x"967c5d",x"977d5f",x"897457",x"927a5c",x"856e53",x"91775d",x"8c7357",x"8e7559",x"8e7559",x"7a6349",x"2f1b0c",x"321e0c",x"301c0c",x"311d0c",x"321c0b",x"311c0c",x"311d0b",x"301c0b",x"301c0c",x"321e0c",x"37200d",x"36200c",x"37200e",x"351f0d",x"38210d",x"36200d",x"341f0c",x"3a240e",x"37220c",x"341f0c",x"321d0c",x"341f0c",x"38210e",x"3b230e",x"36200e",x"39220e",x"3a230f",x"38220e",x"2e1a0a",x"331d0d",x"301d0c",x"311d0c",x"29180b",x"301c0c",x"37210d",x"37210d",x"35200d",x"311d0b",x"331e0c",x"2b190a",x"2f1c0b",x"311d0b",x"321d0b",x"271809",x"321d0c",x"311c0c",x"321d0d",x"3f2511",x"25150a",x"25150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"221409",x"321e0e",x"361d0d",x"261509",x"29170a",x"2b180a",x"3f220f",x"432611",x"412511",x"452611",x"3d220e",x"3b200e",x"361e0d",x"492811",x"331d0d",x"28170a",x"241509",x"201309",x"211409",x"1d1208",x"231409",x"241509",x"201309",x"221409",x"23150a",x"1d1208",x"221409",x"1a1008",x"1c1108",x"170f07",x"1e1208",x"201208",x"1d1208",x"1d1208",x"180f07",x"221409",x"1a1008",x"211409",x"170f07",x"150e07",x"27160a",x"371f0e",x"3b220f",x"3b2210",x"432712",x"412511",x"39200f",x"36200e",x"412511",x"462913",x"3c2310",x"2b190c",x"1e1209",x"1b1108",x"150e07",x"1e1208",x"150e07",x"150e07",x"1b1108",x"1b1108",x"191008",x"150e07",x"1b1008",x"180f08",x"1d1208",x"191008",x"29180b",x"452712",x"2f1a0b",x"301a0b",x"150e07",x"221409",x"221409",x"000000",x"000000",x"482d1a",x"4d301b",x"4e301c",x"4d2f1a",x"482c19",x"472c1b",x"4d301d",x"4b2f1c",x"482b18",x"492d1a",x"472d1a",x"462c19",x"4d301d",x"4c2f1c",x"472d1a",x"462b1a",x"4b2f1b",x"472c1a",x"452a19",x"452a19",x"432817",x"402717",x"452a18",x"472c1a",x"472b19",x"422918",x"432918",x"422816",x"402716",x"442917",x"412717",x"3c2415",x"3a2315",x"412716",x"452916",x"3e2616",x"412816",x"432817",x"482b18",x"422714",x"442816",x"462a16",x"4a2d18",x"4a2c17",x"4b2d18",x"492c18",x"4a2d18",x"4a2d19",x"492b16",x"4a2c17",x"482a16",x"4e2f19",x"4d2e18",x"4b2c16",x"432714",x"442613",x"472814",x"492a15",x"442713",x"422613",x"472914",x"4c2e17",x"4f2f18",x"4a2b16",x"482a17",x"4b2d17",x"4b2d17",x"482a16",x"452916",x"4b2d19",x"492c18",x"4a2d19",x"482c19",x"482b18",x"4d2f1b",x"4c301c",x"4f311d",x"4e311c",x"54341e",x"543520",x"4d301d",x"4c2f1b",x"4a2e1c",x"4d311e",x"4e311e",x"4d311e",x"4c301d",x"4f311d",x"4d311f",x"462c1c",x"452a1a",x"4a2f1d",x"4c2f1d",x"50321f",x"50321d",x"4b2f1c",x"4a2e1b",x"472b1a",x"4b2d1b",x"412819",x"412717",x"472b18",x"4b2e1a",x"4a2d1a",x"482b18",x"492d19",x"4a2d19",x"4f2f18",x"4d2e19",x"503019",x"482b16",x"482b16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"17100a",x"17100a",x"17110a",x"17110a",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"1b1108",x"1f1209",x"2a190b",x"311b0c",x"3a200f",x"3f2310",x"432611",x"442712",x"462813",x"432511",x"442712",x"462813",x"452813",x"452812",x"442712",x"432712",x"412512",x"3e2310",x"3c210f",x"391f0e",x"3a200f",x"3a210f",x"3a210f",x"3d2310",x"3a200f",x"361d0d",x"361d0d",x"3a210f",x"3d2410",x"3f2411",x"3e2410",x"3f2410",x"402511",x"3f2310",x"3d210f",x"3e220f",x"3e220f",x"402310",x"422511",x"432611",x"412411",x"422712",x"422612",x"402511",x"3d2410",x"38200f",x"361f0f",x"331e0d",x"311c0c",x"2e1b0c",x"311c0d",x"37200f",x"38200f",x"38200f",x"361f0e",x"36200e",x"341d0d",x"341c0d",x"321c0c",x"331b0c",x"331c0c",x"391f0e",x"38200e",x"381f0e",x"381f0d",x"391f0d",x"3b200e",x"391f0d",x"381f0d",x"381f0d",x"371d0c",x"371d0c",x"391f0d",x"3b210f",x"3e230f",x"381f0d",x"351d0c",x"341c0c",x"321c0c",x"331c0c",x"341d0d",x"38200e",x"3a210e",x"3c220f",x"3d2310",x"3f2411",x"3b210f",x"39200e",x"351e0d",x"2b190b",x"221409",x"180f07",x"150e07",x"150e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463d34",x"463d34",x"361e0d",x"3a210f",x"3d2310",x"3c2310",x"3d2310",x"39200f",x"38200e",x"311c0c",x"341d0c",x"321c0c",x"311b0c",x"381f0e",x"38200e",x"38200e",x"3a210f",x"341e0d",x"3b2210",x"38200f",x"361f0e",x"331d0d",x"351f0e",x"38200f",x"3b2210",x"3a200f",x"37200f",x"331d0d",x"361f0e",x"361e0d",x"341e0d",x"311c0c",x"301b0c",x"301b0c",x"2c190b",x"2c190b",x"2e1a0b",x"331d0d",x"2d190b",x"321c0c",x"2f1a0b",x"341d0d",x"311b0c",x"2b180b",x"2b180a",x"2d180a",x"2d190b",x"2d190b",x"311c0c",x"321d0c",x"301b0c",x"361e0d",x"2e190b",x"2b180a",x"2d190b",x"2c180b",x"351e0d",x"331d0d",x"361f0e",x"3a210f",x"3f2411",x"412511",x"351e0e",x"371f0e",x"3c210f",x"402511",x"3c2310",x"331d0d",x"341d0d",x"2d190b",x"2e1a0b",x"2b1a0b",x"2b190a",x"271609",x"2d1a0b",x"36200c",x"2e1b0b",x"2c1a0b",x"361f0c",x"301c0c",x"3a220e",x"36200c",x"3b230d",x"351f0c",x"3a230e",x"3c250d",x"39230e",x"341f0b",x"3a220d",x"35200e",x"36200d",x"37210d",x"35200e",x"38210d",x"301c0c",x"321d0c",x"2c1a0b",x"2d1a0b",x"341f0c",x"301c0b",x"341f0d",x"2e1b0b",x"351e0c",x"301b0c",x"2e1b0b",x"301d0b",x"36200e",x"341f0d",x"2d1a0b",x"2d1b0b",x"2a190a",x"331e0c",x"2c1b09",x"2f1b0b",x"29180a",x"301a0b",x"351e0d",x"23150a",x"23150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"2a180b",x"341d0d",x"341c0d",x"331d0c",x"361e0d",x"361e0d",x"351d0d",x"381f0e",x"361e0d",x"371f0d",x"381f0d",x"3a200e",x"311a0b",x"3d220f",x"391f0d",x"3a200e",x"3a200e",x"381f0e",x"3c220f",x"3f2410",x"3c220f",x"3e2310",x"341c0c",x"3e2410",x"3b210f",x"39210f",x"371e0d",x"3c2310",x"351d0d",x"331d0d",x"381f0e",x"371f0e",x"3b210f",x"39200f",x"3d2410",x"38200f",x"371f0e",x"381f0e",x"3a210f",x"39200f",x"38200f",x"39200f",x"3a210f",x"3b2210",x"3a210f",x"3e2410",x"361f0e",x"38200f",x"381f0e",x"311c0c",x"351d0d",x"371e0d",x"381f0e",x"39200f",x"321d0d",x"39200f",x"3a210f",x"39200f",x"3c2311",x"3c2311",x"39210f",x"361f0e",x"3c2310",x"3a210f",x"3e2411",x"3c2311",x"3f2511",x"3a210f",x"321c0c",x"301b0b",x"150e07",x"150e07",x"150e07",x"000000",x"492c18",x"53321c",x"4d2f1b",x"57321b",x"4e2f1a",x"52321c",x"52321c",x"54331d",x"55341d",x"56351d",x"56351d",x"50321c",x"4e2f1b",x"492d1a",x"432818",x"4a2d1a",x"4a2d19",x"4b2d1b",x"4b2d1a",x"492b18",x"412717",x"452817",x"442716",x"452816",x"492b17",x"4c2d19",x"4d2d19",x"53311b",x"53331c",x"54331c",x"512f1a",x"502f1a",x"4f2e1a",x"482b18",x"4a2c19",x"4d2d19",x"4b2d19",x"482b19",x"4b2c18",x"4a2b16",x"4b2c18",x"4f2d17",x"512f1a",x"492b17",x"502e19",x"4d2d18",x"512f1a",x"523019",x"533119",x"512f18",x"462715",x"54311a",x"502f19",x"563319",x"543019",x"533019",x"4b2a14",x"58351b",x"4e2c16",x"4e2d16",x"4f2d17",x"553219",x"58351b",x"56321a",x"553119",x"523018",x"533118",x"56321b",x"55321b",x"55321a",x"512f19",x"56331c",x"54331b",x"55331c",x"57351d",x"56341c",x"4e2f1c",x"53321c",x"53321c",x"51311d",x"51301b",x"52331e",x"563520",x"553620",x"573620",x"55331d",x"5b3821",x"55361e",x"583821",x"53341d",x"53341f",x"52341f",x"4f321e",x"50331f",x"563520",x"56351f",x"4b2e1b",x"4b2d19",x"4a2c1a",x"4f2f1a",x"472a19",x"462918",x"482a17",x"452817",x"452815",x"4c2c17",x"512f19",x"4f2f19",x"4e2f1a",x"57341c",x"53331b",x"4d2e17",x"4d2e17",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"171009",x"171009",x"171009",x"171009",x"17110a",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"1c1108",x"1e1209",x"29180b",x"341d0d",x"3c220f",x"402511",x"432612",x"442712",x"432711",x"452812",x"442712",x"442712",x"412410",x"402410",x"3d210f",x"3a200e",x"3c210f",x"3d2210",x"3b2210",x"3b2210",x"38200f",x"38200f",x"3a2210",x"3b2210",x"3b2210",x"3b2310",x"3d2310",x"3c2310",x"3e2411",x"3f2511",x"3e2511",x"3b210f",x"391f0d",x"391f0d",x"3a200d",x"3c210d",x"3c210d",x"3b200e",x"3c210e",x"3a1f0d",x"381f0d",x"3b210e",x"422611",x"402511",x"3e2310",x"392110",x"351f0e",x"331d0d",x"301c0d",x"2e1b0c",x"301b0c",x"311b0c",x"321c0c",x"321b0c",x"321c0c",x"321c0b",x"311b0b",x"2e1a0a",x"2d190a",x"2d180a",x"2f190a",x"321c0b",x"351d0c",x"39200e",x"39200d",x"3f240f",x"3f2310",x"3e2310",x"3b200e",x"3b200e",x"3b200e",x"3b210d",x"381f0d",x"381f0d",x"3a200d",x"351d0d",x"331c0c",x"321c0c",x"2d180a",x"311b0c",x"321c0c",x"311b0c",x"361e0d",x"371f0e",x"3b210f",x"3d2310",x"3b210f",x"39200e",x"2c180a",x"2c1a0b",x"201309",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503f33",x"503f33",x"462813",x"4b2b15",x"492b14",x"482a14",x"432712",x"3a200e",x"391f0d",x"381d0d",x"391f0d",x"351d0c",x"351d0c",x"381e0d",x"381e0d",x"371e0c",x"3b200e",x"3c220f",x"422611",x"422712",x"432712",x"432712",x"402511",x"442712",x"402410",x"412511",x"3a200e",x"351e0d",x"361d0d",x"3a1f0e",x"3a200e",x"371e0d",x"331c0b",x"30190b",x"31190b",x"30190a",x"341c0b",x"351c0b",x"321c0c",x"361e0d",x"3c210f",x"3c220f",x"3b210f",x"361e0d",x"361e0d",x"361e0d",x"381f0d",x"351d0c",x"371e0d",x"351d0d",x"351d0d",x"341c0c",x"311b0b",x"311b0c",x"2d190b",x"321c0c",x"331c0c",x"361e0d",x"341d0d",x"361e0d",x"3a210f",x"402511",x"351e0d",x"2f1a0b",x"381f0e",x"39200f",x"39210f",x"3a210f",x"39200f",x"351e0d",x"38200f",x"361f0d",x"341d0d",x"361e0d",x"361f0e",x"331d0d",x"38200e",x"39210e",x"38210e",x"3f250f",x"3e240f",x"41270f",x"40260f",x"3c230f",x"3d2410",x"432810",x"3f250f",x"41270f",x"3d230f",x"3a210e",x"3f250f",x"3d240e",x"38200d",x"39210e",x"3a210e",x"38210e",x"301d0c",x"36200d",x"3d240f",x"38210f",x"3a220e",x"351f0e",x"3a210f",x"38200e",x"3c2410",x"38210f",x"3d240f",x"3b220f",x"3d2411",x"381f0d",x"2e1b0b",x"331c0c",x"2c180a",x"2e1a0a",x"301a0b",x"2f1a0b",x"3a1f0d",x"321b0c",x"321b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"1f1208",x"2c180b",x"2e1a0b",x"361e0d",x"351d0d",x"321c0c",x"321c0c",x"321c0c",x"341d0c",x"351d0d",x"351d0d",x"331c0c",x"371f0d",x"351d0d",x"39200e",x"3c220f",x"38200e",x"3b210f",x"38200e",x"3b2210",x"381f0e",x"351e0d",x"3a210f",x"2f190b",x"351e0e",x"311c0d",x"39210f",x"3a220f",x"331d0d",x"341d0d",x"321c0c",x"341d0c",x"311c0c",x"331d0d",x"381f0e",x"3c2310",x"3a2210",x"341f0e",x"3b2210",x"371f0d",x"38210f",x"341e0e",x"321c0d",x"311c0c",x"351e0d",x"331c0c",x"321c0d",x"321c0c",x"331d0d",x"301c0c",x"341c0d",x"341d0d",x"341d0d",x"341d0d",x"371f0e",x"331c0d",x"351e0d",x"311d0d",x"341e0d",x"361f0e",x"371f0e",x"311c0c",x"301b0c",x"351e0e",x"39200f",x"3a220f",x"3a2110",x"341d0d",x"331c0d",x"2a170a",x"150e07",x"150e07",x"150e07",x"000000",x"3e2616",x"492c18",x"4e2e18",x"4c2e19",x"4b2c19",x"55321c",x"4d2f1a",x"502f1a",x"4a2c17",x"4a2b19",x"4a2c19",x"57341d",x"4f301b",x"4c2c1a",x"4c2f1c",x"57351d",x"55341d",x"54321d",x"50301a",x"492b17",x"462917",x"462917",x"482b17",x"4b2c17",x"4f2e18",x"4e2e17",x"523019",x"55321c",x"4d2b16",x"4d2d19",x"512f1b",x"54331b",x"512f1b",x"512f1a",x"4b2c18",x"472a16",x"492b17",x"4a2c17",x"462915",x"472816",x"4e2d18",x"502d18",x"512f19",x"522f19",x"502f18",x"513119",x"522f1a",x"54321a",x"522f19",x"56331a",x"59331b",x"4d2c16",x"5b361a",x"5d371c",x"59351a",x"5a361c",x"58331a",x"543118",x"553118",x"553118",x"522f18",x"4c2b15",x"533018",x"543219",x"5a361b",x"613a1e",x"5c361c",x"5d361c",x"56331a",x"5d381d",x"54321b",x"4f2d18",x"59351b",x"502e18",x"56351d",x"52301b",x"56331c",x"58351d",x"5c381e",x"52301c",x"51301d",x"553520",x"59361f",x"56341e",x"56341f",x"583720",x"573620",x"553520",x"5c3920",x"51331f",x"51331e",x"4c301d",x"4b301c",x"50321d",x"53331d",x"4e311c",x"4c2f1c",x"4f2f1a",x"4c2d18",x"492c19",x"482b19",x"462a18",x"472a19",x"462917",x"462916",x"4c2c19",x"4b2b16",x"4b2c17",x"492c16",x"492b15",x"432714",x"4e2d16",x"4e2d16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"17100a",x"17100a",x"171009",x"17110a",x"17100a",x"17110a",x"171009",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"1d1208",x"201309",x"29180b",x"321c0c",x"3d2410",x"422612",x"3e230f",x"3e230f",x"402410",x"3f230f",x"422611",x"402410",x"422511",x"422611",x"3a200e",x"3b210e",x"3b210f",x"39200e",x"361e0d",x"331c0d",x"351e0e",x"361f0e",x"331d0d",x"351f0e",x"361f0e",x"341d0d",x"331d0d",x"361f0e",x"37200e",x"39220f",x"3c230f",x"3a210e",x"39200e",x"3c210e",x"3b200d",x"3c210e",x"3c220e",x"3d220f",x"3c210e",x"3a200e",x"3a200e",x"3b210e",x"3d220e",x"3a210e",x"361e0e",x"301b0c",x"2e190b",x"2c190b",x"2d190b",x"2c190b",x"2f1b0c",x"321c0c",x"37200e",x"39200f",x"38200f",x"37200e",x"351e0d",x"341e0c",x"331c0b",x"341d0c",x"351d0b",x"38200d",x"371f0c",x"361e0c",x"3b220e",x"3b210e",x"381f0d",x"381f0d",x"3b210e",x"3f230f",x"3c210d",x"3c220e",x"371e0d",x"361f0c",x"37200c",x"321c0c",x"321c0c",x"2e190b",x"2d190b",x"2d190b",x"311b0c",x"341d0d",x"371f0e",x"39200e",x"3a200f",x"3c2210",x"371e0e",x"371f0e",x"331d0d",x"241409",x"201309",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3d31",x"4e3d31",x"402410",x"50331d",x"472a14",x"472a14",x"563821",x"432813",x"533620",x"523520",x"3e230f",x"4c311d",x"381f0d",x"3b210f",x"4f331e",x"3f2411",x"563822",x"4e341e",x"422612",x"513520",x"412612",x"3e2411",x"4f3520",x"402411",x"4e341f",x"3a200e",x"3b210f",x"4a301c",x"39200e",x"3b200e",x"4d321e",x"381f0d",x"462d1a",x"351d0c",x"462d1a",x"361e0c",x"361e0d",x"371e0c",x"452c19",x"361e0d",x"321b0c",x"351d0d",x"331c0c",x"301a0b",x"301a0b",x"311b0b",x"311b0b",x"2e190a",x"452e1b",x"432d1b",x"301b0b",x"412a18",x"2b170a",x"2c180a",x"442d1a",x"422c1a",x"442c18",x"442c1a",x"301b0c",x"331d0c",x"4b321d",x"492f1c",x"432c1a",x"2a180b",x"331c0d",x"482f1c",x"351e0e",x"472d1a",x"3a210f",x"432c1a",x"472e1b",x"472e1b",x"351f0e",x"38200e",x"49301c",x"331e0d",x"39210e",x"48311d",x"36200e",x"4f351e",x"432810",x"4f341d",x"402510",x"51361e",x"3d240f",x"4e341d",x"39220e",x"4b311b",x"37200d",x"4d341f",x"3b230f",x"4f341e",x"3a230e",x"49301b",x"341e0c",x"48311d",x"442f1c",x"331e0c",x"36200d",x"472f1a",x"472f1b",x"472e1b",x"472f1b",x"49311b",x"422c19",x"351f0d",x"432c1a",x"432c1a",x"49311c",x"4b311c",x"311d0c",x"301c0c",x"432d1a",x"29170a",x"2d190b",x"2e190b",x"4e331d",x"351d0d",x"351d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"2c1a0b",x"39200f",x"3a210f",x"3f2310",x"3e2310",x"391f0e",x"3e230f",x"412511",x"3e230f",x"3e2310",x"3e2310",x"432612",x"3d2310",x"3f230e",x"3b200d",x"3b200d",x"3d210e",x"3e220e",x"422612",x"3c210f",x"3d2310",x"351d0d",x"381f0e",x"3a210f",x"381f0e",x"3d220f",x"371f0e",x"361f0e",x"341c0d",x"371e0d",x"3b210f",x"3a210e",x"351d0d",x"30190b",x"3a200e",x"412612",x"3a2210",x"3f2411",x"3f2511",x"3c230f",x"3c220f",x"3a220f",x"3f2411",x"3b2210",x"39200f",x"361e0d",x"381f0e",x"3d2411",x"3a2210",x"3c220f",x"371e0d",x"3a200e",x"412612",x"3e2310",x"3c2310",x"39210f",x"361f0e",x"3d230f",x"3e2310",x"422611",x"3e2310",x"3a210f",x"391f0e",x"3a200e",x"402511",x"3b2310",x"2f1c0d",x"211409",x"150e07",x"150e07",x"150e07",x"150e07",x"321f11",x"452a17",x"301f12",x"402615",x"492c19",x"482d18",x"4e2f1b",x"4e301a",x"57351d",x"54331c",x"50301a",x"5c381f",x"5a381f",x"59361f",x"52321c",x"4b2d18",x"4e2f1a",x"4f2e19",x"4e2f19",x"50301c",x"4e2f1b",x"502f19",x"5a351c",x"4d2d19",x"4c2c19",x"482916",x"462917",x"58341c",x"58361d",x"5b361e",x"5a371f",x"5a371c",x"5a351b",x"56331b",x"57341c",x"58331b",x"502f1a",x"4e2e19",x"4f2f1a",x"4d2c18",x"502f19",x"4b2d18",x"51321a",x"4e2e18",x"4f2e16",x"4d2c16",x"4f2d16",x"4e2d16",x"522f18",x"503119",x"512f18",x"4e2d17",x"5b351b",x"5b361b",x"563219",x"553118",x"512f17",x"502e17",x"523018",x"502d16",x"543118",x"59341a",x"542f17",x"492914",x"452612",x"4a2b16",x"5c371c",x"5d371c",x"5b361c",x"51301a",x"4d2d18",x"4f2f18",x"5b371d",x"5a371d",x"54321b",x"4f2f1b",x"4b2d19",x"5a371e",x"5e3a20",x"643c22",x"512f1b",x"56321c",x"5f3a21",x"583620",x"5a351d",x"553620",x"553520",x"52331e",x"53341f",x"53341f",x"4c301c",x"4e301c",x"482d1b",x"4c2e1c",x"4f311c",x"50321e",x"583820",x"54351e",x"5c3a20",x"51311c",x"4e2e1b",x"432918",x"472b18",x"492b18",x"462917",x"452917",x"4a2c18",x"4b2d17",x"4d2e18",x"4b2d18",x"4a2c18",x"422716",x"4f3017",x"4f3017",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130c",x"1a130c",x"19120c",x"19130c",x"19120b",x"171009",x"17100a",x"17110a",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"1d1208",x"1f1309",x"27170a",x"301c0d",x"371f0e",x"3b210f",x"402511",x"442713",x"422612",x"3f2310",x"3f2310",x"3f2410",x"452813",x"472a15",x"3c220f",x"361d0d",x"38200e",x"39210f",x"331d0d",x"341e0d",x"311c0d",x"2f1b0c",x"2f1b0c",x"301c0d",x"311c0d",x"2f1b0c",x"2f1b0c",x"2d190b",x"2f1a0c",x"351f0e",x"3b230f",x"392210",x"3f2611",x"3f2610",x"3f240f",x"3c220e",x"39200d",x"3b210e",x"3c210f",x"3a210e",x"3c210e",x"3a200f",x"3b220f",x"381f0e",x"351f0e",x"311c0d",x"2f1b0c",x"2d190b",x"2e1b0c",x"2f1c0d",x"331e0e",x"341d0d",x"351e0d",x"351d0d",x"331c0c",x"351e0d",x"361e0d",x"38200e",x"361f0d",x"38210e",x"361f0d",x"38200c",x"361f0c",x"39200e",x"3f2510",x"3f2510",x"3d2310",x"3f2410",x"3f250f",x"3f2510",x"3e230f",x"3e240f",x"3a210e",x"3a200e",x"3b230e",x"351e0d",x"311b0c",x"311c0d",x"2f1b0c",x"2f1b0c",x"2e1a0b",x"301b0b",x"311b0b",x"341d0c",x"371e0d",x"3a210f",x"39210f",x"361e0e",x"2d190b",x"27160a",x"1e1208",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3d31",x"402410",x"50331d",x"472a14",x"472a14",x"563821",x"432813",x"533620",x"523520",x"3e230f",x"4c311d",x"381f0d",x"3b210f",x"4f331e",x"3f2411",x"563822",x"4e341e",x"422612",x"513520",x"412612",x"3e2411",x"4f3520",x"402411",x"4e341f",x"3a200e",x"3b210f",x"4a301c",x"39200e",x"3b200e",x"4d321e",x"381f0d",x"462d1a",x"351d0c",x"462d1a",x"361e0c",x"361e0d",x"371e0c",x"452c19",x"361e0d",x"321b0c",x"351d0d",x"331c0c",x"301a0b",x"301a0b",x"311b0b",x"311b0b",x"2e190a",x"452e1b",x"432d1b",x"301b0b",x"412a18",x"2b170a",x"2c180a",x"442d1a",x"422c1a",x"442c18",x"442c1a",x"301b0c",x"331d0c",x"4b321d",x"492f1c",x"432c1a",x"2a180b",x"331c0d",x"482f1c",x"351e0e",x"472d1a",x"3a210f",x"432c1a",x"472e1b",x"472e1b",x"351f0e",x"38200e",x"49301c",x"331e0d",x"39210e",x"48311d",x"36200e",x"4f351e",x"432810",x"4f341d",x"402510",x"51361e",x"3d240f",x"4e341d",x"39220e",x"4b311b",x"37200d",x"4d341f",x"3b230f",x"4f341e",x"3a230e",x"49301b",x"341e0c",x"48311d",x"442f1c",x"331e0c",x"36200d",x"472f1a",x"472f1b",x"472e1b",x"472f1b",x"49311b",x"422c19",x"351f0d",x"432c1a",x"432c1a",x"49311c",x"4b311c",x"311d0c",x"301c0c",x"432d1a",x"29170a",x"2d190b",x"2e190b",x"4e331d",x"351d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"23150a",x"311c0c",x"37200e",x"361f0e",x"2f1b0c",x"2d190b",x"402511",x"2e1b0c",x"39210f",x"362310",x"37200e",x"37200e",x"331c0c",x"311c0c",x"2b180b",x"261509",x"381f0e",x"3e220f",x"371e0d",x"3e220f",x"3e230f",x"3c220f",x"3a200f",x"2d180a",x"2e190b",x"271609",x"2a180b",x"25160a",x"1d1108",x"1a1008",x"1a1008",x"1d1108",x"1d1108",x"1f1209",x"1f1209",x"1d1208",x"211409",x"1d1208",x"180f07",x"1f1309",x"211409",x"1f1209",x"1e1209",x"1d1209",x"221409",x"24160a",x"24150a",x"25160a",x"28180b",x"2c1a0c",x"26160a",x"2b190c",x"26160a",x"25160a",x"251509",x"26160a",x"231509",x"231509",x"28170a",x"321d0d",x"361e0e",x"321d0d",x"2c190b",x"24150a",x"27170a",x"251509",x"26160a",x"2d1a0c",x"27170a",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2d17",x"402513",x"352012",x"3f2616",x"4d2e19",x"452b19",x"4c2e19",x"53321b",x"4e301a",x"52321c",x"58371e",x"4f301c",x"51321b",x"4e2f19",x"4d301b",x"50311b",x"55341d",x"51321b",x"53321c",x"4d311b",x"54331d",x"4b2d18",x"502f19",x"472b18",x"442815",x"4f2e18",x"472a17",x"4e2f19",x"4f2f1a",x"56331c",x"54321b",x"4f2e19",x"52311a",x"5b371d",x"58331b",x"55331b",x"55321c",x"52311a",x"51301b",x"4f2f1a",x"53321b",x"59351d",x"492b16",x"402412",x"4b2b15",x"442814",x"492a15",x"4f2d17",x"4c2b16",x"3f2412",x"472814",x"58341b",x"4c2c16",x"4c2d17",x"5b361b",x"472814",x"4c2b16",x"5e381c",x"523119",x"4c2d17",x"55331a",x"613b1e",x"55331a",x"533119",x"4d2e18",x"56321a",x"512f19",x"52321a",x"5b381e",x"52331a",x"452815",x"472915",x"4c2c18",x"51311b",x"53321b",x"4d2d1b",x"59361e",x"54321c",x"56351e",x"59381f",x"55341d",x"55331d",x"492c19",x"53311c",x"53331e",x"50311c",x"50311c",x"442c1c",x"4c2f1c",x"50331f",x"573821",x"52321d",x"4e301c",x"4c2f1c",x"4e321e",x"4e311d",x"422919",x"482d1b",x"50321c",x"462c1b",x"492e1b",x"472d1a",x"492d1b",x"462c18",x"3f2717",x"432a19",x"492d1a",x"51321c",x"51311a",x"472c19",x"432816",x"422917",x"301e11",x"482915",x"482915",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19130b",x"19130b",x"19120b",x"19120b",x"19120b",x"1a130d",x"1a130c",x"171009",x"17110a",x"171009",x"17110a",x"150e07",x"150e07",x"1a1008",x"1a1008",x"1c1108",x"1d1208",x"24160a",x"2b190b",x"2d190b",x"361e0d",x"3c2210",x"402512",x"3c220f",x"412512",x"412612",x"412612",x"412612",x"422713",x"3a210f",x"341c0c",x"2f1a0b",x"301c0c",x"2d1a0b",x"2a180b",x"28170a",x"28170a",x"28170b",x"2a190b",x"2b190b",x"2a180b",x"2c1a0c",x"2c1a0c",x"2d1a0c",x"2c190c",x"2f1c0c",x"341f0e",x"38200f",x"3d240f",x"3e2410",x"3c2310",x"3b220f",x"37200e",x"38200e",x"38200f",x"3a2310",x"39220f",x"3a220f",x"361f0e",x"311c0d",x"2d1a0c",x"2b190b",x"29180b",x"28170a",x"28170a",x"2e1a0c",x"331e0e",x"38200f",x"38210f",x"38210f",x"37200f",x"341e0d",x"361f0d",x"361e0d",x"331d0c",x"39210c",x"37200d",x"361f0d",x"371f0d",x"3c230f",x"3c230f",x"3c230f",x"381f0d",x"3c230f",x"3d230f",x"3b220e",x"3a220e",x"37200e",x"3a220e",x"37200e",x"2e1a0b",x"2e1a0c",x"2a180b",x"271609",x"221408",x"28170a",x"2c180a",x"2f1a0b",x"321c0b",x"321c0b",x"2c180a",x"321c0b",x"311c0c",x"2e1b0c",x"25160a",x"1c1108",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"2f1a0c",x"2f1a0c",x"2c190b",x"170f07",x"26160a",x"301c0c",x"341e0d",x"361f0e",x"361f0e",x"341e0d",x"311c0d",x"321d0d",x"2f1a0b",x"341d0c",x"2b180a",x"341d0c",x"2a170a",x"2a1709",x"311b0b",x"2e1a0b",x"2c180a",x"2c190a",x"321c0b",x"291709",x"2d190b",x"2e1a0c",x"2d1a0c",x"29170a",x"382010",x"321d0e",x"2e1a0c",x"301b0c",x"301b0c",x"331d0d",x"2f1a0b",x"2f1a0c",x"311c0d",x"2e1b0c",x"301c0d",x"311c0d",x"301c0d",x"2c1a0c",x"331d0e",x"321d0e",x"2f1c0d",x"301c0d",x"331d0e",x"2c190c",x"341e0e",x"2d1a0c",x"331e0e",x"321d0e",x"2a180b",x"2c190b",x"29170a",x"29170a",x"2b180b",x"2c190b",x"28170a",x"29170a",x"2e1a0b",x"2b180b",x"2e1a0c",x"2d1a0b",x"2d1a0b",x"24150a",x"2c190b",x"2f1b0c",x"321d0d",x"2d1a0c",x"25150a",x"150e07",x"150e07",x"150e07",x"150e07",x"482a15",x"4b2c17",x"442a16",x"4b2d19",x"53331b",x"4e2f1a",x"59361e",x"50301a",x"53321a",x"4d2d19",x"57341c",x"57341c",x"4d2e19",x"56341c",x"54321b",x"51301a",x"59341b",x"502f1a",x"4c2d17",x"4e2e19",x"59341b",x"472a16",x"5b341c",x"4f2d19",x"4d2d19",x"53301a",x"55311a",x"53321b",x"55331b",x"4a2b17",x"4b2b18",x"533119",x"57341c",x"58351d",x"54331c",x"53321b",x"5a361e",x"51301a",x"55341c",x"492b17",x"462815",x"402512",x"492b15",x"4a2b15",x"402513",x"422714",x"452814",x"412512",x"3e2210",x"452712",x"472814",x"442712",x"543119",x"513017",x"502d16",x"4c2e16",x"513017",x"553219",x"563217",x"553117",x"512e16",x"4c2c15",x"4e2d15",x"4b2b13",x"513016",x"533017",x"56341a",x"57341a",x"543119",x"4c2f19",x"533219",x"53321a",x"533019",x"53321a",x"57351c",x"57351c",x"52321b",x"58351d",x"5b3a20",x"58351d",x"53311b",x"50301b",x"52311b",x"50301b",x"54321c",x"482c1a",x"4e2f1a",x"482c1a",x"492c1a",x"51321d",x"50311d",x"55341e",x"53331d",x"4d2f1c",x"492c1a",x"51311c",x"54331d",x"4f311c",x"482b18",x"492b18",x"52321c",x"52331c",x"56351d",x"4a2d19",x"51321a",x"51321b",x"57351d",x"52311a",x"4f2f19",x"4d2e17",x"482b16",x"492b16",x"3e2413",x"362010",x"482915",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130b",x"1a130b",x"19120b",x"19120b",x"19130c",x"1a130c",x"19130c",x"1a130c",x"171009",x"17110a",x"171009",x"150e07",x"150e07",x"1c1108",x"1c1108",x"201309",x"23150a",x"28170b",x"301c0d",x"38210f",x"3d2411",x"3c2210",x"3f2512",x"412512",x"402511",x"3f2511",x"422713",x"3e2310",x"3b210f",x"381f0e",x"341d0d",x"321c0c",x"311b0c",x"2f1a0b",x"2c190b",x"2b180b",x"29170a",x"29170a",x"2a180b",x"2a180b",x"2a180b",x"29180b",x"28170a",x"28170a",x"2a190b",x"37220d",x"2d1a0b",x"2d1a0b",x"321d0c",x"39220f",x"3c2410",x"3a230f",x"3a210f",x"38210f",x"3b2410",x"3a220f",x"3a220f",x"3a210f",x"38200f",x"331d0d",x"2c190b",x"2a180b",x"2a180b",x"2a190b",x"2a180b",x"2d1a0b",x"311c0c",x"341d0d",x"351e0e",x"351e0e",x"341e0d",x"341d0c",x"351e0d",x"341d0c",x"331d0c",x"38200d",x"3a210d",x"39210e",x"361f0d",x"371f0d",x"371f0d",x"38200e",x"37200d",x"38200e",x"39210e",x"3e2510",x"3b220f",x"39210e",x"37200e",x"38210f",x"2d190b",x"2b180a",x"221308",x"251509",x"221409",x"211308",x"261609",x"29170a",x"29170a",x"2a1709",x"311b0b",x"2d190a",x"2e190b",x"2b190b",x"231509",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3b210f",x"3b210f",x"38200e",x"28170a",x"36200e",x"3a2110",x"37200f",x"3b2210",x"37200f",x"3a2210",x"2f1a0c",x"2d190b",x"321c0c",x"2f1a0b",x"311b0b",x"2e190a",x"331c0c",x"331c0c",x"321c0b",x"331c0c",x"311b0b",x"2f1a0b",x"2e190a",x"331c0c",x"2d190a",x"301c0d",x"2b180b",x"38200f",x"321d0d",x"311c0c",x"2e1b0c",x"301b0c",x"331d0d",x"321c0d",x"341d0d",x"2d190b",x"311c0c",x"341e0d",x"341e0d",x"331d0d",x"341e0e",x"321d0e",x"321d0e",x"2f1b0c",x"311c0d",x"2f1b0c",x"311c0d",x"2a180b",x"311c0d",x"27170a",x"2d190b",x"2a180b",x"29170a",x"251409",x"271509",x"221308",x"241409",x"251509",x"1e1007",x"1c1008",x"221208",x"261409",x"2a170a",x"281609",x"251409",x"251409",x"231308",x"261409",x"2b180a",x"281609",x"1f1208",x"180f08",x"150e07",x"150e07",x"150e07",x"492b16",x"452815",x"4d2d17",x"523119",x"53311a",x"55331c",x"53311a",x"502f19",x"513019",x"5a361c",x"54321a",x"58351c",x"513019",x"512f1a",x"55321b",x"52301a",x"54311b",x"54321b",x"53311b",x"56341b",x"59351c",x"502f1a",x"4e2e19",x"502e17",x"4c2c19",x"4a2b16",x"4d2d18",x"513019",x"56341b",x"54321a",x"54321b",x"57351c",x"55341d",x"52311b",x"53321b",x"54331d",x"50301a",x"522f19",x"442714",x"4c2c16",x"422512",x"502d16",x"3f2312",x"4a2b15",x"4f2d17",x"4b2b14",x"4e2c14",x"4e2d15",x"4b2b14",x"412512",x"4c2c15",x"402412",x"4f2d15",x"512f17",x"533118",x"543218",x"4b2b14",x"522f17",x"523016",x"513017",x"533017",x"533017",x"4b2a13",x"4e2d15",x"533118",x"593519",x"553218",x"563218",x"58341a",x"57351b",x"563118",x"533118",x"55331a",x"59341b",x"523119",x"553219",x"4e2d19",x"4d2e19",x"512f1a",x"4c2d18",x"472715",x"452817",x"472918",x"452917",x"452917",x"422618",x"331f15",x"3f2516",x"402718",x"472a19",x"4a2c1a",x"472b19",x"442717",x"432516",x"432615",x"4b2b18",x"482b18",x"4d2e1a",x"4e2d18",x"55341c",x"54331d",x"54331c",x"4e2f1a",x"54311b",x"4c2d19",x"56341b",x"4e2f19",x"54321b",x"4d2d18",x"4a2b16",x"4c2c17",x"502f18",x"462914",x"382111",x"382111",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"1b150e",x"1b150e",x"19130c",x"1a130c",x"19120c",x"1a130c",x"19120c",x"171009",x"171009",x"150e07",x"1e1209",x"1e1209",x"241509",x"29180b",x"2e1b0d",x"351f0f",x"39200f",x"402511",x"3e230f",x"3b200e",x"412410",x"412511",x"402410",x"3e220f",x"3e220f",x"381d0c",x"371c0c",x"351c0c",x"351b0b",x"351b0b",x"341b0b",x"251107",x"2f170a",x"2f1709",x"311a0a",x"321a0b",x"341c0c",x"311a0b",x"2e180a",x"2a1509",x"2e180a",x"331d0b",x"37200c",x"3a210c",x"3c230f",x"3e250f",x"412610",x"442811",x"422610",x"3f230f",x"3e2310",x"442812",x"432712",x"422611",x"3c220f",x"3b210e",x"3c220f",x"38200e",x"38200f",x"37200e",x"361f0e",x"361e0d",x"38200e",x"3a200e",x"3c220f",x"3b210f",x"3c220f",x"3a210f",x"3c230f",x"351e0c",x"371e0d",x"341d0c",x"3b220e",x"361e0d",x"37200c",x"39210e",x"3b220f",x"39210e",x"3e240f",x"3d240f",x"3d240f",x"3c220f",x"3d2410",x"3e2510",x"3c240f",x"3b220e",x"341d0c",x"331c0c",x"2a170a",x"301b0b",x"281609",x"2f1a0b",x"321c0c",x"321c0b",x"331c0b",x"351d0c",x"331c0b",x"2e190a",x"391f0d",x"2d1a0c",x"341e0f",x"2b180b",x"27170b",x"1f1309",x"191008",x"160e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3a200f",x"3a200f",x"351c0c",x"29170a",x"351e0d",x"38200f",x"39200f",x"3a210f",x"371f0e",x"381f0e",x"38200e",x"351e0d",x"2e190a",x"341d0c",x"301b0b",x"331c0c",x"331c0c",x"291709",x"2e190a",x"321b0b",x"331c0c",x"341c0c",x"2b180a",x"351d0c",x"2e1a0a",x"331d0d",x"351e0e",x"361f0e",x"341d0d",x"311b0c",x"2f1b0c",x"351d0d",x"331c0c",x"321c0c",x"311c0c",x"321b0c",x"3a210f",x"341d0d",x"301b0c",x"301a0b",x"311b0c",x"361e0d",x"351e0e",x"351f0e",x"37200f",x"351f0f",x"37200f",x"341d0d",x"311c0c",x"2d190b",x"301b0c",x"2e1a0b",x"301b0c",x"2d190b",x"2d190b",x"301c0c",x"2d1a0b",x"331d0d",x"381f0e",x"321c0d",x"331d0d",x"361f0e",x"392110",x"361e0e",x"321c0d",x"2f1a0b",x"311b0c",x"331d0d",x"331d0d",x"331d0d",x"301c0c",x"27170a",x"150e07",x"150e07",x"150e07",x"543117",x"59341b",x"4d2f18",x"4c2d17",x"4b2c17",x"462715",x"452713",x"452613",x"402412",x"442613",x"462814",x"472814",x"462814",x"462814",x"4b2c15",x"462814",x"432614",x"442713",x"462915",x"462914",x"4c2d17",x"4e2f18",x"4f2f18",x"4b2c16",x"4c2d17",x"442713",x"452714",x"482915",x"492a16",x"442713",x"402311",x"472914",x"482a15",x"462a15",x"432815",x"3f2413",x"422714",x"402513",x"422613",x"3d2211",x"412512",x"3a2110",x"422512",x"3c2211",x"3c2211",x"331c0d",x"3a200e",x"412410",x"452612",x"3a200e",x"422511",x"3d220f",x"442611",x"452814",x"422612",x"422511",x"402410",x"422512",x"482914",x"472912",x"402311",x"402411",x"3f230f",x"432613",x"432612",x"4a2b14",x"442612",x"422411",x"432612",x"482914",x"472a15",x"502f17",x"502f18",x"513019",x"4e2d17",x"492c16",x"472916",x"482a16",x"4c2c18",x"4c2e19",x"492b17",x"482b17",x"4e2f1a",x"4b2d19",x"4e301a",x"4d2e1a",x"51311c",x"50311b",x"51311a",x"55341d",x"54321c",x"4c2e1a",x"4d2d19",x"4c2d18",x"50301a",x"54331c",x"54331c",x"54331c",x"54341b",x"56341c",x"56351d",x"56341c",x"54331c",x"53311b",x"52311a",x"4b2d18",x"4b2c17",x"472a14",x"422612",x"422613",x"412513",x"422511",x"482914",x"3e2411",x"3e2411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"1c150e",x"1c150e",x"1b140d",x"1b140d",x"1a130c",x"19120b",x"19130c",x"1a130c",x"171009",x"150e07",x"1e1209",x"1e1209",x"211309",x"251509",x"331d0d",x"3b210f",x"432712",x"452813",x"472914",x"482a14",x"452712",x"432611",x"422411",x"432511",x"442611",x"452611",x"422410",x"432511",x"472912",x"492a14",x"482913",x"462712",x"472813",x"462812",x"4a2b14",x"4a2b14",x"452711",x"412410",x"3d220f",x"3c210f",x"412511",x"402510",x"482a13",x"4a2b13",x"472a12",x"4b2c14",x"4c2c14",x"4e2f15",x"4c2d15",x"4c2b14",x"4a2b14",x"482913",x"462712",x"40230f",x"3f230f",x"3d210e",x"3b200d",x"3d210e",x"3d210f",x"3d210f",x"3e230f",x"3f230f",x"3d220f",x"3e230f",x"3e220f",x"40240f",x"412411",x"402410",x"442811",x"472a14",x"452812",x"432711",x"432611",x"3f240e",x"3e230f",x"3f250f",x"3f240f",x"3d230e",x"3d220e",x"432711",x"432611",x"442811",x"482a13",x"422610",x"432710",x"412510",x"432611",x"341c0b",x"3e220e",x"321b0b",x"3c210e",x"3b200e",x"351d0c",x"331c0b",x"371e0c",x"3e220e",x"3f230f",x"371d0c",x"41240f",x"371e0d",x"3f2412",x"3d2310",x"371f0e",x"2d190b",x"1d1108",x"160f07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"38200e",x"38200e",x"3c220f",x"301b0c",x"392110",x"412611",x"482a13",x"482812",x"472712",x"432511",x"462712",x"442610",x"452610",x"3c200d",x"40230f",x"44260f",x"3b200c",x"381e0c",x"371e0b",x"3b200d",x"43240f",x"41230f",x"321b0b",x"341d0c",x"321c0b",x"321c0c",x"331c0d",x"2e190b",x"361e0d",x"341c0c",x"311b0b",x"2d190b",x"311b0b",x"3a1f0d",x"3c210e",x"3b200e",x"3e220f",x"402310",x"412410",x"462812",x"472812",x"452712",x"432511",x"432611",x"3f2410",x"3e2310",x"402511",x"432611",x"452712",x"412511",x"432611",x"412511",x"3c220f",x"402410",x"412410",x"3e2410",x"3f2410",x"3f2410",x"402410",x"331d0d",x"371f0e",x"39210f",x"39200f",x"3c220f",x"391f0d",x"351e0d",x"2c190b",x"301b0c",x"311c0c",x"2c190b",x"221409",x"1f1208",x"150e07",x"150e07",x"150e07",x"452711",x"3c220f",x"321d0d",x"2f1a0d",x"301a0d",x"311c0d",x"321c0d",x"301b0d",x"311c0d",x"331c0e",x"331c0d",x"301c0d",x"311b0d",x"321b0d",x"301c0d",x"321c0d",x"331c0d",x"331d0e",x"331d0e",x"321d0e",x"321d0e",x"321d0e",x"382010",x"372010",x"361e0f",x"3b2211",x"392110",x"382010",x"3a2111",x"392110",x"3a2210",x"392111",x"382011",x"361f10",x"321d0f",x"301c0e",x"2e1b0d",x"2c1a0d",x"301b0d",x"2a190b",x"2d1a0c",x"2a190c",x"2c1a0c",x"25160b",x"21150a",x"25160b",x"23150b",x"241509",x"2a170a",x"261609",x"2e190b",x"251509",x"28170a",x"28170a",x"29160a",x"26150a",x"241409",x"271509",x"28160a",x"2c180a",x"2b180a",x"2a170a",x"2a170a",x"2b180a",x"2f1b0c",x"311c0c",x"311c0c",x"311c0c",x"331d0d",x"311d0e",x"361f0f",x"341e0f",x"351e0f",x"351e0f",x"382010",x"351f0f",x"382112",x"382111",x"3a2211",x"3b2312",x"372011",x"372011",x"3b2312",x"3c2514",x"372012",x"392213",x"432816",x"402714",x"422716",x"442916",x"442915",x"3f2414",x"422715",x"3e2412",x"422613",x"422614",x"3f2413",x"402513",x"432613",x"412614",x"442914",x"432814",x"432814",x"402412",x"371e0f",x"361d0e",x"321b0d",x"301a0d",x"2e1a0c",x"2e1b0c",x"2c1a0c",x"2f1c0d",x"3c210e",x"402411",x"402411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1610",x"1d1610",x"1d1710",x"1b150e",x"1b140d",x"1b140d",x"1b150e",x"1c150f",x"19130c",x"19130c",x"19120b",x"171009",x"150e07",x"1d1108",x"1d1108",x"231509",x"29170b",x"321d0d",x"3b210f",x"412410",x"432611",x"422511",x"452712",x"452711",x"472812",x"472812",x"472912",x"472812",x"462711",x"472712",x"462712",x"492a13",x"462712",x"472712",x"492a14",x"472812",x"452812",x"462813",x"482a14",x"422511",x"3f220f",x"3e220f",x"3d210f",x"412410",x"3c210e",x"422610",x"452711",x"462911",x"472912",x"492a12",x"482913",x"482912",x"41240f",x"3f220f",x"391e0d",x"3b200c",x"3b200d",x"3c200d",x"3a1f0d",x"3d210e",x"3d220f",x"3a1f0d",x"371d0c",x"391e0d",x"381e0d",x"381e0d",x"3a1f0d",x"3f220f",x"3f230f",x"40230f",x"40240f",x"3d220f",x"432610",x"432711",x"422611",x"492b12",x"472a12",x"452811",x"432711",x"432811",x"422610",x"472911",x"442812",x"4a2c14",x"482a12",x"452811",x"442710",x"3f230e",x"442711",x"44260f",x"3c210e",x"3b200d",x"3c210d",x"3d210e",x"361e0c",x"331c0b",x"341c0b",x"361e0c",x"3e220e",x"42240f",x"371d0b",x"43250f",x"39200e",x"3b2110",x"3a200e",x"2f1a0b",x"2d190b",x"1b1008",x"1b1008",x"190f08",x"190f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"432611",x"432611",x"402411",x"321c0d",x"3f2512",x"3e230f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"381f0d",x"150e07",x"331c0c",x"271509",x"150e07",x"150e07",x"150e07",x"150e07",x"371e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"391f0d",x"251509",x"180f07",x"301a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"2b180a",x"1f1208",x"150e07",x"221409",x"1d1108",x"150e07",x"150e07",x"150e07",x"462911",x"3f240f",x"2d1a0b",x"2c1a0a",x"28160a",x"28160a",x"2a180a",x"261609",x"27160a",x"28160a",x"29170a",x"28160a",x"271609",x"29170a",x"2a180a",x"2a180a",x"28160a",x"28160a",x"29170a",x"28170a",x"28160a",x"28170a",x"2b180b",x"2c180b",x"2e1a0b",x"301b0c",x"301b0c",x"301b0c",x"2f1b0c",x"2f1b0c",x"2d1a0b",x"2c190b",x"2c190b",x"2b190b",x"2a180b",x"26160a",x"231409",x"231409",x"241509",x"201308",x"201308",x"1d1108",x"1e1208",x"1c1108",x"1a1008",x"190f07",x"190f07",x"190f07",x"180f07",x"180f07",x"190f07",x"190f07",x"180f07",x"191008",x"180f07",x"180f07",x"180f07",x"190f07",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"211309",x"201309",x"231409",x"24150a",x"24150a",x"24150a",x"211309",x"221409",x"231409",x"241509",x"251509",x"241509",x"241409",x"261509",x"28160a",x"28170a",x"29170a",x"2a170a",x"2a180a",x"2c180a",x"2f1a0b",x"311b0b",x"331c0c",x"341d0c",x"351d0d",x"341c0c",x"311b0b",x"311b0b",x"321b0c",x"321b0b",x"351d0c",x"351d0d",x"371e0d",x"371e0d",x"341c0c",x"331c0c",x"331c0c",x"331c0c",x"321c0c",x"311b0c",x"2d190b",x"2a170a",x"28160a",x"27160a",x"231409",x"1e1208",x"1d1108",x"2e1a0b",x"432511",x"432511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1d1610",x"1d1710",x"1c160f",x"1c160f",x"1b150e",x"1c150e",x"1b140d",x"1b150e",x"19130c",x"17110a",x"150e07",x"1e1208",x"1e1208",x"221409",x"2a180b",x"321d0d",x"38200f",x"361e0d",x"351d0d",x"3a200e",x"3c210f",x"3d210f",x"3c210e",x"3a1f0d",x"381e0c",x"3b200d",x"3e220f",x"3f230f",x"3f230f",x"3e220e",x"3e220f",x"3e210e",x"3f230f",x"3f230f",x"40230f",x"402310",x"3f220f",x"3b200e",x"391e0d",x"381d0c",x"361d0c",x"371e0d",x"3a200d",x"3d220e",x"41260e",x"3f240e",x"40240f",x"40240f",x"412510",x"3f240e",x"40240f",x"3c200e",x"40230f",x"3b200e",x"3e220e",x"40240f",x"361d0c",x"381f0d",x"3a200e",x"3b210e",x"361d0c",x"351c0c",x"381e0d",x"3b200e",x"3b200e",x"361e0c",x"3b200e",x"3c210f",x"3b210e",x"3b220e",x"3d230f",x"42260f",x"38200d",x"40250f",x"3c230e",x"3b220f",x"3c230e",x"361f0d",x"3c220f",x"3b220e",x"3c220e",x"3c220f",x"422610",x"462a11",x"3d230e",x"3a1f0d",x"3b210e",x"3d230e",x"371e0d",x"371f0e",x"391f0e",x"3b200d",x"361d0c",x"341c0b",x"331c0b",x"381e0d",x"3e220e",x"361e0c",x"3a200d",x"3a200f",x"3f2310",x"3e2311",x"3b2211",x"2d180b",x"28150a",x"1c1108",x"160f07",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"442611",x"442611",x"442712",x"321c0d",x"3e2411",x"381e0d",x"211308",x"2c190b",x"2b180b",x"2d190b",x"2c180b",x"2c180a",x"2a170a",x"2a170a",x"261509",x"241509",x"211309",x"251509",x"2d190b",x"29170a",x"271609",x"2c190a",x"1f1208",x"150e07",x"150e07",x"150e07",x"38200e",x"180f07",x"1e1108",x"211309",x"1e1208",x"150e07",x"150e07",x"502d14",x"2c190b",x"201309",x"251509",x"261509",x"28160a",x"251509",x"28170a",x"26160a",x"2d190b",x"2d1a0b",x"28170a",x"29180b",x"2b190b",x"2c1a0b",x"27170a",x"221409",x"221308",x"251409",x"221309",x"27160a",x"26160a",x"261609",x"251509",x"201309",x"150e07",x"150e07",x"2f1a0b",x"422510",x"150e07",x"1d1108",x"27160a",x"211409",x"150e07",x"150e07",x"4b2b14",x"150e07",x"1b1008",x"1f1208",x"150e07",x"150e07",x"150e07",x"3f240f",x"2d1b0b",x"2d1b0b",x"2c190b",x"2e1b0b",x"29170a",x"271609",x"271509",x"261509",x"251509",x"261509",x"281609",x"2a180a",x"2c190b",x"2d190b",x"2d1a0b",x"2c190b",x"2a170a",x"29170a",x"29170a",x"29170a",x"29170a",x"29160a",x"2a170a",x"2d180a",x"2d190a",x"2e190b",x"311b0b",x"311c0c",x"2f1a0b",x"2f1a0b",x"2d190b",x"2d190b",x"2c180a",x"2b180a",x"2e1a0b",x"2a170a",x"2c190b",x"2a180a",x"231409",x"28170a",x"211308",x"241509",x"241509",x"221409",x"201309",x"1f1208",x"1d1108",x"1c1108",x"1f1208",x"1d1108",x"201309",x"1d1108",x"1e1208",x"1f1208",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"201309",x"221409",x"231509",x"231409",x"221409",x"231409",x"231409",x"241509",x"26160a",x"27160a",x"28170a",x"28170a",x"28170a",x"2a180b",x"2b190b",x"2b190b",x"2b190b",x"29170a",x"241409",x"251409",x"271509",x"28170a",x"2c190b",x"2d190b",x"2f1b0c",x"321c0c",x"361f0e",x"361e0d",x"371e0d",x"381f0d",x"3b210e",x"3b200e",x"3a200e",x"3c210f",x"3c210f",x"3c210e",x"3e2310",x"3f2310",x"3d220f",x"3d220f",x"3d2210",x"3b210f",x"371e0d",x"39200e",x"371f0e",x"341d0d",x"311c0c",x"301b0c",x"2c190b",x"261509",x"221309",x"1f1208",x"1b1008",x"180f07",x"381f0f",x"381f0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d160f",x"1d160f",x"1e1711",x"1c160f",x"1d1710",x"1d160f",x"1e1811",x"1b140d",x"1b150e",x"1b140d",x"19130c",x"171009",x"150e07",x"1e1209",x"1e1209",x"231409",x"29170a",x"2d190b",x"341d0d",x"38200e",x"38200e",x"3a220f",x"3e2310",x"3d2310",x"3e2310",x"341b0b",x"33190a",x"361c0c",x"3a1f0d",x"3e230f",x"402310",x"3f230f",x"422511",x"432611",x"452711",x"412410",x"40230f",x"422410",x"412410",x"3f230f",x"402310",x"3e230f",x"3a200e",x"3b210f",x"3e2410",x"412610",x"422710",x"452711",x"442811",x"412510",x"452810",x"3f240f",x"3f230f",x"3f230f",x"3f230f",x"3c210e",x"3b210d",x"381e0c",x"3a200d",x"341c0b",x"321a0b",x"341b0b",x"331c0b",x"341d0c",x"361e0d",x"371e0d",x"371e0d",x"351d0d",x"341c0c",x"351d0c",x"381f0d",x"331c0b",x"361f0c",x"361f0b",x"36200b",x"36200c",x"341f0b",x"351f0c",x"331d0c",x"2b190a",x"2d1a0b",x"2f1a0b",x"2e1a0a",x"311b0b",x"311c0b",x"371f0d",x"3c220e",x"341d0b",x"38200c",x"39200d",x"311c0d",x"351e0e",x"2e1b0d",x"361e0e",x"351d0c",x"381f0d",x"311b0b",x"331c0c",x"301b0b",x"331c0b",x"371e0d",x"371e0e",x"3b2312",x"381f10",x"392110",x"321c0c",x"251509",x"1e1208",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"522f16",x"4a2a13",x"472812",x"452711",x"432510",x"432510",x"452712",x"422511",x"432611",x"482912",x"442611",x"3f230f",x"3b200d",x"3d210e",x"3f220f",x"3f220f",x"412410",x"3b200e",x"3f230f",x"3f230f",x"3f230f",x"3c210e",x"3d220f",x"3d220f",x"3c210e",x"3d220f",x"3e220f",x"3e220f",x"3f2310",x"3e230f",x"3c210f",x"3f230f",x"3f230f",x"3c210e",x"3d220e",x"3a1f0e",x"39200d",x"371e0d",x"381e0d",x"371d0c",x"361d0c",x"361d0c",x"361d0c",x"381e0d",x"381f0d",x"391f0e",x"391f0d",x"391f0d",x"391f0d",x"361d0d",x"361d0d",x"361d0c",x"371e0d",x"351c0c",x"2f1a0b",x"341c0c",x"371e0d",x"371e0d",x"371e0c",x"381f0d",x"361e0d",x"371d0c",x"331b0b",x"321a0b",x"381f0d",x"3c210f",x"381f0d",x"3b200e",x"3c210e",x"391f0d",x"3f2310",x"3e230f",x"381f0c",x"39200d",x"3b200d",x"391f0d",x"391f0d",x"381f0d",x"3b210e",x"3b200e",x"381f0c",x"3c210e",x"351d0d",x"3c220f",x"391f0e",x"3b210e",x"371f0d",x"381f0e",x"3c210e",x"3b200e",x"371e0d",x"351d0c",x"361d0d",x"381f0d",x"371e0d",x"3a200e",x"3a200e",x"3a200f",x"3a200e",x"3a210f",x"3a200e",x"39200e",x"3b220f",x"38200f",x"3d220f",x"39200e",x"381f0d",x"39200e",x"3a200e",x"3a210f",x"3a200e",x"3a210f",x"3d220f",x"39200e",x"361d0d",x"361d0c",x"341c0c",x"361e0d",x"39200e",x"39200e",x"361e0d",x"38200e",x"371f0e",x"311b0c",x"331c0c",x"3a210e",x"39200e",x"3a200e",x"3b200e",x"3a200e",x"3a200e",x"391f0e",x"351d0d",x"361e0d",x"3a200f",x"371f0e",x"3a200e",x"381f0e",x"351d0d",x"361e0d",x"341d0d",x"331c0c",x"331c0c",x"351d0c",x"361d0d",x"351d0d",x"371f0d",x"361e0d",x"371f0d",x"371f0d",x"341d0c",x"331c0c",x"351d0d",x"361d0d",x"341c0c",x"331c0c",x"361e0d",x"331d0c",x"3a200e",x"422511",x"371e0e",x"000000"),
(x"442712",x"442712",x"452813",x"321c0d",x"402511",x"432611",x"2e1b0c",x"321c0d",x"321c0c",x"331c0d",x"2e190b",x"2d190b",x"2b180a",x"301b0b",x"2d190b",x"281609",x"261509",x"2c180a",x"281609",x"2c190a",x"321c0b",x"281609",x"2c180a",x"1d1108",x"150e07",x"3f220e",x"28170a",x"231409",x"241409",x"261509",x"261509",x"1d1108",x"150e07",x"150e07",x"442711",x"1f1309",x"29180a",x"28170a",x"28160a",x"29170a",x"301b0c",x"2e1a0b",x"321c0d",x"321c0c",x"2e1a0b",x"2e1a0c",x"2c190b",x"2d1a0b",x"2e1a0c",x"2e1a0c",x"29180a",x"2c190b",x"2c190b",x"29180b",x"28170a",x"2a180b",x"29170a",x"26160a",x"231509",x"150e07",x"3b200e",x"311b0c",x"231509",x"25150a",x"2c190b",x"29180a",x"25150a",x"150e07",x"150e07",x"3b2210",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301d0c",x"311c0c",x"2d190b",x"301c0c",x"2f1a0b",x"2c180a",x"2b170a",x"29160a",x"271509",x"2b170a",x"2c190b",x"2c180a",x"2a170a",x"2b170a",x"2d190b",x"2f1a0b",x"2d190b",x"2d190b",x"2e1a0b",x"301b0b",x"351d0d",x"39210f",x"3a210f",x"3b210f",x"3a200e",x"381e0d",x"371e0d",x"3a200e",x"351c0c",x"361e0c",x"38200e",x"3b210f",x"3c220f",x"3c220f",x"3a210f",x"2e180a",x"371f0d",x"371f0e",x"331c0c",x"301a0b",x"331c0c",x"2d190a",x"291709",x"291709",x"271609",x"291709",x"2e1a0b",x"2c180a",x"2d190a",x"2b180a",x"2d190b",x"2a170a",x"2d190b",x"29170a",x"271509",x"281609",x"271609",x"28160a",x"27160a",x"29170a",x"2a180b",x"2b180b",x"2b190b",x"2b180b",x"2b180b",x"2b180b",x"2e1a0c",x"2c190b",x"2f1b0c",x"2e1a0b",x"2e1a0c",x"2f1b0c",x"301b0c",x"2d190b",x"301c0c",x"2f1b0c",x"301b0c",x"2f1b0c",x"2e1a0b",x"2f1b0c",x"311c0c",x"311b0c",x"341d0d",x"331c0c",x"39200e",x"3a210e",x"361e0d",x"391f0e",x"3d220f",x"3e2310",x"3d220f",x"3d220f",x"3f2310",x"3f2410",x"412411",x"422611",x"432612",x"432612",x"422611",x"3e2310",x"391f0e",x"361d0d",x"351c0c",x"361d0d",x"361e0d",x"351d0d",x"311b0c",x"2a170a",x"251509",x"211308",x"1d1108",x"1a1008",x"3f2411",x"26160a",x"28170a",x"2d1a0b",x"2e1a0c",x"2e1a0b",x"2e190b",x"311c0d",x"321d0d",x"2f1c0d",x"2a180b",x"29180b",x"29170a",x"28170a",x"26160a",x"241509",x"201309",x"1d1108",x"1c1008",x"1c1008",x"1e1108",x"241509",x"28170a",x"2d190b",x"311c0c",x"321d0d",x"301b0c",x"29170a",x"2d1a0b",x"29170a",x"29170a",x"241509",x"211308",x"211308",x"201308",x"231409",x"27160a",x"221409",x"201309",x"190f07",x"502f18",x"1e1711",x"1e1711",x"1f1912",x"1f1812",x"1d1710",x"1d1610",x"1d1710",x"1d1710",x"1c150f",x"1b150e",x"1c150f",x"17110a",x"150e07",x"22160d",x"22160d",x"29190e",x"2d1b0f",x"311e10",x"341f11",x"341f10",x"382212",x"3a2212",x"3b2211",x"3e2513",x"402513",x"412514",x"3f2512",x"402513",x"3e2312",x"432815",x"432714",x"442814",x"3f2412",x"422613",x"442814",x"412512",x"3d2312",x"432714",x"422614",x"422713",x"3f2412",x"3e2412",x"3d2313",x"3d2412",x"412613",x"402713",x"432914",x"462b15",x"442815",x"442914",x"3f2412",x"3b2211",x"3e2412",x"3e2413",x"412612",x"3f2512",x"3b2211",x"382010",x"3a2211",x"38200f",x"392010",x"361f10",x"371f0f",x"341f0f",x"311c0f",x"311c10",x"362011",x"392111",x"372010",x"382011",x"3c2211",x"3c2310",x"38200f",x"392210",x"3c2410",x"39220f",x"3a220f",x"301d0c",x"2b1c0c",x"2c1b0c",x"26170b",x"2d1b0f",x"2e1c0f",x"331e0e",x"382110",x"3a2210",x"37200f",x"341e0d",x"362010",x"392110",x"311d0f",x"362011",x"362012",x"311e11",x"2c1a0f",x"2d1a0c",x"29180b",x"2d1a0c",x"321c0d",x"2e1b0c",x"361e0e",x"2f1c0f",x"382215",x"352013",x"362012",x"2c190c",x"241409",x"1e1208",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"3d230f",x"522f16",x"4a2a13",x"472812",x"452711",x"432510",x"432510",x"452712",x"422511",x"432611",x"482912",x"442611",x"3f230f",x"3b200d",x"3d210e",x"3f220f",x"3f220f",x"412410",x"3b200e",x"3f230f",x"3f230f",x"3f230f",x"3c210e",x"3d220f",x"3d220f",x"3c210e",x"3d220f",x"3e220f",x"3e220f",x"3f2310",x"3e230f",x"3c210f",x"3f230f",x"3f230f",x"3c210e",x"3d220e",x"3a1f0e",x"39200d",x"371e0d",x"381e0d",x"371d0c",x"361d0c",x"361d0c",x"361d0c",x"381e0d",x"381f0d",x"391f0e",x"391f0d",x"391f0d",x"391f0d",x"361d0d",x"361d0d",x"361d0c",x"371e0d",x"351c0c",x"2f1a0b",x"341c0c",x"371e0d",x"371e0d",x"371e0c",x"381f0d",x"361e0d",x"371d0c",x"331b0b",x"321a0b",x"381f0d",x"3c210f",x"381f0d",x"3b200e",x"3c210e",x"391f0d",x"3f2310",x"3e230f",x"381f0c",x"39200d",x"3b200d",x"391f0d",x"391f0d",x"381f0d",x"3b210e",x"3b200e",x"381f0c",x"3c210e",x"351d0d",x"3c220f",x"391f0e",x"3b210e",x"371f0d",x"381f0e",x"3c210e",x"3b200e",x"371e0d",x"351d0c",x"361d0d",x"381f0d",x"371e0d",x"3a200e",x"3a200e",x"3a200f",x"3a200e",x"3a210f",x"3a200e",x"39200e",x"3b220f",x"38200f",x"3d220f",x"39200e",x"381f0d",x"39200e",x"3a200e",x"3a210f",x"3a200e",x"3a210f",x"3d220f",x"39200e",x"361d0d",x"361d0c",x"341c0c",x"361e0d",x"39200e",x"39200e",x"361e0d",x"38200e",x"371f0e",x"311b0c",x"331c0c",x"3a210e",x"39200e",x"3a200e",x"3b200e",x"3a200e",x"3a200e",x"391f0e",x"351d0d",x"361e0d",x"3a200f",x"371f0e",x"3a200e",x"381f0e",x"351d0d",x"361e0d",x"341d0d",x"331c0c",x"331c0c",x"351d0c",x"361d0d",x"351d0d",x"371f0d",x"361e0d",x"371f0d",x"371f0d",x"341d0c",x"331c0c",x"351d0d",x"361d0d",x"341c0c",x"331c0c",x"361e0d",x"331d0c",x"3a200e",x"422511",x"371e0e",x"371e0e"),
(x"462813",x"462813",x"4b2c15",x"361f0f",x"3c2311",x"391f0d",x"28170a",x"321c0c",x"301b0c",x"2f1a0b",x"2b170a",x"301b0c",x"321d0c",x"311b0b",x"2c180a",x"2c180a",x"301a0b",x"2f1a0b",x"2e1a0b",x"2b170a",x"27160a",x"2b180a",x"2d190b",x"1a1008",x"150e07",x"150e07",x"29170a",x"251509",x"2a170a",x"29170a",x"261609",x"1d1208",x"150e07",x"150e07",x"1f1208",x"412511",x"191008",x"221409",x"2d1a0b",x"2d190b",x"311c0c",x"361f0e",x"351e0d",x"2f1b0c",x"2a180a",x"28170a",x"2f1b0c",x"301b0c",x"2d190b",x"2b180a",x"2a170a",x"301b0c",x"2a180b",x"1f1209",x"28170a",x"27160a",x"28170a",x"251509",x"201208",x"150e07",x"150e07",x"2d190b",x"211309",x"28160a",x"251509",x"231409",x"211308",x"150e07",x"150e07",x"3c210f",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"361e0d",x"331c0c",x"331c0c",x"2f1a0b",x"341d0d",x"311b0c",x"311b0c",x"301b0c",x"2d190b",x"2e1a0b",x"311c0c",x"341d0d",x"301b0c",x"341d0d",x"321c0c",x"321c0c",x"321c0c",x"321c0d",x"341d0d",x"36200e",x"371f0e",x"371e0d",x"381f0e",x"351d0c",x"371e0c",x"361d0c",x"361d0c",x"2f180a",x"231006",x"221006",x"251107",x"361d0c",x"371e0d",x"3a200e",x"3b210f",x"351d0c",x"39200e",x"3d2310",x"381f0e",x"3a200d",x"301a0a",x"361d0c",x"391f0d",x"381f0d",x"371e0c",x"311b0b",x"341c0c",x"381f0d",x"361e0d",x"381f0e",x"3a200e",x"381f0d",x"361d0d",x"321c0c",x"321b0b",x"301a0b",x"301a0b",x"2d190b",x"2e1a0b",x"2d190b",x"2f1a0c",x"311c0c",x"331d0d",x"321c0d",x"321d0d",x"301b0c",x"301b0c",x"321c0d",x"321d0d",x"331d0d",x"301b0c",x"2f1a0b",x"2f1a0b",x"321c0d",x"301b0c",x"2e1a0b",x"2d190b",x"2d190b",x"2f1a0b",x"301b0c",x"301b0c",x"2f1a0b",x"301b0b",x"321c0c",x"321b0c",x"341c0c",x"361d0d",x"381f0e",x"381f0d",x"381f0d",x"361d0c",x"371f0d",x"361d0c",x"371e0d",x"3b200e",x"3c220f",x"3d220f",x"3b200e",x"391f0d",x"381f0d",x"3b200e",x"3a200e",x"371f0d",x"361d0d",x"331c0c",x"331c0c",x"331d0d",x"2d190b",x"28170a",x"25150a",x"201309",x"1f1208",x"24150a",x"26160a",x"28170a",x"2d1a0b",x"2e1a0c",x"2e1a0b",x"2e190b",x"311c0d",x"321d0d",x"2f1c0d",x"2a180b",x"29180b",x"29170a",x"28170a",x"26160a",x"241509",x"201309",x"1d1108",x"1c1008",x"1c1008",x"1e1108",x"241509",x"28170a",x"2d190b",x"311c0c",x"321d0d",x"301b0c",x"29170a",x"2d1a0b",x"29170a",x"29170a",x"241509",x"211308",x"211308",x"201308",x"231409",x"27160a",x"221409",x"201309",x"190f07",x"502f18",x"1f1811",x"1f1811",x"1f1912",x"1f1811",x"201912",x"1f1811",x"1d1710",x"1d1710",x"1e1711",x"1b150e",x"1b150e",x"171009",x"150e07",x"23160b",x"23160b",x"28190d",x"2f1c0e",x"341e0f",x"36200f",x"351e0f",x"341d0e",x"351d0e",x"3a2110",x"3d2312",x"3e2414",x"3c2314",x"3c2211",x"402513",x"412613",x"412613",x"3f2413",x"3c2211",x"3e2412",x"3b2111",x"3c2211",x"3d2212",x"3e2412",x"3f2413",x"3c2211",x"3a2110",x"3c2211",x"3b2111",x"361f10",x"382011",x"3b2312",x"3e2512",x"3e2413",x"3f2511",x"3d2411",x"3f2512",x"412713",x"412612",x"3d2311",x"3d2312",x"3d2513",x"412714",x"432813",x"402614",x"422712",x"3f2512",x"3d2412",x"3b2212",x"3c2312",x"3c2412",x"382011",x"3c2312",x"3e2413",x"3d2413",x"402512",x"3f2614",x"402714",x"402716",x"3e2615",x"3c2615",x"3a2412",x"372212",x"3a2614",x"362212",x"2d1e12",x"2b1c11",x"291c10",x"25180f",x"2b1c12",x"331f12",x"362113",x"372213",x"3a2413",x"362112",x"392312",x"3f2816",x"3a2516",x"392416",x"382417",x"382416",x"382315",x"372416",x"372315",x"2f1f14",x"331f12",x"2f1e12",x"352013",x"331f13",x"392518",x"3a2619",x"372215",x"311f13",x"2b1b11",x"23170d",x"1c140c",x"1c140d",x"1c140d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"37200e",x"37200e",x"4b2b14",x"39200e",x"351d0d",x"311b0c",x"331d0d",x"311b0c",x"2d190b",x"2a170a",x"2c190b",x"2a180b",x"2c190b",x"2d190b",x"26160a",x"29170a",x"28160a",x"28160a",x"28160a",x"251509",x"231409",x"1f1208",x"201309",x"241409",x"251509",x"221309",x"221409",x"26150a",x"2a180a",x"27160a",x"231509",x"251509",x"241409",x"241509",x"221409",x"231409",x"1e1208",x"221409",x"221409",x"211309",x"180f07",x"221409",x"201309",x"201309",x"1c1108",x"231509",x"25150a",x"221409",x"211409",x"241509",x"28170a",x"241509",x"28170a",x"26160a",x"28170a",x"29180b",x"26160a",x"1e1208",x"211309",x"1f1208",x"211308",x"1e1108",x"1d1108",x"190f07",x"190f07",x"1a0f07",x"1f1208",x"221309",x"27160a",x"27160a",x"251509",x"28160a",x"2d1a0b",x"2a180b",x"2d190b",x"201308",x"1b1108",x"28170a",x"2b180a",x"28160a",x"2b180a",x"2a180a",x"341d0c",x"28170a",x"28170a",x"241509",x"241509",x"1c1108",x"180f07",x"170f07",x"1c1108",x"221409",x"231409",x"241509",x"26160a",x"251509",x"211409",x"211409",x"221409",x"26160a",x"211409",x"1a1008",x"27160a",x"211309",x"24150a",x"1f1309",x"241509",x"221409",x"241509",x"25160a",x"231409",x"211309",x"211309",x"241509",x"27170a",x"201309",x"231409",x"211309",x"231409",x"201208",x"211309",x"211309",x"1f1208",x"170f07",x"1b1108",x"150e07",x"1d1108",x"1c1108",x"1c1108",x"1d1108",x"1f1208",x"211409",x"231409",x"1d1108",x"221409",x"1e1208",x"180f08",x"1d1108",x"1b1108",x"1d1108",x"1f1208",x"1f1309",x"201309",x"1e1208",x"1f1208",x"221409",x"241509",x"1d1108",x"231509",x"201309",x"241509",x"241509",x"25150a",x"1f1208",x"27160a",x"201309",x"26160a",x"28170b",x"211309",x"231409",x"211309",x"2f1a0b",x"2d180b",x"2d180b"),
(x"452712",x"452712",x"492a15",x"371f0e",x"3b2210",x"472913",x"361f0e",x"331d0d",x"361f0e",x"38200f",x"351e0e",x"2a170a",x"291609",x"341d0d",x"2e1b0c",x"2f1a0b",x"2e1a0b",x"2a180a",x"2d190b",x"2f1b0c",x"2a180b",x"2f1b0c",x"1d1108",x"150e07",x"150e07",x"371e0d",x"2f1b0c",x"241509",x"271609",x"29170a",x"1e1208",x"150e07",x"150e07",x"2d1a0c",x"412511",x"180f07",x"412511",x"27160a",x"150e07",x"2a180b",x"2b190b",x"27160a",x"28160a",x"241409",x"211309",x"27160a",x"27160a",x"251509",x"29170a",x"29170a",x"261509",x"29170a",x"251509",x"27160a",x"2c190b",x"25150a",x"221309",x"221409",x"150e07",x"150e07",x"2c180a",x"2f1a0b",x"170f07",x"251509",x"251509",x"211309",x"150e07",x"150e07",x"231509",x"191008",x"26160a",x"1a1008",x"150e07",x"150e07",x"150e07",x"321c0c",x"39200e",x"351e0d",x"341c0c",x"3a200e",x"402511",x"3e230f",x"3f2410",x"3c220f",x"39200f",x"361f0e",x"301b0c",x"321c0d",x"331c0d",x"331d0d",x"321c0c",x"2f1a0b",x"2d190b",x"301b0c",x"321d0d",x"321d0d",x"2b190b",x"231509",x"25160a",x"2b190b",x"311b0c",x"2e1a0b",x"301b0c",x"361f0e",x"341e0d",x"2c190b",x"2f1b0c",x"38200f",x"39210f",x"351e0d",x"38200e",x"3a210f",x"3e2411",x"3b220f",x"381f0e",x"3c2210",x"3a210f",x"3a200e",x"3b200e",x"3a200d",x"381f0d",x"381f0e",x"3f2310",x"391f0d",x"3f2310",x"39200e",x"361e0d",x"341d0d",x"321c0c",x"321d0d",x"2d190b",x"2f1a0b",x"331b0b",x"3b210e",x"402410",x"412612",x"402511",x"3e2410",x"3c2210",x"371f0e",x"361d0d",x"381f0d",x"3a210f",x"381f0e",x"351d0d",x"381e0d",x"381f0d",x"381f0d",x"351d0d",x"341d0c",x"2f190b",x"2e190b",x"29170a",x"261509",x"27160a",x"29170a",x"2e1a0b",x"331c0d",x"311b0c",x"2d180a",x"2d190b",x"29170a",x"231409",x"381f0e",x"371e0d",x"231309",x"29170a",x"2e190b",x"2e190b",x"321c0c",x"311b0b",x"331c0c",x"361e0e",x"39200f",x"39200e",x"3a210f",x"3b220f",x"38200e",x"311b0c",x"2b190b",x"27160a",x"2c180b",x"321c0d",x"301b0c",x"2f1a0c",x"2d190b",x"2a180b",x"29170a",x"26160a",x"27170a",x"2a180b",x"2e1a0c",x"2f1b0c",x"2f1a0b",x"2f1a0b",x"2f1a0c",x"311c0d",x"311c0d",x"2f1b0c",x"2d1a0c",x"2b180b",x"2d1a0b",x"2c190b",x"29170a",x"25150a",x"25160a",x"25160a",x"25160a",x"27160a",x"2b190b",x"2e1a0c",x"301b0c",x"331d0d",x"321c0d",x"321c0d",x"2e1a0b",x"28170a",x"27160a",x"29170b",x"28170a",x"261609",x"261509",x"261609",x"251509",x"27170a",x"25150a",x"201309",x"1a1008",x"4b2d16",x"1f1811",x"1f1811",x"1e1710",x"1f1811",x"1f1812",x"1f1811",x"1f1912",x"1d1610",x"1d1710",x"1b150e",x"1b150e",x"17100a",x"150e07",x"231409",x"231409",x"29180b",x"301c0e",x"2e1a0d",x"331c0e",x"301a0b",x"321c0c",x"341d0d",x"351d0d",x"351d0e",x"3a2111",x"3a2213",x"3b2211",x"3c2211",x"3c210f",x"3e230e",x"412410",x"432711",x"381d0c",x"3e220f",x"3e220f",x"3d210e",x"3d220e",x"3b200e",x"3a1f0d",x"391e0d",x"3d2210",x"3c2110",x"3b2110",x"371f0f",x"3e2311",x"3b220f",x"422713",x"402511",x"422612",x"452813",x"452813",x"442712",x"412612",x"3d2312",x"3e2411",x"442813",x"462a14",x"422713",x"432813",x"402511",x"402611",x"3f2412",x"3b2010",x"3d2311",x"3e2412",x"3e2411",x"3e2311",x"3d2211",x"3b2010",x"3f2513",x"462c17",x"452b17",x"402918",x"432917",x"422917",x"3e2616",x"422a17",x"372314",x"3c2715",x"352214",x"372414",x"3b2616",x"3d2718",x"3c2617",x"3c2616",x"3e2715",x"422916",x"3c2515",x"412815",x"3e2714",x"372215",x"402918",x"412b1a",x"3e2718",x"3b2517",x"392416",x"342114",x"362317",x"362215",x"311f13",x"382214",x"382417",x"39271a",x"3c281b",x"3d281c",x"372214",x"28180b",x"21140b",x"1a110a",x"191109",x"191109",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38281d",x"38281d",x"3d210e",x"321c0c",x"2e190b",x"2b180a",x"27160a",x"251509",x"221309",x"201208",x"1c1108",x"1e1108",x"1f1208",x"201308",x"211409",x"201309",x"1b1108",x"1d1108",x"1e1108",x"191008",x"1b1008",x"1a1008",x"1a1008",x"1c1108",x"150e07",x"1b1008",x"150e07",x"180f07",x"1f1208",x"1c1108",x"1f1209",x"211409",x"201309",x"1d1108",x"1d1208",x"1d1108",x"1c1108",x"150e07",x"150e07",x"191008",x"150e07",x"1f1309",x"201309",x"1d1208",x"1d1108",x"170f07",x"170f07",x"170f07",x"150e07",x"1c1108",x"1e1208",x"180f07",x"1c1108",x"150e07",x"1b1108",x"211409",x"150e07",x"150e07",x"170f07",x"1b1108",x"150e07",x"150e07",x"180f07",x"1b1108",x"150e07",x"201309",x"150e07",x"1b1108",x"1c1108",x"201309",x"1c1108",x"201309",x"1c1108",x"1f1208",x"201309",x"1d1108",x"1c1108",x"1a1008",x"1d1108",x"150e07",x"856e53",x"856d51",x"94785e",x"977c5c",x"8b7358",x"8f7758",x"8e7458",x"93785d",x"937b5d",x"876f54",x"846e54",x"957a5d",x"7f694d",x"93795c",x"816d52",x"150e07",x"150e07",x"180f07",x"150e07",x"180f07",x"180f07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"180f08",x"170f07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1008",x"170f07",x"180f07",x"150e07",x"150e07",x"191008",x"191008",x"1d1108",x"1e1208",x"191008",x"321c0c",x"311c0c",x"311c0c"),
(x"422712",x"422712",x"472914",x"311b0c",x"38200f",x"3a200e",x"28160a",x"29170a",x"2d190a",x"2f1a0b",x"2d190b",x"2d190b",x"2e1b0d",x"321d0d",x"2e1a0b",x"2c190b",x"2c190b",x"2c190b",x"2a180a",x"2a180b",x"2b180b",x"28170a",x"150e07",x"150e07",x"4c2a13",x"150e07",x"422510",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"492912",x"311c0d",x"1a1008",x"150e07",x"150e07",x"26160a",x"351e0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"381f0e",x"150e07",x"2c190b",x"271609",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200d",x"211308",x"150e07",x"211409",x"1c1108",x"150e07",x"150e07",x"150e07",x"331c0c",x"2d190a",x"341c0c",x"361e0d",x"3c210f",x"412511",x"412410",x"422611",x"3b210f",x"361e0d",x"321c0c",x"311c0d",x"2e1a0b",x"311c0d",x"301b0c",x"321c0c",x"311c0c",x"321c0c",x"311b0c",x"2f1a0b",x"2e1a0b",x"2a180b",x"27170a",x"27160a",x"2d190b",x"311b0c",x"321c0d",x"331d0d",x"351d0d",x"321c0c",x"2b180a",x"2e1a0b",x"331c0c",x"321b0b",x"301a0b",x"331c0c",x"351d0c",x"381f0d",x"3c220f",x"412612",x"3d2310",x"3c220f",x"3a200e",x"391f0d",x"39200d",x"3b210f",x"3b200f",x"412511",x"452712",x"432611",x"3e230f",x"3b210f",x"39200e",x"351d0d",x"341d0d",x"2f1a0b",x"311c0c",x"361f0d",x"361d0d",x"381f0d",x"402511",x"3e2310",x"3d2310",x"3d2410",x"3d2310",x"3b2210",x"3a210f",x"371f0e",x"341d0d",x"361d0d",x"3b210f",x"3f2310",x"3e220f",x"3b210e",x"39200e",x"39200e",x"351e0d",x"2e1a0b",x"2a180a",x"28160a",x"271609",x"29170a",x"2d190b",x"2f1a0b",x"301b0b",x"2e1a0b",x"2c190b",x"251509",x"301b0c",x"351d0d",x"251509",x"29170a",x"2c180a",x"2d180a",x"2f1a0b",x"311a0b",x"321b0b",x"331c0b",x"351c0c",x"381f0d",x"39200e",x"3a200e",x"381f0d",x"311c0c",x"2c190b",x"2c190b",x"2f1a0b",x"341d0d",x"351d0d",x"361e0e",x"361f0e",x"331d0d",x"331d0d",x"311c0c",x"301b0c",x"2e1a0c",x"2f1a0c",x"311c0c",x"321c0d",x"321c0d",x"331d0d",x"2f1a0b",x"2d190b",x"2b180a",x"2d1a0b",x"301c0c",x"2f1a0b",x"2f1b0c",x"2e1a0c",x"29170a",x"27160a",x"251509",x"241509",x"251509",x"27160a",x"28160a",x"2a170a",x"2d190a",x"2e190b",x"301b0b",x"331c0c",x"351e0e",x"37200f",x"351f0e",x"301b0b",x"301b0b",x"2c190b",x"2c190b",x"29170a",x"29170b",x"251509",x"211309",x"2b190b",x"4e2d17",x"201912",x"201912",x"201a13",x"1f1812",x"1f1812",x"1f1812",x"1f1912",x"1f1912",x"1d1610",x"1d1710",x"1b150e",x"17110a",x"150e07",x"231409",x"231409",x"2a180d",x"2f1c0f",x"311d0f",x"341f10",x"361f0f",x"382010",x"38200e",x"3a200e",x"3f2512",x"412615",x"3e2615",x"3c2313",x"3c2313",x"3b2010",x"3b200d",x"3d220e",x"3b210d",x"3c210e",x"3d220e",x"3f230f",x"3f230f",x"3c200d",x"3b200d",x"391f0d",x"381e0d",x"3a200f",x"381f0f",x"371e0e",x"361e0e",x"371e0e",x"371e0e",x"381f0e",x"3a210f",x"3e220f",x"3c2210",x"3f2411",x"3f2412",x"3d2312",x"3c2212",x"3e2412",x"432713",x"432813",x"412514",x"432813",x"412613",x"402612",x"3e2313",x"3d2512",x"382010",x"3e2312",x"3d2310",x"3f2412",x"402412",x"412511",x"412614",x"422715",x"402816",x"3f2918",x"412a19",x"402919",x"422918",x"432b19",x"3e2818",x"3d281a",x"382416",x"3a2517",x"3a2719",x"3d271a",x"3a2619",x"382417",x"3b2717",x"3c2718",x"3e2717",x"3e2615",x"412a18",x"442c1a",x"442d1d",x"452e1d",x"3e2a1c",x"3a271a",x"3b271a",x"3a2719",x"372519",x"382517",x"392516",x"372316",x"392518",x"3c2a1c",x"3c291c",x"3c291d",x"39261a",x"2b1a0e",x"201309",x"190f08",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422e21",x"422e21",x"452611",x"2b180b",x"2a180b",x"231409",x"211409",x"1f1209",x"1c1108",x"191008",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"180f07",x"1d1108",x"150e07",x"170f07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"967c5d",x"8e735a",x"977d5f",x"987c5e",x"997d5e",x"987f60",x"977d5f",x"9a7e60",x"9a7e60",x"977e60",x"997e60",x"977f60",x"8b7359",x"7e664e",x"977d5d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"2e1a0c",x"2c190b",x"2c190b"),
(x"462913",x"462913",x"452813",x"341e0d",x"3c2311",x"3a200e",x"432510",x"43240f",x"43240f",x"3d1f0d",x"3d1f0c",x"43240f",x"3e1f0d",x"4b2a13",x"4b2a13",x"4b2a13",x"4a2a14",x"432611",x"442611",x"452712",x"432511",x"432611",x"3c200d",x"43240f",x"412410",x"341d0d",x"311c0c",x"422510",x"3f220f",x"311b0b",x"3f210e",x"381f0d",x"2d1a0b",x"321c0c",x"39200e",x"371e0d",x"2f1a0b",x"321b0b",x"321a0b",x"40220e",x"3f210e",x"3d200d",x"3f220e",x"412611",x"412511",x"472812",x"4a2812",x"492912",x"462611",x"4c2a13",x"4a2913",x"4f2d15",x"4d2c15",x"4e2d14",x"472812",x"452611",x"422511",x"412410",x"432510",x"371f0e",x"341d0d",x"2a180a",x"341c0c",x"422510",x"2b180b",x"3c210e",x"301b0c",x"311b0c",x"351d0d",x"311b0c",x"2a180b",x"1f1208",x"150e07",x"150e07",x"150e07",x"4a2b15",x"351e0b",x"351d0e",x"371f0f",x"3d2312",x"422713",x"422613",x"3f2514",x"3b2313",x"372112",x"331f12",x"331f11",x"321f11",x"321f11",x"2f1c10",x"331f10",x"341f10",x"311c0e",x"321c0e",x"331d0f",x"331d0e",x"321c0d",x"331d0d",x"301b0c",x"311b0c",x"2f1a0b",x"311b0c",x"311b0c",x"341d0c",x"351e0d",x"321b0c",x"361e0d",x"3b210e",x"381f0d",x"331c0c",x"2f190b",x"2f190b",x"30190a",x"31190a",x"30190a",x"351d0d",x"3c230f",x"3b210f",x"3c220f",x"3e2410",x"3c220f",x"3e230f",x"412511",x"432611",x"3b200e",x"381d0c",x"391f0d",x"3c220f",x"3c220f",x"3b210f",x"3a200e",x"361d0c",x"341c0c",x"381f0d",x"3b200f",x"3d220f",x"3c220f",x"3a200e",x"341c0c",x"331b0c",x"2e170a",x"311a0b",x"321b0b",x"2f190b",x"311a0b",x"3b220f",x"3f2411",x"412511",x"3a200e",x"39200e",x"371e0d",x"371e0d",x"361e0e",x"321c0d",x"2e1b0c",x"2b190b",x"2c190b",x"301c0c",x"311b0c",x"331d0d",x"321c0c",x"2f1a0b",x"2a180b",x"29170a",x"361e0d",x"2f1a0c",x"2f1a0b",x"341d0c",x"351d0d",x"39200e",x"3a200e",x"3a200e",x"38200e",x"381f0d",x"3a200e",x"3b210f",x"3a200e",x"39200e",x"2e1a0b",x"2c180b",x"2d190b",x"2e1a0b",x"321c0c",x"341d0d",x"351e0d",x"341d0d",x"361f0e",x"331d0d",x"331d0d",x"321c0d",x"311b0c",x"2d190b",x"321c0c",x"331d0d",x"321c0c",x"331c0c",x"321c0c",x"2f1a0c",x"311c0c",x"341d0d",x"301b0c",x"321c0c",x"2f1a0b",x"2e1a0b",x"2f1a0b",x"2a180a",x"2a190c",x"2a190c",x"29180c",x"2e1c0f",x"301d0f",x"301d11",x"321e11",x"311d11",x"2f1d11",x"2f1c12",x"311e11",x"2f1d11",x"382214",x"382214",x"352012",x"342012",x"331f12",x"301d0f",x"342011",x"2b1a0d",x"27180c",x"301a0b",x"512f19",x"201a13",x"201a13",x"201a13",x"211a13",x"211a14",x"1f1812",x"1e1811",x"1f1812",x"1d1711",x"1d1610",x"1b140e",x"171009",x"150e07",x"201309",x"201309",x"25160b",x"2c1a10",x"2f1e12",x"382213",x"3a2415",x"3a2212",x"3b2212",x"3b2110",x"3e2412",x"3d2514",x"402715",x"412716",x"432918",x"422813",x"442812",x"3e230f",x"3d210f",x"402410",x"412411",x"40230f",x"412410",x"402310",x"3e220f",x"3c210e",x"412512",x"3f2311",x"3d2110",x"3f2411",x"3f2512",x"3c2312",x"3c2212",x"3a2111",x"3b2211",x"3b2211",x"3d2311",x"402512",x"3e2412",x"3b2211",x"3b2111",x"3d2312",x"3e2513",x"3f2614",x"422714",x"432815",x"412714",x"402614",x"3d2412",x"3d2412",x"3b2211",x"3b2111",x"3b2111",x"412613",x"412514",x"3f2312",x"432916",x"442a17",x"432b18",x"422a19",x"462c1c",x"412919",x"422b1b",x"41291a",x"3f2919",x"3a2618",x"372518",x"3d281a",x"3b2719",x"3e291a",x"3f291b",x"3e281a",x"3d281b",x"3d281a",x"3b2719",x"392519",x"3d2719",x"3c2a1d",x"422d1d",x"462f1f",x"3e2a1d",x"3f2b1d",x"3b291c",x"3a281b",x"3d2a1d",x"3c291c",x"3a261a",x"342318",x"35251a",x"3a291d",x"3e2c1f",x"3d2b1f",x"372619",x"2a1b10",x"1d1108",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"433328",x"433328",x"472912",x"2c1a0b",x"24150a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"8e755a",x"947b5c",x"937a5d",x"997e60",x"997e60",x"9a7e60",x"947a5e",x"967c5e",x"997e60",x"987d5f",x"957c5d",x"967c5e",x"947a5e",x"947b5e",x"977a5e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1a0b",x"2a180b",x"2a180b"),
(x"442712",x"442712",x"432611",x"331d0d",x"3d2411",x"381f0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442712",x"221409",x"2f1b0c",x"341d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"422410",x"301a0c",x"25150a",x"241509",x"2a180a",x"2e1a0c",x"29180b",x"231509",x"150e07",x"150e07",x"3f2410",x"27170a",x"150e07",x"150e07",x"150e07",x"311c0c",x"27160a",x"351e0d",x"231509",x"231409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"361e0d",x"3c220f",x"150e07",x"351f0e",x"39200e",x"351e0d",x"321d0d",x"311b0c",x"2f1b0b",x"39200f",x"3c210f",x"371f0e",x"150e07",x"2d1a0c",x"241509",x"150e07",x"150e07",x"150e07",x"4a2b15",x"38200e",x"361e0e",x"3e2311",x"412614",x"412513",x"422615",x"3a2213",x"331f12",x"301d12",x"301e12",x"2f1e12",x"311e12",x"342013",x"2f1d11",x"2e1c10",x"2f1c0f",x"321e10",x"321d0e",x"311c0e",x"2f1b0d",x"2e1a0b",x"2e190b",x"2e1a0b",x"2f1a0b",x"311b0c",x"331d0d",x"351e0d",x"341d0d",x"351d0d",x"361e0d",x"371e0d",x"3a200e",x"381f0e",x"341d0e",x"341d0e",x"392010",x"392010",x"39200f",x"371e0f",x"392010",x"3a2010",x"3b2211",x"3f2413",x"412714",x"422814",x"402614",x"422713",x"432713",x"422613",x"3e2312",x"3a2111",x"3a2111",x"39200f",x"3b2110",x"3d2311",x"3c2110",x"3c2110",x"3e2411",x"412613",x"422713",x"412613",x"412613",x"3e2411",x"3b2211",x"3b2211",x"3c2312",x"3b2211",x"351e0f",x"321c0d",x"351f0f",x"3b2211",x"3d2311",x"3a210e",x"39200e",x"39210f",x"371f0e",x"38200e",x"351f0e",x"301c0d",x"2d1a0c",x"2f1b0c",x"321d0d",x"351f0e",x"341e0d",x"331d0d",x"2f1b0c",x"2b190b",x"311c0c",x"3b210f",x"26160a",x"2c190b",x"301b0c",x"351e0d",x"371f0e",x"38200f",x"39200f",x"39200f",x"39200e",x"39200e",x"39200e",x"371f0d",x"351e0d",x"301a0c",x"2a170a",x"2e1a0b",x"311c0c",x"321c0c",x"341d0d",x"321b0c",x"2d180a",x"2b170a",x"2c180a",x"2d190b",x"2c180b",x"2f1a0c",x"2d190b",x"2b180a",x"2d190b",x"301b0c",x"311c0c",x"2f1b0c",x"2c190b",x"2a170a",x"2b180a",x"2c180b",x"2d1a0b",x"2f1a0b",x"2e1a0c",x"2c1a0d",x"29190f",x"2a1b10",x"2b1c11",x"2c1e14",x"2f1f15",x"312014",x"342217",x"362317",x"382518",x"392418",x"382519",x"382518",x"382517",x"392619",x"382519",x"342316",x"352316",x"352418",x"322114",x"302116",x"2c1e14",x"261a11",x"24180f",x"4e2e18",x"201a13",x"201a13",x"201a13",x"201a13",x"201a13",x"211a14",x"1f1912",x"1f1811",x"1d1710",x"1d160f",x"1b150e",x"171009",x"150e07",x"221409",x"221409",x"2c1c10",x"332114",x"342114",x"372316",x"392315",x"3a2414",x"392313",x"3d2413",x"3f2715",x"3f2615",x"432a19",x"432a18",x"412916",x"432915",x"432815",x"432813",x"432712",x"422611",x"412410",x"422510",x"402310",x"452712",x"432713",x"442813",x"452814",x"432713",x"432714",x"442814",x"422715",x"412715",x"402615",x"412615",x"3f2514",x"3e2513",x"3f2514",x"3e2616",x"3e2515",x"3a2214",x"3f2514",x"402716",x"432815",x"412715",x"402715",x"3d2515",x"371f12",x"362010",x"372111",x"392112",x"392213",x"3d2413",x"382112",x"3b2213",x"3d2313",x"422916",x"432917",x"422817",x"402817",x"412919",x"442c1b",x"462d1c",x"412b1c",x"422b1c",x"402a1a",x"3b271a",x"3b271a",x"3e291b",x"3e291c",x"3d291c",x"422c1e",x"3f291c",x"412a1c",x"452e1e",x"412b1b",x"412a1b",x"462e1e",x"432d1f",x"442f21",x"432e20",x"402b1d",x"422d1f",x"3e2a1d",x"3d2b1e",x"3b291c",x"3a2a1e",x"3a281c",x"39281c",x"37261b",x"3a2a1e",x"3b2b1f",x"3b2a1f",x"37271d",x"2c1d13",x"1d1108",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"46382d",x"46382d",x"432511",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1107",x"180f07",x"181007",x"181007",x"191007",x"1a1107",x"191007",x"8d7357",x"94795d",x"967d5e",x"947a5d",x"957c5d",x"977e5f",x"967c5f",x"977a5d",x"957b5b",x"957b5e",x"997e60",x"997e60",x"8c7255",x"8a7156",x"8a6f55",x"1a1107",x"1a1107",x"191007",x"170f07",x"160f07",x"181007",x"191007",x"191007",x"191007",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"231509",x"231509"),
(x"452712",x"452712",x"432611",x"311c0d",x"3a210f",x"472813",x"211409",x"311d0d",x"2d1b0c",x"311c0d",x"2e1a0b",x"29170a",x"2d1a0b",x"27170a",x"29180b",x"28170a",x"1c1108",x"150e07",x"150e07",x"150e07",x"391f0e",x"150e07",x"26160a",x"251509",x"1f1208",x"150e07",x"150e07",x"150e07",x"402310",x"2d190b",x"241509",x"1b1108",x"150e07",x"150e07",x"341d0d",x"381f0e",x"170f07",x"231509",x"2a190b",x"26170a",x"150e07",x"150e07",x"402410",x"2f1b0c",x"3d2411",x"150e07",x"211409",x"37210f",x"150e07",x"1c1208",x"26160a",x"27170a",x"2c190b",x"21150a",x"29180b",x"24150a",x"150e07",x"150e07",x"150e07",x"150e07",x"452812",x"150e07",x"402511",x"3a210f",x"341d0d",x"321d0e",x"150e07",x"25160a",x"28170b",x"150e07",x"2b180b",x"1d1108",x"150e07",x"150e07",x"150e07",x"422613",x"331f12",x"392313",x"3d2516",x"3e2516",x"3c2516",x"3c2517",x"342114",x"2f1f14",x"291c13",x"211811",x"201710",x"1f170f",x"201810",x"1f160f",x"21170e",x"27190e",x"2e1c0f",x"301c0e",x"311c0e",x"321d0e",x"321c0c",x"331d0d",x"311c0c",x"321c0c",x"321c0c",x"321c0d",x"351e0d",x"38200f",x"371f0e",x"371f0f",x"3b2212",x"412715",x"412715",x"3f2717",x"3e2717",x"402818",x"3e2818",x"3d2617",x"402819",x"412a19",x"422a1a",x"3f2818",x"3a2518",x"362317",x"342217",x"362316",x"3d2617",x"412819",x"422918",x"3f2617",x"3c2517",x"3b2517",x"3b2415",x"3c2516",x"3c2617",x"3a2415",x"382214",x"382215",x"3a2314",x"3d2415",x"3e2616",x"3e2514",x"3d2515",x"382213",x"372215",x"362113",x"352112",x"311f12",x"271a0f",x"1c140d",x"19120c",x"1a130c",x"1c120a",x"25180c",x"311d0d",x"37210f",x"35210f",x"351f0e",x"2f1b0c",x"2a190b",x"2a190b",x"301c0d",x"361f0f",x"36200e",x"331d0d",x"2e1a0c",x"26160a",x"1b1108",x"3a210f",x"1b1108",x"24150a",x"2e1b0c",x"331e0e",x"361f0e",x"37200f",x"37200f",x"371f0e",x"361f0e",x"341d0d",x"341d0d",x"341d0d",x"341c0d",x"311c0c",x"2d190b",x"2a180b",x"2a170a",x"2c180b",x"301b0c",x"2f1a0b",x"301b0b",x"301b0b",x"311c0c",x"301b0c",x"2e1a0b",x"2d190b",x"2c190b",x"2d1a0b",x"2f1a0c",x"301b0c",x"301b0c",x"2d1a0b",x"2c190b",x"2a180b",x"2b190b",x"2c190b",x"2e1a0b",x"2f1b0c",x"2d1a0b",x"2c1a0d",x"2b1b0f",x"2b1c11",x"2c1d11",x"2d1e14",x"302116",x"352418",x"382619",x"3b2719",x"3d291a",x"3c281b",x"372317",x"3a2619",x"3c2719",x"3c2718",x"3b271a",x"382619",x"332116",x"322217",x"2f1f15",x"302016",x"2b1d13",x"251a11",x"1f160f",x"4d2e18",x"201a14",x"201a14",x"201a13",x"201a13",x"201912",x"211a14",x"1e1710",x"1f1811",x"1f1812",x"1d160f",x"1b140d",x"17110a",x"150e07",x"201208",x"201309",x"2a1c11",x"312013",x"362416",x"3a2517",x"3b2618",x"3b2718",x"372415",x"382314",x"3c2615",x"402a17",x"3d2817",x"3e2716",x"412817",x"3f2615",x"3c2615",x"3c2312",x"412713",x"432712",x"412511",x"3f2410",x"3f2410",x"452814",x"452814",x"462a15",x"462b16",x"452a16",x"482c17",x"462b17",x"462b18",x"442a17",x"442a18",x"452b18",x"3f2717",x"3f2816",x"412916",x"3f2716",x"3f2616",x"3f2717",x"402817",x"3d2616",x"402817",x"422a16",x"3d2515",x"3d2515",x"3f2714",x"3b2515",x"3d2414",x"3e2513",x"3d2516",x"402615",x"402615",x"422815",x"452916",x"452b17",x"462b19",x"452c1b",x"472d1a",x"442919",x"482f1d",x"442c1c",x"462d1b",x"442d1c",x"412a1b",x"402c1d",x"3f2a1a",x"3f2a1d",x"402a1c",x"402a1c",x"442d1d",x"432d1d",x"472f1f",x"4a311f",x"472f1e",x"412c1e",x"453020",x"452f1f",x"462f1f",x"463121",x"432e1f",x"3f2c1e",x"39291e",x"3a291d",x"38291e",x"39281c",x"38291d",x"36261a",x"34261c",x"382a1f",x"3b2a1d",x"382a20",x"35271d",x"291d13",x"1b1008",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d3228",x"3d3228",x"432611",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191007",x"1e1308",x"1a1107",x"1b1108",x"1b1108",x"1d1308",x"1e1308",x"1d1308",x"1a1107",x"1c1208",x"1c1208",x"1c1208",x"1b1108",x"1c1208",x"1e1308",x"221508",x"201508",x"1f1408",x"211508",x"221508",x"211508",x"241708",x"211508",x"1e1308",x"1f1408",x"1d1308",x"191107",x"180f07",x"1c1208",x"1d1308",x"1c1208",x"1c1208",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"2d1a0b",x"2d1a0b"),
(x"432712",x"432712",x"442712",x"351f0e",x"3c2210",x"3d220e",x"28170a",x"311c0c",x"2d1a0b",x"301c0c",x"311b0c",x"2f1a0b",x"311b0c",x"331d0d",x"2c190b",x"2d1a0b",x"28170a",x"221409",x"150e07",x"3c210f",x"2a180b",x"201309",x"2d1a0b",x"2b180b",x"27160a",x"241509",x"180f07",x"150e07",x"150e07",x"432511",x"371f0d",x"2a180b",x"150e07",x"311c0d",x"3b210e",x"1e1208",x"2f1b0c",x"2a180b",x"28160a",x"2c180b",x"29170a",x"150e07",x"190f07",x"201108",x"2f1a0b",x"371f0e",x"150e07",x"150e07",x"4b2a13",x"2f1a0b",x"150e07",x"2d1a0c",x"2e1b0c",x"2c1a0b",x"331d0d",x"311c0d",x"331d0d",x"27170b",x"23150a",x"150e07",x"150e07",x"452812",x"150e07",x"29180b",x"3f2410",x"2f1b0c",x"472813",x"311c0d",x"27170a",x"150e07",x"2b190b",x"1f1309",x"150e07",x"150e07",x"150e07",x"402613",x"332011",x"382415",x"3d2616",x"442a18",x"412817",x"412919",x"392516",x"312015",x"2a1e14",x"221912",x"1d160f",x"1c160f",x"1d1710",x"1b150e",x"1b150e",x"1c140c",x"25180e",x"2b1a0c",x"301c0e",x"321c0e",x"321c0c",x"301b0b",x"2f1b0c",x"29170a",x"28170b",x"29180b",x"261609",x"2a180a",x"351f0d",x"402411",x"3d2312",x"3e2312",x"3e2514",x"392313",x"3b2515",x"3a2415",x"422a19",x"432a18",x"3d2617",x"402819",x"422919",x"402919",x"3f2819",x"3b2518",x"3a2518",x"3d2819",x"432918",x"472d1a",x"492d1a",x"482c1a",x"462a19",x"442b1a",x"402718",x"3f2516",x"3e2516",x"432817",x"422816",x"442a18",x"452b18",x"392214",x"392314",x"352113",x"352113",x"322012",x"2d1d12",x"2d1c12",x"2d1d12",x"2a1a10",x"1e150e",x"1c150e",x"19130c",x"19130c",x"191109",x"21150a",x"2d190b",x"331c0c",x"371f0e",x"361f0e",x"301c0c",x"2c190b",x"2d1a0c",x"2f1c0c",x"331d0d",x"351e0e",x"341e0e",x"2e1b0c",x"25160a",x"1a1008",x"381e0d",x"191008",x"211309",x"2b190b",x"311c0d",x"331d0d",x"351e0d",x"351f0e",x"351d0d",x"341d0d",x"331c0c",x"361f0e",x"351e0d",x"341d0d",x"311b0c",x"2c180b",x"2a180b",x"2b180b",x"2c190b",x"2b170a",x"2e1a0b",x"2f1a0b",x"311b0c",x"321c0d",x"301b0c",x"2d190b",x"2b190b",x"2b190b",x"2b190b",x"2e1a0c",x"2e1a0c",x"2e1a0b",x"2d190b",x"2c190b",x"29180b",x"2a180b",x"2c190b",x"2e1a0b",x"2e1a0c",x"2e1a0c",x"2b190d",x"2a1a0f",x"2b1c10",x"2c1d11",x"2f2015",x"322216",x"342317",x"382518",x"382518",x"3b2719",x"3a2618",x"3d281b",x"3a2719",x"372518",x"392518",x"382619",x"342318",x"322217",x"312116",x"2d1e14",x"2c1e15",x"281c12",x"231911",x"1f150e",x"513018",x"201a13",x"201a13",x"201913",x"201912",x"201913",x"201a13",x"1e1711",x"1e1711",x"1f1912",x"1d160f",x"1b140d",x"171009",x"150e07",x"1e130a",x"1d130a",x"25180f",x"2c1e14",x"2f2116",x"2d1f15",x"332317",x"382517",x"372315",x"342115",x"3c2515",x"402917",x"422a17",x"3f2716",x"3e2717",x"3d2616",x"3d2514",x"3d2514",x"3b2412",x"3f2614",x"422614",x"422614",x"422713",x"412613",x"412814",x"422716",x"482b18",x"462b18",x"462c1a",x"472c1a",x"422918",x"422a18",x"412919",x"432c19",x"402918",x"432b18",x"432a19",x"442b1a",x"402918",x"422917",x"3f2818",x"412917",x"432a19",x"412918",x"432a19",x"412917",x"442a17",x"402817",x"412715",x"3e2515",x"3f2615",x"3f2717",x"3f2715",x"412816",x"432917",x"412818",x"442a1a",x"462d1b",x"462c1b",x"462d1b",x"472e1d",x"472f1d",x"472e1c",x"452d1d",x"432d1c",x"3b281b",x"39281c",x"3e291a",x"422c1e",x"412c1e",x"402a1c",x"412c1e",x"45301f",x"422c1d",x"412c1c",x"432d1d",x"472f1e",x"432e1f",x"432e20",x"412d20",x"3f2c1e",x"3e2c1e",x"3c2b20",x"3a2b20",x"3b2b20",x"3a2a1e",x"37291e",x"392a20",x"34281e",x"372a1f",x"3d2d20",x"392c21",x"35271c",x"281d15",x"1c120a",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2e25",x"3d2e25",x"331a0a",x"2f1a0b",x"351c0c",x"381f0d",x"3f230f",x"3d220f",x"3d220f",x"3a200e",x"3b200e",x"3a210f",x"38200e",x"3c220f",x"361f0d",x"3c220f",x"3c2310",x"3e2310",x"402511",x"3b2210",x"3f2411",x"3f2411",x"39210f",x"3c220f",x"3e2310",x"3c2210",x"3d2310",x"3f2410",x"402511",x"432711",x"432612",x"3f2410",x"3f2410",x"3d230f",x"3f2410",x"3b200e",x"381f0e",x"281509",x"221308",x"3b210e",x"3f230f",x"3c220f",x"371f0d",x"381f0e",x"301b0b",x"241409",x"261509",x"261509",x"29170a",x"251509",x"2b180a",x"241509",x"2f1a0b",x"3b200e",x"3b210e",x"3a200e",x"3a1f0e",x"351d0d",x"39200e",x"221409",x"2c190b",x"231409",x"29170a",x"231409",x"2b190a",x"3a200e",x"3a200e",x"3d230f",x"402410",x"3f2310",x"3d220f",x"442712",x"432611",x"442711",x"412610",x"432710",x"41250f",x"442711",x"40240f",x"422510",x"3d220e",x"3d220e",x"3f230e",x"432610",x"3c220e",x"3f250f",x"3d220e",x"432710",x"3f240e",x"40250f",x"3e240e",x"412610",x"432711",x"41250f",x"422610",x"432711",x"432712",x"402510",x"402510",x"3e2410",x"432712",x"3b220e",x"3f2410",x"341c0b",x"381f0e",x"3b220f",x"3e2310",x"3a200e",x"3e2411",x"422612",x"422612",x"3d2310",x"3f2411",x"3e2410",x"3c2310",x"3d2310",x"3e2310",x"3e2411",x"3f2411",x"412611",x"412511",x"422611",x"432712",x"412611",x"402511",x"3f2410",x"402511",x"412512",x"422612",x"422612",x"422612",x"412611",x"3f2511",x"3d2310",x"3a210f",x"402411",x"452813",x"402511",x"3d2310",x"3d2310",x"3e2410",x"3d2310",x"3c220f",x"39200f",x"3a200e",x"39200e",x"381f0f",x"361f0d",x"361e0d",x"371e0e",x"3b210f",x"3a200e",x"3d220f",x"3f2410",x"402411",x"3e2310",x"402511",x"402510",x"3f2411",x"341d0d",x"2c190b",x"251509",x"361e0d",x"361e0d"),
(x"422712",x"422712",x"462813",x"311c0d",x"3d2310",x"452812",x"29180b",x"281609",x"2f1a0b",x"2f1a0b",x"2b180a",x"2e1a0b",x"2a170a",x"2e1a0b",x"2a170a",x"281609",x"241409",x"1d1108",x"150e07",x"150e07",x"2b180a",x"29170a",x"231308",x"1d0f07",x"1d0f07",x"1f1208",x"1b1008",x"150e07",x"150e07",x"1e1108",x"3f210e",x"2b170a",x"150e07",x"442610",x"331c0c",x"27160a",x"2a180a",x"2e1a0b",x"321c0c",x"2f1b0c",x"2e190b",x"2b180a",x"180f08",x"150e07",x"150e07",x"1f1209",x"4b2b14",x"150e07",x"150e07",x"28170a",x"422410",x"211309",x"26160a",x"2e1a0b",x"2f1b0c",x"2e1b0c",x"2d1a0b",x"311c0d",x"2c1a0c",x"2a190b",x"150e07",x"150e07",x"37200f",x"2c1a0b",x"150e07",x"371f0e",x"29170b",x"26160a",x"311d0d",x"150e07",x"29180b",x"211409",x"150e07",x"150e07",x"150e07",x"452914",x"402613",x"342213",x"3a2415",x"3b2516",x"3e2718",x"3d2617",x"382316",x"311f14",x"2a1c13",x"241a12",x"1d1610",x"1c160f",x"1d1710",x"1b150e",x"1b140d",x"1c140d",x"1f150d",x"26180e",x"2b190c",x"2d1a0c",x"2d190b",x"2d190b",x"2b180b",x"29170a",x"26160a",x"25150a",x"27160a",x"2b190b",x"2f1b0c",x"341e0f",x"341e0f",x"362011",x"352013",x"2d1d11",x"2d1e13",x"311f13",x"352216",x"352215",x"352316",x"352317",x"342217",x"322116",x"2d1f15",x"2b2017",x"2a1e15",x"2d1f15",x"342115",x"392315",x"3a2417",x"311e14",x"2a1b12",x"352115",x"321f14",x"362013",x"352013",x"341f12",x"362014",x"362114",x"322014",x"342114",x"342013",x"342012",x"321f11",x"301f13",x"2f1f12",x"2f1e12",x"2f1e12",x"2a1b10",x"25180f",x"22170f",x"19120b",x"19120b",x"25170b",x"311d0e",x"3b220f",x"3c220f",x"331c0c",x"2e190b",x"2b180b",x"28170a",x"2c190b",x"311c0d",x"321c0d",x"341d0d",x"331e0e",x"2c1a0c",x"201409",x"1b1108",x"361d0d",x"2b1c11",x"2b1c11",x"2c1d12",x"2d1e13",x"302014",x"322115",x"342215",x"332114",x"332014",x"311f14",x"312014",x"352215",x"382113",x"392214",x"3b2415",x"372213",x"311f13",x"2b1c11",x"281b11",x"281b11",x"2a1b12",x"2d1d12",x"2d1b10",x"2f1c0f",x"341f11",x"392112",x"3a2111",x"3a2111",x"371f10",x"311c0f",x"29190e",x"20150d",x"1a120b",x"19120c",x"19120b",x"19130c",x"1a140c",x"1f150c",x"26180e",x"2c1c11",x"301d11",x"2f1d12",x"311f14",x"311f12",x"301f14",x"342216",x"342216",x"352317",x"362418",x"342218",x"332117",x"362317",x"392416",x"3c2517",x"3b2416",x"392315",x"382315",x"321f12",x"2e1c11",x"2a190f",x"26180e",x"24180f",x"1e140d",x"432713",x"211a13",x"211a13",x"201a13",x"201913",x"211a14",x"201a13",x"201913",x"1e1711",x"1f1811",x"1d160f",x"1b140d",x"171009",x"150e07",x"1f140a",x"20140a",x"2b1d11",x"2c1e14",x"312216",x"362517",x"382516",x"3b2718",x"402a17",x"3e2817",x"3d2617",x"432b18",x"422a17",x"3c2616",x"382214",x"3b2415",x"3b2314",x"3d2515",x"3f2714",x"3f2514",x"432815",x"442815",x"462a15",x"442915",x"452a16",x"462a18",x"482d17",x"462c18",x"472b18",x"462a17",x"472b1a",x"442a19",x"3e2717",x"412a19",x"442b19",x"3f2717",x"452c1a",x"452d1c",x"462c19",x"452b19",x"432a19",x"432a19",x"3f2817",x"432b19",x"412a1a",x"402817",x"412916",x"3d2414",x"3e2615",x"432a17",x"3e2515",x"3b2414",x"3e2516",x"3e2616",x"3d2515",x"3e2717",x"41291a",x"402918",x"422a1a",x"402a1b",x"432c1c",x"442b1c",x"422a1b",x"442c1b",x"452d1d",x"422b1c",x"422c1d",x"412c1d",x"442e1f",x"412b1c",x"432d1e",x"442d1d",x"402b1c",x"452e1f",x"452e1f",x"422c1e",x"452f1f",x"422e20",x"422e20",x"3f2c1f",x"3d2b1f",x"3c2a1f",x"392a1f",x"38291d",x"36271d",x"35271c",x"39281d",x"36291f",x"30251b",x"31281f",x"382a1e",x"34271e",x"37291e",x"291f18",x"1a110a",x"160e07",x"160e07",x"452e1e",x"452f20",x"442f21",x"3f2b1f",x"412d20",x"433022",x"422e21",x"412e20",x"3f2e21",x"3b2d20",x"3c2c20",x"3b2b1e",x"392a1e",x"37291f",x"36291f",x"35291f",x"32281d",x"30271d",x"372a1f",x"35291f",x"35291f",x"36291d",x"2c2118",x"1e150d",x"170f07",x"3c2310",x"3e2310",x"402511",x"3b2210",x"3f2411",x"3f2411",x"39210f",x"3c220f",x"3e2310",x"3c2210",x"3d2310",x"3f2410",x"402511",x"432711",x"432612",x"3f2410",x"3f2410",x"3d230f",x"3f2410",x"3b200e",x"381f0e",x"281509",x"221308",x"3b210e",x"3f230f",x"3c220f",x"371f0d",x"381f0e",x"301b0b",x"241409",x"261509",x"261509",x"29170a",x"251509",x"2b180a",x"241509",x"2f1a0b",x"3b200e",x"3b210e",x"3a200e",x"3a1f0e",x"351d0d",x"39200e",x"221409",x"2c190b",x"231409",x"29170a",x"231409",x"2b190a",x"3a200e",x"3a200e",x"3d230f",x"402410",x"3f2310",x"3d220f",x"442712",x"432611",x"442711",x"412610",x"432710",x"41250f",x"442711",x"40240f",x"422510",x"3d220e",x"3d220e",x"3f230e",x"432610",x"3c220e",x"3f250f",x"3d220e",x"432710",x"3f240e",x"40250f",x"3e240e",x"412610",x"432711",x"41250f",x"422610",x"432711",x"432712",x"402510",x"402510",x"3e2410",x"432712",x"3b220e",x"3f2410",x"341c0b",x"381f0e",x"3b220f",x"3e2310",x"3a200e",x"3e2411",x"422612",x"422612",x"3d2310",x"3f2411",x"3e2410",x"3c2310",x"3d2310",x"3e2310",x"3e2411",x"3f2411",x"412611",x"412511",x"422611",x"432712",x"412611",x"402511",x"3f2410",x"402511",x"412512",x"422612",x"422612",x"422612",x"412611",x"3f2511",x"3d2310",x"3a210f",x"402411",x"452813",x"402511",x"3d2310",x"3d2310",x"3e2410",x"3d2310",x"3c220f",x"39200f",x"3a200e",x"39200e",x"381f0f",x"361f0d",x"361e0d",x"371e0e",x"3b210f",x"3a200e",x"3d220f",x"3f2410",x"402411",x"3e2310",x"402511",x"402510",x"3f2411",x"341d0d",x"2c190b",x"251509",x"361e0d",x"000000"),
(x"442712",x"442712",x"452712",x"341e0d",x"3b2210",x"452712",x"1e1208",x"2a180a",x"2e1a0b",x"2e1a0b",x"29170a",x"281609",x"221409",x"1f1208",x"29170a",x"28170a",x"241509",x"150e07",x"150e07",x"27160a",x"331d0d",x"26160a",x"2a180a",x"211309",x"231409",x"150e07",x"150e07",x"150e07",x"371f0d",x"150e07",x"150e07",x"3f230f",x"150e07",x"3e220f",x"2d190b",x"301b0c",x"2d1a0b",x"301b0c",x"2d1a0b",x"2f1b0c",x"341e0d",x"321d0d",x"311c0c",x"28170a",x"1d1208",x"150e07",x"381f0e",x"311c0d",x"191008",x"150e07",x"150e07",x"4c2913",x"29170a",x"211409",x"331d0d",x"341e0e",x"2f1c0d",x"2f1b0c",x"2c190b",x"2a180b",x"180f07",x"150e07",x"38200e",x"150e07",x"361e0d",x"150e07",x"331d0d",x"1d1108",x"2c190b",x"150e07",x"26160a",x"1e1209",x"150e07",x"150e07",x"150e07",x"3e2413",x"301f13",x"241409",x"231409",x"241409",x"29170a",x"2e1a0b",x"301a0b",x"2e1a0b",x"2d190b",x"2b180a",x"2a170a",x"29170a",x"28170a",x"271609",x"261509",x"241509",x"211309",x"201208",x"201309",x"201309",x"1a1008",x"170f07",x"1b1108",x"1d1108",x"1c1108",x"1b1108",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"201309",x"1e1209",x"231409",x"28160a",x"2e1a0b",x"321c0c",x"2e190b",x"291609",x"2a170a",x"2e190b",x"2e1a0b",x"2c190b",x"2a180a",x"301b0c",x"331d0d",x"331d0d",x"341d0d",x"361e0d",x"341e0d",x"311b0c",x"2d190b",x"2c190a",x"2e1a0b",x"2f1a0b",x"301b0c",x"311c0c",x"321d0d",x"321c0c",x"311c0c",x"2d190b",x"2d190b",x"311b0c",x"331c0c",x"331d0d",x"341d0d",x"351e0d",x"371f0e",x"39200f",x"361f0e",x"2f1b0c",x"28170a",x"28170a",x"27160a",x"221409",x"1f1309",x"1f1309",x"231509",x"27160a",x"2a170a",x"2b180b",x"2c190b",x"2b190b",x"2b190b",x"351f0e",x"311c0d",x"28180b",x"1d1208",x"1a1008",x"2f1e13",x"2f1f13",x"311e12",x"322013",x"342015",x"362214",x"372315",x"372315",x"372215",x"342114",x"332014",x"332115",x"372214",x"3b2415",x"3d2415",x"3c2414",x"372214",x"321e12",x"2c1c11",x"291b11",x"291c11",x"2c1d12",x"2e1e12",x"2f1c11",x"311e11",x"352012",x"382112",x"382010",x"3a2011",x"371f10",x"311d0f",x"29190e",x"1f150d",x"1a120b",x"19130c",x"19130c",x"19130c",x"1b130b",x"21160c",x"28190e",x"2f1d11",x"301d11",x"311f12",x"352013",x"372215",x"372416",x"382517",x"382418",x"3b2619",x"3d2719",x"3e2819",x"382417",x"382317",x"3c2517",x"412818",x"412818",x"3f2616",x"402817",x"3c2516",x"3a2415",x"341f11",x"2e1d11",x"281a10",x"1f150d",x"432612",x"201a13",x"201a13",x"201a13",x"211a14",x"201912",x"211b14",x"201912",x"1e1710",x"1f1912",x"1c160f",x"1b150e",x"17110a",x"150e07",x"20140a",x"20140b",x"271b11",x"2e1f15",x"322317",x"372517",x"372517",x"3b2617",x"3e2817",x"3c2617",x"412919",x"492d1a",x"442b18",x"402817",x"3b2515",x"3c2415",x"3d2515",x"3f2715",x"412716",x"402816",x"3f2513",x"3f2512",x"432815",x"412714",x"432816",x"432817",x"412817",x"422917",x"452917",x"442b17",x"432a18",x"412818",x"412918",x"412817",x"422918",x"422a19",x"3f2718",x"3f2819",x"412919",x"422919",x"412919",x"3d2719",x"3d2718",x"3e2819",x"3e2716",x"3b2517",x"3d2616",x"402716",x"3f2616",x"402716",x"3b2415",x"3c2415",x"3a2313",x"3d2615",x"3e2616",x"422818",x"432a1a",x"462c1c",x"492e1c",x"422a1b",x"452d1b",x"452c1c",x"462d1d",x"472f1d",x"432b1b",x"432b1c",x"3a271b",x"432c1d",x"442d1e",x"452f1e",x"452e1f",x"442d1f",x"422d1f",x"442f20",x"472f1f",x"3f2b1e",x"402b1e",x"402c1f",x"462f21",x"432e21",x"412f22",x"402d1f",x"3d2b1e",x"3c2c20",x"3a2a1f",x"3b2a1f",x"38291f",x"38291e",x"34281e",x"382a1f",x"3f2f20",x"38291e",x"372a1f",x"291d15",x"1b120b",x"160f07",x"422d1f",x"452e1e",x"452f20",x"442f21",x"3f2b1f",x"412d20",x"433022",x"422e21",x"412e20",x"3f2e21",x"3b2d20",x"3c2c20",x"3b2b1e",x"392a1e",x"37291f",x"36291f",x"35291f",x"32281d",x"30271d",x"372a1f",x"35291f",x"35291f",x"36291d",x"2c2118",x"1e150d",x"170f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"412511",x"412511",x"412511",x"361f0e",x"412612",x"3d230f",x"150e07",x"1c1108",x"180f07",x"180f07",x"180f07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4f2c14",x"150e07",x"472912",x"29170a",x"150e07",x"150e07",x"150e07",x"150e07",x"462611",x"231409",x"170f07",x"150e07",x"150e07",x"422410",x"331c0b",x"281509",x"2b170a",x"29160a",x"2d180a",x"2e1a0b",x"321c0d",x"351f0e",x"2d1a0c",x"331d0d",x"321d0d",x"2e1a0c",x"2b190b",x"150e07",x"150e07",x"432711",x"201309",x"25160a",x"150e07",x"150e07",x"38200e",x"3b220f",x"150e07",x"301c0c",x"301b0c",x"2c190b",x"2a180b",x"2a180b",x"1c1108",x"150e07",x"231409",x"150e07",x"231409",x"2c190b",x"2e1a0b",x"2d190b",x"27160a",x"150e07",x"1d1208",x"1a1108",x"150e07",x"150e07",x"150e07",x"2d1a0d",x"391f0f",x"231409",x"241409",x"2a170a",x"2f190b",x"321c0c",x"311b0b",x"2d190a",x"29170a",x"271509",x"271509",x"28160a",x"281609",x"261509",x"261509",x"251509",x"231409",x"231409",x"231409",x"221409",x"1e1208",x"1c1108",x"1e1208",x"201309",x"1f1209",x"201309",x"231509",x"25150a",x"231509",x"24150a",x"25160a",x"231509",x"241509",x"2b180b",x"2e1a0b",x"341e0d",x"341d0d",x"331d0d",x"311b0c",x"2f1a0b",x"2f1a0b",x"2f1a0b",x"2d1a0b",x"2e1a0b",x"331c0c",x"361e0e",x"38200e",x"381f0e",x"371f0e",x"39210e",x"3a210f",x"371f0e",x"301b0b",x"2c180a",x"2b170a",x"2d190a",x"2f1a0b",x"311b0b",x"2d190a",x"2b170a",x"2b170a",x"2d180a",x"2e190b",x"311b0c",x"351e0d",x"39210f",x"3c2311",x"3b220f",x"3a210f",x"361f0e",x"321d0d",x"2d1b0c",x"2d1a0c",x"2b190b",x"26160a",x"211409",x"211309",x"25150a",x"29170a",x"2f1b0c",x"2f1b0c",x"2e1b0c",x"2c190b",x"311c0c",x"3b200e",x"3b200e",x"1d1208",x"39200e",x"402615",x"342012",x"321f12",x"321f13",x"342013",x"362113",x"362113",x"362113",x"352114",x"352114",x"382315",x"3e2616",x"402614",x"412614",x"412614",x"3c2313",x"362011",x"341f10",x"351f10",x"341f11",x"341f11",x"331e11",x"311d10",x"301d10",x"2f1b0e",x"331d0f",x"372010",x"382010",x"371d0e",x"341d0e",x"301c0d",x"2b190c",x"26170c",x"25170b",x"25170b",x"26160b",x"28180c",x"2b1a0d",x"2e1c0d",x"341f11",x"362011",x"362112",x"362012",x"372314",x"372315",x"382314",x"3b2617",x"3c2617",x"3d2719",x"412819",x"452c1a",x"452b1a",x"422918",x"412818",x"412818",x"412716",x"432917",x"3f2615",x"3f2515",x"3d2515",x"382312",x"311e12",x"28190e",x"331f10",x"422511",x"221c15",x"221c15",x"201912",x"201913",x"201a13",x"1f1811",x"201912",x"1e1711",x"1f1811",x"1d1710",x"1b140d",x"171009",x"150e07",x"1c120a",x"1c120a",x"312110",x"342313",x"2a1e15",x"2d1f15",x"342417",x"322417",x"332417",x"342417",x"352416",x"3b2718",x"3a2717",x"392617",x"372416",x"3c2818",x"382517",x"3a2619",x"382517",x"362316",x"382315",x"392417",x"362317",x"352215",x"382414",x"382315",x"382315",x"362113",x"3a2313",x"382112",x"3e2514",x"3e2616",x"3d2617",x"3f2715",x"402817",x"432a19",x"432a17",x"402818",x"3e2717",x"3d2716",x"3b2617",x"372417",x"382517",x"372418",x"392618",x"3b2619",x"3a2719",x"362317",x"382518",x"392518",x"3a2517",x"392618",x"3b2719",x"392517",x"3b2718",x"3e2818",x"3f2819",x"3e281a",x"3e2818",x"3f2817",x"402819",x"3d2718",x"402717",x"422a19",x"452c1a",x"432b19",x"3e2718",x"422918",x"422b1a",x"422918",x"422b19",x"442b19",x"432a1b",x"422a1b",x"472e1c",x"472e1d",x"442c1b",x"412a1a",x"432b1b",x"442c1c",x"482f1c",x"402a1b",x"402a1c",x"3e291c",x"3d291c",x"3f2b1c",x"432d1d",x"432c1d",x"442e1d",x"462f1f",x"442f20",x"402c1f",x"3c2a1e",x"3c291d",x"402e20",x"422d20",x"402c1f",x"412d1f",x"402d1e",x"3f2c20",x"3d2a1f",x"3d2b20",x"402d21",x"402d1f",x"453222",x"433021",x"3b2b1f",x"3b2b1f",x"3b2c20",x"382a1f",x"37291f",x"35281e",x"35281e",x"31271d",x"2f261d",x"312820",x"332920",x"35281f",x"34281d",x"2c2119",x"1d140c",x"170f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"412511",x"412511",x"402310",x"361f0e",x"3e2410",x"3b2210",x"3a210f",x"3f2410",x"3a210f",x"3c220f",x"351d0d",x"351d0c",x"341c0c",x"361d0d",x"341c0c",x"331c0c",x"3e220f",x"452611",x"381f0e",x"2b180b",x"321c0c",x"462711",x"40240f",x"432611",x"3f2310",x"412510",x"150e07",x"1c1108",x"241509",x"1c1108",x"150e07",x"150e07",x"3c210e",x"2b180a",x"452712",x"2e1a0c",x"361e0d",x"331d0d",x"361f0e",x"331d0d",x"311c0d",x"301c0d",x"321d0d",x"2f1b0c",x"2b190b",x"150e07",x"150e07",x"4f2f17",x"2a190b",x"2c1a0b",x"2e1b0d",x"1d1208",x"150e07",x"25160a",x"4d2d15",x"25160a",x"25160a",x"2e1b0d",x"23150a",x"25160a",x"150e07",x"150e07",x"3d2310",x"150e07",x"150e07",x"301c0d",x"211409",x"412611",x"36200e",x"150e07",x"1b1108",x"1d1209",x"150e07",x"150e07",x"150e07",x"39200f",x"2d1a0d",x"301c0e",x"37200f",x"3a2211",x"3d2412",x"3c2413",x"3c2514",x"372113",x"372213",x"362213",x"372213",x"332012",x"331f11",x"311e10",x"2e1c0f",x"2b1a0e",x"29190c",x"29190c",x"28170a",x"27160a",x"271609",x"261609",x"241509",x"241509",x"221409",x"231509",x"28170b",x"2b190b",x"301b0c",x"321c0d",x"2f1b0c",x"29180b",x"29180b",x"301c0c",x"351f0e",x"371f0e",x"331c0c",x"311b0b",x"2f1a0b",x"311b0b",x"311b0b",x"301a0b",x"2f1a0b",x"301b0c",x"331d0c",x"371f0e",x"39200f",x"39200e",x"39200e",x"381f0e",x"391f0e",x"3c220f",x"3b210f",x"3a200e",x"39200e",x"341d0c",x"341d0c",x"341d0c",x"321b0c",x"331c0c",x"331d0d",x"351e0d",x"361e0d",x"38200e",x"3b2210",x"38200e",x"3a210f",x"3d2310",x"3e2411",x"3d2310",x"38200f",x"341e0d",x"331e0e",x"331e0e",x"301c0d",x"29180b",x"25160a",x"26160a",x"29180b",x"2f1b0c",x"321d0d",x"321d0d",x"331d0e",x"301c0d",x"3b200e",x"3d200e",x"3f230f",x"3f230f",x"492a14",x"412613",x"3d2411",x"3c2311",x"3e2412",x"402512",x"402513",x"422713",x"442814",x"432713",x"442814",x"492a14",x"492a14",x"492b15",x"4a2b16",x"472915",x"472914",x"432713",x"442713",x"402412",x"432613",x"432713",x"422613",x"432813",x"452914",x"442813",x"442711",x"472913",x"432611",x"3d220f",x"3a200e",x"381f0e",x"371f0e",x"341d0d",x"321b0c",x"331c0c",x"361e0d",x"351e0d",x"392010",x"392010",x"392110",x"3a2211",x"3c2412",x"3b2312",x"3b2312",x"3e2615",x"3c2413",x"432815",x"452915",x"4a2c18",x"432815",x"412514",x"3e2413",x"3e2312",x"402512",x"402411",x"432614",x"402512",x"402411",x"3e2311",x"3a2110",x"351e0f",x"301d0e",x"3d220f",x"3e210f",x"221c15",x"221c15",x"221c15",x"1f1912",x"201a13",x"201912",x"211a14",x"1f1811",x"1f1811",x"1d1710",x"1b150e",x"171009",x"150e07",x"1c120a",x"1c120a",x"2d1e0f",x"2c2013",x"2e2015",x"352516",x"352618",x"332417",x"322417",x"392718",x"392819",x"3c2817",x"392717",x"3b2819",x"3b2818",x"3d2919",x"3b2719",x"3b2619",x"3e2819",x"3c2819",x"402a1a",x"3c2719",x"3b2718",x"3a2417",x"3f2918",x"3b2517",x"3e2717",x"452b16",x"3f2615",x"3e2616",x"442a18",x"472c18",x"452c1a",x"452b19",x"4e321d",x"4c301b",x"472c1a",x"452b1a",x"412a19",x"452c1a",x"452c19",x"422a1a",x"3f281a",x"3f2819",x"402a1b",x"422b1a",x"412a19",x"432c1c",x"462e1d",x"432b1a",x"432b1b",x"452d1b",x"442b19",x"422b1b",x"41291a",x"412918",x"422a1b",x"432c1a",x"3d2819",x"3f2818",x"402819",x"402818",x"432b19",x"412919",x"432a1a",x"432c1a",x"452b1a",x"452c1a",x"442a19",x"452c1a",x"442c1a",x"482e1c",x"462d1b",x"482f1d",x"462d1c",x"452c1c",x"402a1c",x"3f2819",x"442c1c",x"412a1b",x"472e1c",x"422a1b",x"432b1b",x"402a1c",x"3e2a1c",x"3f2b1d",x"432d1e",x"432d1f",x"432e20",x"452f20",x"462f1f",x"452e20",x"432d20",x"422d1f",x"402d1f",x"422c1e",x"412c1e",x"452f20",x"432c1b",x"453021",x"422e20",x"432f22",x"442f21",x"432e1f",x"432f21",x"402e22",x"3f2e20",x"402e20",x"3d2b1f",x"3c2c20",x"382a1f",x"382b20",x"362a20",x"33281f",x"30271f",x"332920",x"30261d",x"33291f",x"36291f",x"2d231a",x"1f150d",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"402410",x"402410",x"402310",x"3c2311",x"3f2511",x"402511",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331d0d",x"3d220f",x"150e07",x"2d190b",x"381f0d",x"150e07",x"150e07",x"170f07",x"472711",x"2c190b",x"150e07",x"231409",x"1b1108",x"150e07",x"241409",x"3b200d",x"29170a",x"3c220f",x"26160a",x"2f1a0b",x"2d190b",x"301a0b",x"2c190b",x"2e1a0c",x"2d190b",x"2e190b",x"2e1b0c",x"211409",x"150e07",x"150e07",x"472914",x"27170a",x"2c1a0b",x"2b190c",x"25160a",x"1d1208",x"150e07",x"150e07",x"4e2c15",x"331d0d",x"150e07",x"150e07",x"150e07",x"432510",x"150e07",x"180f07",x"1c1108",x"150e07",x"150e07",x"2b190b",x"150e07",x"3e2411",x"150e07",x"2a180b",x"1d1208",x"150e07",x"150e07",x"150e07",x"372113",x"381f0f",x"2f1c0f",x"341e0f",x"382112",x"3a2212",x"392111",x"372113",x"311e12",x"2e1d11",x"2e1d13",x"2e1d12",x"2e1d11",x"301d11",x"311e11",x"311e10",x"2f1d0f",x"2a190c",x"27170b",x"28160a",x"2b180a",x"2c190b",x"2a180b",x"27170a",x"26160a",x"26160a",x"26160a",x"2e1a0b",x"29170a",x"311c0c",x"341e0f",x"331d0e",x"2d1b0d",x"2f1c0e",x"301d0f",x"351f11",x"3a2312",x"3b2414",x"382212",x"362113",x"321d11",x"342012",x"331f11",x"311d10",x"331f11",x"382213",x"3b2413",x"3c2313",x"3a2313",x"392212",x"392212",x"3a2312",x"3c2313",x"3c2313",x"3b2212",x"382212",x"372112",x"341e0f",x"341e0f",x"331e0f",x"341f10",x"372010",x"382011",x"382111",x"331d0f",x"331e0f",x"331e10",x"341f10",x"362011",x"341d0e",x"382010",x"3c2311",x"37200f",x"361f0f",x"37200f",x"321d0d",x"2b190b",x"27170a",x"27170b",x"2a190b",x"2f1b0c",x"301b0c",x"321c0d",x"361f0e",x"351f0e",x"462712",x"371f0e",x"371f0e",x"38200f",x"3d210f",x"38210f",x"38200f",x"331d0e",x"311c0d",x"331d0d",x"36200e",x"37200f",x"341e0d",x"331d0d",x"341d0d",x"371e0d",x"381e0d",x"3b200e",x"3d210f",x"3a200d",x"3a200d",x"361d0c",x"391f0d",x"391f0d",x"3b200e",x"361d0c",x"351c0c",x"331b0b",x"341c0c",x"381f0d",x"3a200e",x"412410",x"422511",x"3f2410",x"371f0d",x"301a0b",x"2f1a0b",x"2d190b",x"2f1a0b",x"321c0d",x"321d0d",x"321d0d",x"331d0d",x"331d0d",x"321d0d",x"311c0c",x"311c0c",x"311c0c",x"301b0c",x"311c0c",x"351f0e",x"371f0e",x"371e0d",x"3c210f",x"3e2410",x"3e2310",x"3c210e",x"381e0d",x"391f0d",x"3b200e",x"3a200e",x"3a200e",x"3b210f",x"38200e",x"331d0c",x"2b180b",x"231409",x"1c1108",x"361d0d",x"221b15",x"221b15",x"221b15",x"211a14",x"201913",x"201912",x"201a13",x"1e1711",x"1e1711",x"1c150f",x"1b140d",x"19120c",x"150e07",x"1a110a",x"1a110a",x"2e1f11",x"332315",x"2a2017",x"2e2115",x"382717",x"352518",x"3b2818",x"3e2a19",x"3b2818",x"3e2a19",x"3e2918",x"412a19",x"432c19",x"402a1a",x"3e2819",x"3e2819",x"3e2819",x"442b1b",x"422a1a",x"3c2719",x"3b2618",x"3d2718",x"412a1a",x"3c2515",x"462b19",x"422a18",x"432a18",x"402715",x"442a18",x"472d1a",x"482e1b",x"432b19",x"452c1a",x"462c19",x"432a19",x"3f2818",x"3f2718",x"3f2817",x"3d2818",x"3e2719",x"3e2819",x"3c2517",x"422a1a",x"3d2719",x"402919",x"3d2719",x"3c2718",x"3d2719",x"412a1a",x"452d1c",x"472e1b",x"422c1b",x"432c1c",x"3e2819",x"3f2819",x"402a1a",x"40291a",x"452c1b",x"482d1c",x"482e1c",x"4a2f1c",x"482e1c",x"472d1a",x"482d1c",x"432b1b",x"472d1c",x"452c1a",x"452c1a",x"492f1d",x"4a2f1c",x"442b1b",x"482f1c",x"472e1d",x"4a301d",x"482f1d",x"432b1a",x"422b1b",x"442d1c",x"472e1d",x"40291a",x"472e1d",x"432b1b",x"442e1d",x"422b1d",x"442c1c",x"422d1e",x"432d1f",x"462f20",x"452f20",x"462f20",x"452f20",x"463122",x"442f20",x"442f20",x"422e20",x"452f20",x"473020",x"483122",x"432d1f",x"422f21",x"3e2c1f",x"422f21",x"442e1f",x"432e21",x"3f2c20",x"3d2b1f",x"402d20",x"433023",x"3f2c1f",x"3c2d20",x"3d2e21",x"35291f",x"34291f",x"382b21",x"32271e",x"352920",x"33271d",x"2b2018",x"20170f",x"180f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"412511",x"412511",x"422411",x"39210f",x"412512",x"482a13",x"231509",x"29170b",x"2a180a",x"2e1b0c",x"29180b",x"28170a",x"201309",x"29180b",x"28170a",x"211309",x"150e07",x"150e07",x"442611",x"150e07",x"432712",x"150e07",x"170f07",x"1a1008",x"150e07",x"150e07",x"150e07",x"472811",x"180f08",x"150e07",x"150e07",x"42240f",x"150e07",x"150e07",x"29170a",x"2d190b",x"311b0c",x"321c0c",x"2d190b",x"2d190a",x"2b180a",x"2d190b",x"2d1a0b",x"2a180b",x"24150a",x"150e07",x"3c220f",x"29180b",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"462811",x"3a200e",x"331c0c",x"432611",x"311b0c",x"2d1a0b",x"2f1b0c",x"2a180b",x"180f07",x"150e07",x"351e0d",x"2a180b",x"150e07",x"29180b",x"1f1309",x"150e07",x"150e07",x"150e07",x"3a2110",x"362010",x"332115",x"3d2718",x"3f2818",x"3f2919",x"372316",x"2f1f15",x"281c14",x"211912",x"1d1610",x"1d1610",x"1d1610",x"1c150e",x"1c150e",x"1a140c",x"20150d",x"24160b",x"29180c",x"2d1b0d",x"2d190b",x"2d1a0b",x"2b190b",x"27160a",x"221409",x"221409",x"211309",x"241509",x"2a190b",x"301c0e",x"341e0f",x"352011",x"2f1e11",x"2c1d12",x"312115",x"342014",x"3a2517",x"3b2719",x"3c271a",x"3b2619",x"3a2618",x"352316",x"2f2117",x"261c14",x"251c15",x"2c1f15",x"362417",x"402919",x"3f291a",x"3f2819",x"3e2617",x"3e2617",x"3e2718",x"3f2718",x"412819",x"3d2515",x"3b2515",x"382214",x"352215",x"2d1c12",x"2d1d12",x"332014",x"332115",x"301f14",x"2f1e13",x"2f1e12",x"2a1a0f",x"24190f",x"1d160f",x"1c150e",x"19120b",x"181109",x"24160c",x"2d1a0b",x"321d0d",x"301c0d",x"2b190b",x"25150a",x"241509",x"231308",x"1f1107",x"201107",x"251408",x"261509",x"211309",x"351e0d",x"381f0e",x"381f0e",x"38200f",x"371e0d",x"361e0c",x"371f0e",x"341d0d",x"2d1a0b",x"2d1a0b",x"301b0c",x"2f1a0b",x"2e1a0b",x"311c0c",x"331d0d",x"39200f",x"3e230f",x"422511",x"422511",x"422510",x"422611",x"432612",x"432612",x"422611",x"3f2410",x"3e230f",x"3f2310",x"3d220f",x"3b200e",x"3c210f",x"3d210f",x"422511",x"432611",x"3f230f",x"3c210f",x"361e0d",x"361f0e",x"341d0d",x"321c0c",x"321c0d",x"311b0c",x"301b0c",x"301b0c",x"311b0c",x"2f1b0b",x"301b0c",x"301b0c",x"2d1a0c",x"2b190b",x"2b190b",x"2e1b0c",x"361f0e",x"381f0e",x"39200e",x"3a210f",x"3a210f",x"3b210f",x"3c220f",x"3c220f",x"381f0e",x"371e0d",x"371f0e",x"371f0e",x"361f0e",x"341e0d",x"2c190b",x"241509",x"1c1108",x"3d2210",x"221b14",x"221b14",x"221c15",x"231c16",x"211a14",x"1f1812",x"211a14",x"1f1811",x"1f1912",x"1d1710",x"1b140e",x"19120b",x"150e07",x"20140a",x"1d130a",x"271b0f",x"302215",x"2c2017",x"2f2016",x"362516",x"392719",x"392718",x"3c2818",x"3b2818",x"3f2b19",x"342416",x"392718",x"3c2717",x"322216",x"312115",x"2e2016",x"362417",x"3a2517",x"3a2517",x"3a2518",x"3b2518",x"3f2817",x"3d2717",x"3d2717",x"3a2517",x"3c2515",x"402817",x"3d2515",x"412816",x"402817",x"422918",x"462c19",x"4a2f1b",x"4a301c",x"492e1b",x"472d1b",x"432b19",x"462d1b",x"442d1a",x"452d1a",x"452d1c",x"452d1d",x"452e1d",x"422b1c",x"482e1b",x"442d1c",x"422b1b",x"442c1c",x"412a1c",x"452c1b",x"442b1a",x"432b1c",x"442d1c",x"422c1c",x"452c1b",x"482f1d",x"452d1a",x"422a1a",x"482d1b",x"452c1a",x"492f1c",x"452d1b",x"432b1b",x"432b1a",x"442c1a",x"462d1a",x"452c1a",x"482e1c",x"452e1d",x"4a2f1c",x"472e1c",x"432a1b",x"452c1c",x"472e1b",x"482f1c",x"472e1b",x"4b311e",x"472e1c",x"462d1d",x"422b1c",x"452d1d",x"422c1c",x"432c1d",x"462f1f",x"442d1c",x"452f1f",x"442e1e",x"452f20",x"483021",x"473020",x"472e1d",x"473021",x"463020",x"462f1f",x"432d1f",x"3e2b1d",x"432e1f",x"412d1f",x"432f21",x"433022",x"412e20",x"412f21",x"3e2d20",x"3f2d21",x"3c2b1e",x"412e22",x"3f2d21",x"3d2b1f",x"3e2d21",x"392a20",x"382c22",x"35281e",x"352a21",x"31281f",x"332921",x"362b20",x"31271f",x"281f18",x"1e150e",x"170f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3e220f",x"3e220f",x"3f2310",x"38200f",x"402612",x"462812",x"29180b",x"321c0d",x"351f0d",x"311c0d",x"311c0d",x"2f1b0c",x"311c0d",x"2e1a0b",x"2e1a0b",x"2c1a0c",x"2b190b",x"150e07",x"150e07",x"462812",x"2d1a0b",x"27170a",x"2d1a0b",x"2a190b",x"2c190b",x"1c1108",x"150e07",x"150e07",x"4a2a13",x"150e07",x"3c210e",x"1a1008",x"150e07",x"3a210f",x"2c190b",x"311b0c",x"331d0d",x"331c0c",x"2e1a0b",x"311c0c",x"2e1a0b",x"2b180b",x"231409",x"150e07",x"150e07",x"150e07",x"3b210f",x"150e07",x"150e07",x"150e07",x"432511",x"422510",x"432410",x"371d0c",x"3d200d",x"3c200e",x"341d0c",x"150e07",x"321c0c",x"251509",x"371d0c",x"1c1108",x"251509",x"27160a",x"27160a",x"211309",x"150e07",x"150e07",x"150e07",x"150e07",x"2b180b",x"211409",x"150e07",x"150e07",x"150e07",x"362010",x"362113",x"221911",x"2f1f14",x"362316",x"3a2516",x"362316",x"332216",x"2b1d14",x"241a12",x"201811",x"1d1710",x"1d1711",x"1d160f",x"1b150e",x"1b140d",x"1c150f",x"1a130c",x"1f150c",x"25170b",x"2b190d",x"2b180c",x"27170b",x"22150b",x"19110a",x"171009",x"171009",x"19110a",x"22160d",x"2c1b0f",x"321f11",x"2d1d12",x"231a12",x"251c15",x"2c1f15",x"352418",x"3a2619",x"3c281b",x"3b271a",x"3c291c",x"39271b",x"342419",x"2e2319",x"282019",x"261f18",x"2c221a",x"31251b",x"332419",x"35251a",x"34241a",x"362519",x"38271c",x"36261a",x"38281d",x"3a291d",x"35261b",x"2e231a",x"272019",x"28211a",x"28211a",x"29221b",x"29221b",x"27211a",x"29221c",x"29231c",x"2b241d",x"2a231c",x"2a241d",x"2a241c",x"2a231c",x"2a241d",x"29221b",x"2b221a",x"32261d",x"32241a",x"2f2219",x"281f18",x"261f17",x"292019",x"2a221a",x"2a211a",x"2c221a",x"2f251d",x"352d25",x"2e261e",x"3b1f0d",x"2b180b",x"26160a",x"221409",x"221409",x"331c0c",x"331c0c",x"2b180a",x"251509",x"261509",x"271609",x"271509",x"271509",x"29160a",x"301b0b",x"361f0d",x"3b210f",x"3e230f",x"3e230f",x"412410",x"3f2310",x"3e230f",x"3f2310",x"3f2310",x"3e2410",x"3e230f",x"3f2410",x"3f2410",x"3c220f",x"3c210f",x"412411",x"412510",x"3f230f",x"412510",x"3c220f",x"351d0d",x"321c0c",x"301b0c",x"2d190b",x"2c180a",x"301b0c",x"301b0c",x"311c0d",x"311c0d",x"321d0d",x"311c0d",x"311c0d",x"2d1a0c",x"29180b",x"26150a",x"28160a",x"2d190b",x"331c0c",x"351e0d",x"371f0e",x"361e0e",x"361e0d",x"351d0d",x"331c0c",x"311b0b",x"301a0b",x"301a0b",x"341d0d",x"361f0e",x"331d0d",x"2c1a0c",x"231509",x"1b1108",x"422511",x"221c15",x"221c15",x"211b14",x"231c16",x"201a13",x"1f1811",x"211b14",x"1f1811",x"1e1711",x"1d1610",x"1b150e",x"19120b",x"150e07",x"20150a",x"21160b",x"2b1d0f",x"302115",x"291e14",x"2c2016",x"332416",x"332417",x"382717",x"372718",x"342416",x"402b19",x"362519",x"352315",x"382617",x"372517",x"362518",x"342215",x"372417",x"372517",x"372416",x"3a2417",x"392518",x"3b2717",x"382416",x"352215",x"3a2516",x"3a2415",x"3b2515",x"382315",x"372214",x"3b2515",x"3e2818",x"3f2918",x"452b19",x"482e19",x"452d1a",x"432a19",x"432a1a",x"452d1c",x"462e1c",x"432b1a",x"402919",x"442d1d",x"422b1c",x"432c1d",x"422c1c",x"3e291b",x"3d2719",x"432b1a",x"3d2819",x"442c1a",x"442c1b",x"432b1b",x"412a1a",x"452d1d",x"482f1c",x"442c1c",x"462d1c",x"402919",x"402919",x"432b1b",x"432a19",x"40291b",x"422b1a",x"412a1a",x"442c1b",x"432c1c",x"442c1b",x"442c1b",x"432b19",x"462d1c",x"462e1c",x"452d1b",x"452d1c",x"4b311e",x"472e1d",x"462e1c",x"492f1d",x"472f1e",x"4b321f",x"482f1e",x"452e1e",x"432c1c",x"462d1e",x"493020",x"452e1d",x"452f20",x"4a3322",x"4a3322",x"483020",x"483120",x"462e1c",x"483121",x"483221",x"473021",x"473121",x"4b3322",x"4a3222",x"443021",x"432f1f",x"453022",x"443023",x"453123",x"402d1f",x"402e21",x"412e21",x"3f2d20",x"3c2b1f",x"3d2c20",x"3a2b1f",x"3a2c21",x"3b2c21",x"3a2b21",x"352a20",x"332920",x"33281f",x"31261c",x"342920",x"2c231b",x"1f160f",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3c210e",x"3c210e",x"412410",x"361f0e",x"3f2411",x"4c2d15",x"2a180b",x"371f0e",x"361f0e",x"351e0d",x"341e0e",x"28170b",x"371f0f",x"361f0e",x"211409",x"28160a",x"29180b",x"1e1209",x"150e07",x"150e07",x"321d0d",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"2d1a0c",x"2c190b",x"1c1108",x"150e07",x"150e07",x"4f2e16",x"311c0d",x"1e1209",x"150e07",x"2b180b",x"341c0c",x"27160a",x"2d190b",x"311c0c",x"2f1c0c",x"321d0d",x"2b190c",x"1e1209",x"150e07",x"27170b",x"2f1c0d",x"211409",x"150e07",x"472711",x"3b210e",x"311c0c",x"3a200e",x"3f230f",x"361f0e",x"321c0d",x"321c0c",x"3c210e",x"2d190b",x"211309",x"2d190b",x"3d220f",x"462711",x"201309",x"241509",x"301c0c",x"2c190b",x"2b190b",x"1d1108",x"150e07",x"39200f",x"150e07",x"2a180b",x"1c1108",x"150e07",x"150e07",x"150e07",x"28180c",x"25170b",x"2f1d0f",x"201912",x"251b12",x"2c1f15",x"2f2015",x"2c1e14",x"281d15",x"201811",x"1e1811",x"1d160f",x"1d160f",x"1d1610",x"20170f",x"1b140d",x"1c130c",x"20150d",x"171009",x"181109",x"1f130b",x"27170a",x"2c190b",x"25160a",x"180f07",x"190f08",x"150e07",x"150e07",x"180f08",x"27190d",x"321e0f",x"2f1d10",x"22180f",x"1f1810",x"241a12",x"271c13",x"2c1f15",x"2d2016",x"2b1f15",x"2e2117",x"2b1e14",x"291f16",x"251c15",x"231c15",x"221b15",x"221b15",x"241c15",x"281e15",x"291e14",x"2f2016",x"37261a",x"392517",x"372417",x"382518",x"3a2617",x"3e2716",x"3d2715",x"3b2515",x"392314",x"3a2414",x"392213",x"362112",x"362011",x"341f12",x"321e12",x"311d10",x"362012",x"362112",x"392314",x"372212",x"362212",x"362111",x"372011",x"362010",x"361f10",x"331d0e",x"2f1b0d",x"301c0d",x"2e1a0d",x"311c0d",x"311b0d",x"2e1a0b",x"27160a",x"2a180b",x"2c190b",x"2e190b",x"2b180b",x"26160a",x"221409",x"221409",x"2a180b",x"2e1b0c",x"311c0d",x"331d0d",x"321d0d",x"301c0c",x"2d1a0c",x"2f1b0c",x"2f1b0c",x"301b0b",x"361f0d",x"3b210f",x"3e230f",x"3e230f",x"412410",x"3f2310",x"3e230f",x"3f2310",x"3f2310",x"3e2410",x"3e230f",x"3f2410",x"3f2410",x"3c220f",x"3c210f",x"412411",x"412510",x"3f230f",x"412510",x"3c220f",x"351d0d",x"321c0c",x"301b0c",x"2d190b",x"2c180a",x"301b0c",x"301b0c",x"311c0d",x"311c0d",x"321d0d",x"311c0d",x"311c0d",x"2d1a0c",x"29180b",x"26150a",x"28160a",x"2d190b",x"331c0c",x"351e0d",x"371f0e",x"361e0e",x"361e0d",x"351d0d",x"331c0c",x"311b0b",x"301a0b",x"301a0b",x"341d0d",x"361f0e",x"331d0d",x"2c1a0c",x"231509",x"1b1108",x"422511",x"211b15",x"211b15",x"211a13",x"221b15",x"201a13",x"201a13",x"1f1811",x"1f1812",x"1f1811",x"1d1610",x"1b150e",x"19130c",x"150e07",x"1d130a",x"1d130a",x"281b10",x"281d12",x"281e15",x"2e2116",x"342618",x"342619",x"342516",x"332417",x"342518",x"362619",x"342517",x"342518",x"332416",x"352416",x"392617",x"372316",x"362317",x"382316",x"392618",x"392619",x"3c2819",x"3e2918",x"3e2919",x"392517",x"412a18",x"412a19",x"3c2617",x"3d2614",x"422817",x"432a18",x"452c1a",x"462d1b",x"492e1b",x"482e1b",x"482d1a",x"472d1a",x"452d1c",x"462d1b",x"472e1b",x"452d1b",x"432b1a",x"412b1b",x"41291a",x"422b1c",x"432b1b",x"422c1c",x"452e1c",x"452c1b",x"432c1d",x"442d1d",x"412b1c",x"402a1a",x"432c1b",x"422b1c",x"432b1b",x"422a1b",x"432b1b",x"452d1c",x"442c1b",x"452d1d",x"412a1a",x"442b1a",x"472e1c",x"452d1b",x"452c1a",x"432c1a",x"432c1b",x"442c1a",x"442d1b",x"452e1b",x"452e1c",x"432b1b",x"432d1d",x"462e1c",x"432c1c",x"462e1c",x"482f1d",x"472e1d",x"422d1d",x"442d1c",x"472f1e",x"472f1f",x"452f20",x"432e1f",x"473020",x"452e1e",x"47301f",x"473120",x"493120",x"4a3120",x"4e3422",x"4c3524",x"503623",x"4b3221",x"4c3423",x"4a3320",x"483222",x"422d1f",x"422f21",x"402c1f",x"422f22",x"483222",x"463121",x"443123",x"422f22",x"443121",x"3f2c1f",x"433022",x"412f21",x"3b2b1f",x"392a20",x"35281f",x"31271e",x"332920",x"342920",x"352a20",x"36281d",x"2d221a",x"20170f",x"180f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3a200e",x"3a200e",x"422511",x"351e0e",x"3c2310",x"452712",x"28170a",x"361f0e",x"2f1b0c",x"301b0c",x"37200f",x"3c2310",x"341e0d",x"2f1a0b",x"2c180b",x"2c180b",x"26160a",x"150e07",x"150e07",x"371f0e",x"2f1b0c",x"2b190b",x"311c0d",x"2d1a0c",x"2d1a0c",x"24150a",x"150e07",x"150e07",x"321d0d",x"201309",x"1e1208",x"2b190b",x"221409",x"150e07",x"4f2c14",x"2f1b0c",x"2a190b",x"2a180b",x"2a190b",x"28170a",x"1d1208",x"150e07",x"3d2411",x"311c0d",x"2c190b",x"482a14",x"2e1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"43240f",x"1b1108",x"3d220e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2a170a",x"3a1f0d",x"170f07",x"1e1208",x"26160a",x"28170a",x"221409",x"150e07",x"150e07",x"150e07",x"29180b",x"1d1108",x"150e07",x"150e07",x"150e07",x"2d1b0d",x"2d1b0d",x"321d0e",x"372011",x"3c2312",x"402614",x"3e2513",x"3c2313",x"3a2314",x"372213",x"332012",x"332013",x"342112",x"352113",x"331f11",x"311e11",x"2f1d11",x"2d1c0f",x"2b1a0e",x"28170c",x"28180b",x"28180c",x"281609",x"271509",x"2b180b",x"2a180b",x"2a190b",x"28180b",x"26170a",x"26160a",x"27170a",x"2c190b",x"2d1a0c",x"311c0d",x"351f0e",x"331d0d",x"2b190b",x"2a180b",x"2f1b0c",x"331d0d",x"331c0d",x"341c0d",x"331c0d",x"341d0d",x"37200e",x"39210f",x"37200e",x"351e0d",x"351e0e",x"331d0d",x"341e0e",x"37200f",x"3d2411",x"3f2411",x"402511",x"412612",x"3f2411",x"3f2410",x"3e2310",x"3d220f",x"3f2410",x"402410",x"3e2310",x"402512",x"3e2411",x"3d2411",x"3c2310",x"3b220f",x"3b2310",x"3c2310",x"3b2210",x"3a2210",x"3a2210",x"3c2310",x"3b220f",x"361e0d",x"341c0d",x"351d0c",x"371e0d",x"361e0d",x"341c0c",x"351d0c",x"321b0c",x"2e190b",x"2d190b",x"2d190b",x"2a170a",x"251509",x"211308",x"241509",x"29170a",x"29170a",x"2f1b0b",x"2f1a0b",x"301b0c",x"2f1a0b",x"301b0c",x"2f1b0c",x"2e1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221b14",x"221b14",x"201912",x"221c15",x"201a13",x"201a13",x"201a13",x"1f1811",x"1e1811",x"1c150f",x"1b140e",x"19120c",x"150e07",x"2d231a",x"2b2119",x"31251a",x"2e2318",x"362819",x"342518",x"322519",x"342518",x"342619",x"352619",x"37271a",x"332519",x"38271a",x"372619",x"3a281a",x"392719",x"3a2719",x"382518",x"382518",x"382619",x"3a2719",x"3b281a",x"372518",x"402a1a",x"3d291a",x"3d2818",x"3e291a",x"432c1c",x"442c1b",x"40291a",x"432a18",x"482e1b",x"472f1e",x"462d1b",x"4a301c",x"4c311d",x"482f1c",x"482f1d",x"492e1c",x"472e1c",x"472e1c",x"412a1a",x"432c1c",x"422c1c",x"452d1d",x"432c1b",x"472e1d",x"452d1c",x"452d1c",x"462d1c",x"452d1b",x"472f1d",x"432d1d",x"432a1a",x"442c1c",x"452d1d",x"462d1c",x"412b1b",x"432b19",x"40291a",x"402a1b",x"3d2819",x"452c1a",x"472e1c",x"462f1c",x"472d1c",x"4a311d",x"452e1d",x"422c1b",x"432d1b",x"432d1d",x"452d1b",x"49301d",x"482f1d",x"462d1c",x"4b321d",x"482f1b",x"4b311d",x"492f1c",x"4b301c",x"432d1c",x"432d1d",x"452f1f",x"48301f",x"462f20",x"453021",x"483121",x"4a3120",x"4b3220",x"4b3321",x"4d3422",x"4b3320",x"4d3422",x"4c3322",x"4d3524",x"4a3222",x"493222",x"4b3322",x"4c3320",x"493221",x"483221",x"4a3220",x"493323",x"473121",x"463223",x"453021",x"453222",x"412e21",x"412e20",x"412d20",x"412e22",x"3b2b1f",x"3a2b1f",x"38291f",x"34291f",x"382c22",x"362b21",x"382b20",x"362a21",x"31251b",x"241910",x"1a110a",x"1a120b",x"1a120b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"391f0e",x"391f0e",x"432611",x"38200f",x"3e2310",x"462711",x"1a1008",x"2d190b",x"2c190b",x"2a180b",x"28170a",x"29180b",x"2c190b",x"150e07",x"1a1008",x"150e07",x"150e07",x"150e07",x"39200f",x"150e07",x"4e2d15",x"28170b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"573419",x"150e07",x"26160a",x"2e1b0c",x"2e1b0c",x"2d1b0c",x"150e07",x"150e07",x"523017",x"2a190b",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0c",x"3b2210",x"482913",x"351e0e",x"1d1208",x"25160a",x"2c1a0c",x"2c190b",x"27160a",x"231409",x"150e07",x"150e07",x"150e07",x"1f1208",x"180f07",x"2a180a",x"29170a",x"251509",x"1d1108",x"150e07",x"150e07",x"3c210f",x"37200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2310",x"25150a",x"1e1108",x"150e07",x"150e07",x"150e07",x"311b0b",x"331d0e",x"351e0f",x"3b2212",x"3e2412",x"402512",x"3f2514",x"3d2513",x"3b2415",x"382214",x"362214",x"331f12",x"342114",x"331f12",x"331f12",x"321f11",x"301e11",x"2d1b0f",x"2c1b0f",x"2c1a0d",x"2d1b0d",x"2e1a0d",x"2d190b",x"2c190b",x"2d1a0b",x"2c1a0b",x"2b190b",x"29180b",x"29180b",x"2a190b",x"2d1a0c",x"2f1b0c",x"2f1a0c",x"301b0c",x"331c0d",x"321c0c",x"2e1a0b",x"2b180b",x"2e1a0c",x"331d0d",x"341d0d",x"331c0c",x"331c0c",x"341d0d",x"331d0d",x"351d0d",x"39210f",x"38210f",x"37200e",x"361f0e",x"371f0e",x"39210f",x"3e2310",x"432712",x"442913",x"442813",x"432712",x"422712",x"422612",x"422612",x"422612",x"412511",x"412611",x"432712",x"3f2511",x"3e2411",x"3d2310",x"3d2310",x"3d2310",x"3c2310",x"39210f",x"39200f",x"3a210f",x"3d2310",x"3e2411",x"3a220f",x"38200e",x"381f0e",x"3b200f",x"3a200e",x"3a200e",x"361e0d",x"341d0d",x"321c0c",x"331c0d",x"331d0d",x"2f1a0b",x"2a180a",x"251509",x"251509",x"2b190b",x"301c0d",x"301b0c",x"341e0d",x"341d0d",x"321c0d",x"311c0c",x"301c0c",x"2e190b",x"2c190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231c15",x"231c15",x"221b15",x"221c15",x"211b15",x"201913",x"201913",x"1f1812",x"1e1711",x"1d160f",x"1a140d",x"17110a",x"150e07",x"53483e",x"53473d",x"4f453a",x"42372d",x"3d3125",x"443528",x"3c3025",x"3e3023",x"3e3025",x"433223",x"3f3125",x"3c2e23",x"3e3024",x"3c2e23",x"413327",x"403125",x"423124",x"423125",x"443327",x"443225",x"453326",x"433123",x"433124",x"453223",x"413024",x"4b3828",x"533c2b",x"503d2d",x"523e2f",x"554131",x"57402f",x"533d2c",x"4f3a2b",x"4e3929",x"513a2a",x"4f3728",x"4f3826",x"503927",x"4d3727",x"4e3524",x"513927",x"4e3625",x"463122",x"463021",x"4a3324",x"463121",x"483223",x"473121",x"4a3323",x"493221",x"4c3524",x"483121",x"4a3221",x"4a3321",x"483121",x"49311e",x"483021",x"4b3321",x"4a3323",x"4a311f",x"472f1d",x"463222",x"493120",x"4a3222",x"483222",x"4a3222",x"4c3523",x"493322",x"483323",x"412e20",x"453122",x"4a3424",x"4a3323",x"473222",x"442e20",x"483220",x"483121",x"483122",x"493221",x"493120",x"493325",x"483425",x"4b3628",x"4a3728",x"4e3929",x"4c3829",x"4d3727",x"4f3827",x"533b2a",x"503827",x"543b28",x"563c29",x"533a29",x"513a29",x"513927",x"4f3828",x"513928",x"4e3827",x"4f3828",x"4b3525",x"503826",x"4d3626",x"4a3323",x"4b3524",x"4a3423",x"463222",x"463120",x"453224",x"443124",x"433122",x"473323",x"413023",x"423123",x"3b2c21",x"382d23",x"36291f",x"3b2d20",x"3f2f20",x"3b2f25",x"433225",x"41362c",x"41382f",x"41382f",x"41382f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3b200e",x"3b200e",x"412511",x"341e0d",x"3a220f",x"351d0d",x"1f1209",x"1c1108",x"1e1208",x"1f1209",x"1f1209",x"1c1108",x"211309",x"150e07",x"1d1208",x"170f07",x"211409",x"432611",x"391f0e",x"28170a",x"2b180a",x"40230f",x"2a180a",x"1d1108",x"381f0e",x"462711",x"150e07",x"150e07",x"2a180b",x"29170a",x"2d190b",x"29170a",x"27160a",x"211409",x"150e07",x"150e07",x"27170a",x"391f0e",x"27160a",x"1e1208",x"39200e",x"311b0c",x"28160a",x"1e1208",x"1a1008",x"251509",x"211308",x"2a170a",x"28160a",x"241409",x"26150a",x"170f07",x"150e07",x"3e210f",x"180f07",x"29170a",x"2c180a",x"251509",x"29170a",x"28170a",x"241509",x"150e07",x"150e07",x"150e07",x"2e1a0b",x"3f2410",x"211309",x"150e07",x"150e07",x"2a180a",x"231509",x"180f07",x"150e07",x"150e07",x"150e07",x"351e0e",x"331d0e",x"392010",x"3f2513",x"3f2412",x"3b2111",x"3c2413",x"3b2313",x"382212",x"331f11",x"311e12",x"2f1d11",x"301d11",x"321f11",x"331f11",x"301d0f",x"2e1c0f",x"2d1b0e",x"2b190c",x"2b180c",x"2c1a0d",x"2e1b0d",x"2e1a0b",x"2d190b",x"2d1a0b",x"2d1a0b",x"2b190b",x"261509",x"28170a",x"28170a",x"2d1a0b",x"2f1b0b",x"301b0c",x"311c0c",x"341d0d",x"361f0e",x"311c0d",x"2d1a0b",x"2f1a0c",x"331d0d",x"361e0d",x"381f0e",x"38200f",x"37200e",x"351d0d",x"331c0c",x"331c0d",x"321c0c",x"311b0b",x"311b0c",x"331c0c",x"361e0d",x"3a200f",x"3b210f",x"3c220f",x"3c220f",x"3c210f",x"3b200e",x"3b200e",x"3a200e",x"3a200e",x"3b210e",x"3c210f",x"3a210e",x"381f0e",x"371e0d",x"381f0e",x"371e0d",x"361e0d",x"341c0c",x"351d0d",x"341d0d",x"321c0c",x"321b0b",x"341d0c",x"341d0c",x"321b0c",x"321b0b",x"341d0c",x"361e0d",x"371e0d",x"361d0d",x"351d0c",x"2f1a0b",x"2e190b",x"321b0c",x"311b0b",x"2d1a0b",x"28170a",x"261609",x"29170a",x"2e1a0c",x"311c0c",x"311b0c",x"301b0b",x"301b0b",x"2e1a0b",x"301b0c",x"2e1a0b",x"2b180a",x"2f1b0c",x"231509",x"231509",x"221409",x"201308",x"1f1308",x"1f1208",x"201308",x"211409",x"211308",x"231409",x"231409",x"241409",x"251509",x"251409",x"251409",x"241409",x"241409",x"241509",x"241509",x"231509",x"221409",x"201308",x"1d1108",x"1a1008",x"190f07",x"1a1008",x"1a1008",x"190f08",x"170f07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221c15",x"221c15",x"231d16",x"221b15",x"201912",x"1f1811",x"201a13",x"1f1811",x"1f1811",x"1d160f",x"1b150e",x"171009",x"150e07",x"574d43",x"564c42",x"4c4136",x"453b31",x"40362c",x"413225",x"433223",x"423326",x"3f3125",x"433224",x"3d2e22",x"443225",x"3d2e22",x"403125",x"3f2f23",x"433225",x"433227",x"443327",x"413226",x"413227",x"433124",x"402f21",x"453122",x"443020",x"433124",x"483424",x"4d3828",x"503b2c",x"523d2c",x"57402e",x"573e2b",x"543e2e",x"523c2b",x"513c2b",x"543b28",x"563d2b",x"543c29",x"4f3928",x"4d3828",x"4b3727",x"4f3928",x"513927",x"483323",x"463122",x"4a3424",x"4b3524",x"4b3523",x"4a3322",x"483221",x"493323",x"4e3621",x"4a3322",x"4b3320",x"473020",x"452f20",x"473120",x"483221",x"452f20",x"483120",x"483121",x"462f20",x"47301f",x"452f1e",x"483120",x"473020",x"3e2b1c",x"453020",x"442f20",x"422f20",x"412d1f",x"422f21",x"453120",x"473221",x"483221",x"46301f",x"432e1e",x"472f1e",x"422c1e",x"463020",x"452f1e",x"463021",x"473223",x"453021",x"443123",x"443124",x"473425",x"463427",x"4b3627",x"4e3725",x"513927",x"563d29",x"523a28",x"533a27",x"513a27",x"523a28",x"4e3929",x"4b3524",x"503929",x"4a3526",x"513927",x"4f3827",x"4a3526",x"4c3625",x"4b3422",x"4b3525",x"4a3322",x"4c3727",x"463224",x"4a3423",x"463223",x"413022",x"433121",x"423122",x"3e2f23",x"403123",x"3a2b1d",x"402f20",x"473322",x"493523",x"443529",x"483a2f",x"473d34",x"453b32",x"453b32",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"391e0d",x"391e0d",x"432712",x"301b0c",x"361f0f",x"39200e",x"190f08",x"190f08",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"170f07",x"201309",x"4c2c14",x"3f2410",x"2a180b",x"341d0d",x"422510",x"29170a",x"150e07",x"331c0d",x"422410",x"150e07",x"150e07",x"2b180b",x"2e1a0b",x"2d190b",x"2c190b",x"221409",x"150e07",x"150e07",x"150e07",x"211308",x"361d0d",x"28170a",x"1f1208",x"3b210f",x"371f0e",x"2b180a",x"27160a",x"180f07",x"2b180b",x"2f1b0c",x"2c190b",x"2a170a",x"2a170a",x"201309",x"150e07",x"150e07",x"361d0c",x"191008",x"1f1208",x"211309",x"251509",x"251509",x"201208",x"1a1008",x"150e07",x"150e07",x"150e07",x"301b0c",x"39200e",x"26160a",x"150e07",x"150e07",x"321c0c",x"26160a",x"1e1208",x"150e07",x"150e07",x"341e0e",x"2f1a0c",x"2f190c",x"331b0d",x"381e0e",x"3c2311",x"3b2111",x"371f10",x"351f10",x"331e0f",x"2f1b0e",x"2d1b0e",x"2d1a0f",x"2c1a0f",x"2d1b0e",x"2e1b0f",x"2a180c",x"2c1a0c",x"2e1a0d",x"2f1b0d",x"2f1c0d",x"2f1c0d",x"2e1a0b",x"2c190b",x"2e1a0b",x"29170a",x"2a180a",x"2c190b",x"2b180b",x"2c190b",x"2c190b",x"301b0c",x"321c0c",x"331c0d",x"341d0d",x"39200f",x"361e0e",x"341d0d",x"311c0c",x"351f0e",x"371f0e",x"3a210f",x"39200f",x"38200e",x"381f0e",x"38200e",x"39200f",x"39200e",x"3a210f",x"371f0e",x"341d0d",x"351d0d",x"39200e",x"3b200e",x"3d220f",x"3f2310",x"3e220f",x"3c210f",x"3b210e",x"3a200e",x"391f0e",x"361d0c",x"341c0c",x"331c0c",x"331b0c",x"351d0c",x"39200e",x"3a210f",x"381f0d",x"39200e",x"371e0d",x"361e0d",x"361e0d",x"361e0d",x"381f0e",x"39200e",x"351d0d",x"341c0c",x"341d0d",x"351d0d",x"331b0b",x"331a0b",x"351d0c",x"341d0c",x"341d0c",x"331c0d",x"331d0d",x"2f190b",x"2c180a",x"29170a",x"251509",x"231409",x"2a180b",x"2f1a0c",x"311b0c",x"321c0c",x"2f1a0b",x"2f1a0b",x"2c180a",x"2c190b",x"2e1a0b",x"241509",x"231509",x"231509",x"221409",x"201308",x"1f1308",x"1f1208",x"201308",x"211409",x"211308",x"231409",x"231409",x"241409",x"251509",x"251409",x"251409",x"241409",x"241409",x"241509",x"241509",x"231509",x"221409",x"201308",x"1d1108",x"1a1008",x"190f07",x"1a1008",x"1a1008",x"190f08",x"170f07",x"150e07",x"3e2412",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"221c15",x"231c15",x"201913",x"211b14",x"201a13",x"1f1912",x"1f1812",x"1d1610",x"1b140d",x"171009",x"150e07",x"594e43",x"574d42",x"564b41",x"4a3f35",x"41362b",x"41342a",x"413226",x"433226",x"463426",x"4c3727",x"493424",x"463425",x"473527",x"443225",x"443325",x"423126",x"453327",x"473527",x"473528",x"493629",x"4a3629",x"463426",x"433022",x"463326",x"463223",x"493628",x"493627",x"513a29",x"563d29",x"553e2c",x"58412f",x"563f2d",x"523b2a",x"503a2a",x"513a28",x"563d28",x"523b28",x"4e3928",x"4f3927",x"4a3526",x"4e3928",x"503926",x"4d3726",x"4e3826",x"4c3624",x"4f3724",x"4d3725",x"4f3827",x"453121",x"473222",x"4a3525",x"4b3421",x"473121",x"453022",x"453021",x"453020",x"493322",x"4a3424",x"473120",x"4a3321",x"4a3323",x"4b3420",x"483220",x"47301e",x"4c3422",x"4c3422",x"4d3521",x"473221",x"4c3521",x"483422",x"453123",x"483221",x"4b3320",x"463120",x"4b3422",x"4a3320",x"4b331f",x"47301f",x"4a3321",x"4a3320",x"4b3420",x"493322",x"473123",x"483222",x"4b3524",x"4b3626",x"4d3727",x"523b29",x"523a27",x"513925",x"553b27",x"543b28",x"553b27",x"553c27",x"543c29",x"503a29",x"503929",x"4b3626",x"503929",x"4c3727",x"4e3827",x"4b3728",x"4f3827",x"553c28",x"503928",x"533b28",x"523925",x"4e3722",x"4d3827",x"493424",x"473425",x"483627",x"4d3825",x"453322",x"423121",x"3f3022",x"433121",x"4b3724",x"4b3725",x"493a2d",x"4c4035",x"4c4138",x"4c4238",x"4c4238",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"402410",x"402410",x"432712",x"29180b",x"3b2210",x"412411",x"170f07",x"2b190b",x"2e1a0b",x"2c190b",x"26160a",x"29180b",x"201309",x"2a180b",x"24150a",x"1d1108",x"150e07",x"150e07",x"361e0d",x"150e07",x"462712",x"201309",x"150e07",x"191008",x"150e07",x"150e07",x"150e07",x"543117",x"150e07",x"29180b",x"2d1a0c",x"29180b",x"2a180b",x"150e07",x"150e07",x"492912",x"1f1208",x"150e07",x"1c1108",x"150e07",x"150e07",x"29180b",x"361f0e",x"472913",x"301b0c",x"24150a",x"26160a",x"2d1a0c",x"2c190b",x"2a180b",x"1f1208",x"150e07",x"150e07",x"150e07",x"2d1a0c",x"241509",x"29170a",x"251509",x"221409",x"150e07",x"150e07",x"150e07",x"402510",x"341d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a200e",x"25160a",x"211409",x"150e07",x"150e07",x"351d0e",x"37200f",x"3a2110",x"271c15",x"332c24",x"362f27",x"342d25",x"352d26",x"362e26",x"382e26",x"372d24",x"3a2f27",x"392f27",x"362c24",x"3e352c",x"3b3229",x"3a3028",x"362e26",x"393129",x"383129",x"383028",x"362e27",x"1d160f",x"1d1710",x"1d160f",x"1c160f",x"1c150e",x"1c150e",x"1e150e",x"1d150d",x"1d140d",x"1d140d",x"1b140c",x"1a130c",x"19120c",x"19130c",x"19130c",x"19130c",x"19120b",x"19120b",x"19120c",x"19130c",x"1a130c",x"1f160f",x"241910",x"291c12",x"2e1e14",x"2d1f14",x"2a1e16",x"251c15",x"241d17",x"221b14",x"241e17",x"221c15",x"241d16",x"221b13",x"271d15",x"2b1f16",x"2f2015",x"302116",x"291d14",x"20170f",x"1d160f",x"1b150e",x"1b150e",x"1b150e",x"27190e",x"3c210f",x"29180b",x"26160a",x"231509",x"231509",x"23150a",x"26160a",x"26160a",x"27170a",x"27170a",x"29180b",x"2a180b",x"27160a",x"27160a",x"231509",x"221409",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1c1108",x"190f08",x"1a1008",x"1a1008",x"1b1108",x"1e1208",x"201309",x"211309",x"221409",x"241509",x"27160a",x"27160a",x"261509",x"25150a",x"231409",x"211309",x"201308",x"211309",x"211309",x"201309",x"201309",x"201309",x"221409",x"221309",x"221409",x"231409",x"241509",x"261509",x"251509",x"241308",x"231308",x"231409",x"241509",x"241409",x"231409",x"231409",x"211309",x"1e1208",x"1b1108",x"1a1008",x"1b1108",x"1b1108",x"1a1008",x"170f07",x"26160a",x"3d2311",x"3d2311",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221c15",x"221c15",x"221b14",x"201913",x"201913",x"201a13",x"211b14",x"1f1812",x"1f1811",x"1d160f",x"1b140d",x"171009",x"150e07",x"594f44",x"584e43",x"594d41",x"4d4136",x"4d3f34",x"45372c",x"45362a",x"443327",x"4f3a29",x"503b2a",x"493627",x"4a3628",x"4d392a",x"493629",x"473528",x"4a3628",x"4f3a2a",x"4e392a",x"4c392b",x"4d3a2d",x"513c2f",x"4e3a2b",x"483427",x"523c2b",x"543e2d",x"533d2c",x"533c2c",x"533c2b",x"513927",x"503c2c",x"513c2d",x"513c2d",x"533e2e",x"503a29",x"523b29",x"533c29",x"4e3927",x"4e3a29",x"503a29",x"503a28",x"4f3927",x"513927",x"503926",x"503928",x"4c3727",x"493527",x"4c3626",x"4f3827",x"493525",x"483323",x"493423",x"483324",x"483424",x"4a3524",x"4a3526",x"4b3525",x"4a3525",x"503a27",x"503827",x"4b3524",x"4b3624",x"493424",x"483222",x"483323",x"4a3422",x"493423",x"493423",x"473424",x"493524",x"473323",x"483423",x"473221",x"483525",x"463222",x"473323",x"453021",x"493321",x"483221",x"4a3220",x"4b3422",x"513823",x"493322",x"483323",x"4b3422",x"4b3524",x"4b3626",x"513a28",x"533b28",x"543c28",x"563d28",x"553b26",x"553b27",x"553c29",x"583f2b",x"59412e",x"573e2b",x"573f2d",x"59402d",x"543f2e",x"553f2e",x"533d2e",x"513b2d",x"523c2c",x"523c2c",x"533d2d",x"513c2c",x"543e2c",x"4f3b2b",x"4e3a2c",x"4a3728",x"4f3b2b",x"4a3829",x"4d392a",x"503c2a",x"423326",x"413123",x"493727",x"483626",x"4e3c2d",x"534234",x"50453b",x"52473d",x"53493f",x"53493f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"432712",x"432712",x"442712",x"341d0d",x"39200f",x"422510",x"1f1208",x"2d1a0b",x"321c0c",x"301b0c",x"2c190b",x"2f1b0c",x"301b0c",x"2d190b",x"29180a",x"201309",x"1f1309",x"150e07",x"150e07",x"371f0e",x"301b0c",x"2a180b",x"2c190b",x"2b180b",x"29180b",x"1d1208",x"150e07",x"150e07",x"321c0d",x"331d0d",x"1e1208",x"27170a",x"1f1309",x"150e07",x"4e2b14",x"231409",x"221409",x"29180b",x"2c190b",x"2b190b",x"150e07",x"150e07",x"331c0d",x"2f1a0b",x"241509",x"412511",x"2b180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a1f0d",x"1b1008",x"391e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2a170a",x"3c210e",x"180f07",x"1d1108",x"27160a",x"29170a",x"211309",x"150e07",x"150e07",x"150e07",x"251509",x"1f1309",x"150e07",x"150e07",x"150e07",x"281a11",x"1d160f",x"1e1711",x"1f1912",x"1f1912",x"1f1811",x"201912",x"231a11",x"271b12",x"281c13",x"271b13",x"271a13",x"291b11",x"2d1d12",x"2f1d12",x"2f1f13",x"2b1c11",x"271910",x"22170f",x"1f170f",x"1e170f",x"201710",x"221810",x"251910",x"2a1a10",x"2e1c10",x"321e11",x"331e10",x"331f11",x"2f1d10",x"2b1b0f",x"23160c",x"1f150d",x"1c140c",x"1a130c",x"1a130c",x"19120c",x"19130c",x"19120b",x"1a130c",x"1e140c",x"24180f",x"28190f",x"2e1d13",x"2f1e14",x"2d1e14",x"2c1e14",x"281e16",x"231c15",x"231c16",x"241d16",x"241e17",x"231c16",x"221b14",x"241c15",x"291e15",x"2d1f15",x"312016",x"2d1e13",x"281c12",x"1e150e",x"1c160f",x"1c150e",x"1b150e",x"402614",x"4c2c17",x"2b190b",x"2a180b",x"28170a",x"27160a",x"28170a",x"2a180b",x"2d190b",x"2e1a0c",x"2d190b",x"2d190b",x"2d190b",x"2d190b",x"2b180b",x"241509",x"201308",x"1d1108",x"1e1208",x"211309",x"221409",x"211309",x"201208",x"1e1208",x"1d1108",x"1b1008",x"1a1008",x"1b1108",x"1e1208",x"201309",x"221409",x"231409",x"251509",x"251509",x"221409",x"1d1108",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"180f07",x"1a1008",x"1c1108",x"1d1208",x"1e1208",x"1f1208",x"201208",x"231308",x"251409",x"281609",x"28160a",x"29170a",x"27160a",x"251509",x"251509",x"241409",x"211308",x"201208",x"1f1208",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"180f07",x"3f2411",x"3f2411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221b15",x"221b15",x"221b14",x"201913",x"201a13",x"201912",x"201a13",x"1f1811",x"1e1711",x"1d1710",x"1b140e",x"171009",x"150e07",x"584c41",x"5a4f44",x"54493d",x"55493e",x"4e4034",x"493c31",x"4a3b2e",x"4b3c31",x"4e3d31",x"503e30",x"4d3c2f",x"4f3d2e",x"4e3c2e",x"4c382a",x"49362a",x"47362a",x"4f3d2f",x"4e3d30",x"534134",x"554336",x"554236",x"4f3d31",x"503e31",x"523f30",x"544132",x"533f30",x"513d2e",x"523c2c",x"503928",x"4f3a29",x"523d2d",x"523c2d",x"4f3a29",x"503a2a",x"513c2c",x"4e3927",x"4d3927",x"4d3a2a",x"4b3827",x"4b3625",x"4d3826",x"4c3624",x"4c3726",x"4b3625",x"4b3625",x"483425",x"493423",x"463222",x"443225",x"433225",x"453325",x"493525",x"453224",x"483424",x"493424",x"443122",x"493524",x"493627",x"493628",x"473527",x"493626",x"483524",x"483526",x"473425",x"473425",x"483626",x"4b392a",x"483727",x"493729",x"453527",x"433122",x"483628",x"483524",x"443224",x"443225",x"453427",x"433022",x"433124",x"432f20",x"433022",x"493423",x"463224",x"473222",x"453222",x"483426",x"473426",x"503a29",x"513a29",x"523b2a",x"513a29",x"573e2b",x"563e2c",x"553e2c",x"563e2b",x"563f2d",x"5b4534",x"5a4332",x"574130",x"574334",x"554132",x"544132",x"533e30",x"574436",x"544133",x"544234",x"544235",x"524032",x"534133",x"514032",x"524134",x"524135",x"4d3e31",x"4c3d30",x"493a2d",x"4b3e32",x"483a2e",x"4a3c2e",x"4d3d2f",x"4b3d32",x"4d4236",x"4b4036",x"564b40",x"52483e",x"52483e",x"4c2f1b",x"492914",x"4e301b",x"492a14",x"4a2a14",x"4c2e1a",x"4a3120",x"4d3424",x"482913",x"4c311f",x"483121",x"412511",x"4e311e",x"4d321f",x"4a301f",x"4b3222",x"452712",x"4b301e",x"3f2310",x"402410",x"452b18",x"452812",x"452712",x"482d1b",x"442712",x"422511",x"472c1b",x"432611",x"5f4c3f",x"614c3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3c210f",x"3c210f",x"3e2411",x"331d0d",x"3c2310",x"472812",x"2a180b",x"2e190b",x"2e1a0b",x"301b0b",x"2d190b",x"29170a",x"321c0c",x"2b180b",x"2e1a0b",x"27160a",x"1e1208",x"1e1208",x"150e07",x"150e07",x"2b180a",x"27160a",x"2c190b",x"29170a",x"2d190b",x"27160a",x"1c1108",x"150e07",x"150e07",x"4c2b13",x"2e1a0c",x"150e07",x"150e07",x"25160a",x"321c0c",x"221409",x"2a170a",x"28170a",x"2a170a",x"241409",x"241409",x"150e07",x"150e07",x"1d1108",x"231409",x"1c1108",x"150e07",x"472812",x"3e2310",x"2c190b",x"311b0c",x"361d0d",x"2e190b",x"2f1a0b",x"311b0c",x"371e0d",x"231309",x"211309",x"2a180a",x"39200e",x"432611",x"231509",x"211309",x"28160a",x"2f1b0c",x"2b180b",x"1c1108",x"150e07",x"341c0c",x"150e07",x"29180b",x"1d1108",x"150e07",x"150e07",x"150e07",x"402412",x"331f12",x"241911",x"22170f",x"261b12",x"271a12",x"291c11",x"291b11",x"291b10",x"2e1c12",x"2d1c11",x"301e12",x"321f13",x"331f12",x"362013",x"341f12",x"332013",x"332013",x"2f1d12",x"301e12",x"332013",x"331f11",x"341f11",x"341f11",x"372012",x"3b2112",x"3b2011",x"432713",x"452814",x"3e2311",x"382010",x"321c0e",x"2c1b0f",x"29190e",x"27180c",x"26170c",x"27170d",x"2b190c",x"2a190c",x"2c1b0f",x"2d1b0f",x"2d1b0f",x"2e1d11",x"2f1e13",x"301d12",x"312014",x"301f14",x"2d1e14",x"302118",x"2f2015",x"322217",x"302016",x"322317",x"2f2016",x"312015",x"332115",x"342116",x"3a2417",x"362214",x"332013",x"311f13",x"2d1c10",x"271910",x"2a1a0f",x"2b1a0e",x"462813",x"311a0b",x"2f190b",x"2e190b",x"301a0b",x"331c0c",x"321b0b",x"341c0c",x"371e0d",x"381f0e",x"3c2310",x"3c2310",x"3a200e",x"361d0d",x"2c180a",x"2d190b",x"2e1a0b",x"2e1a0b",x"28160a",x"29160a",x"2e190b",x"2a180a",x"2f1b0c",x"321c0d",x"311b0c",x"29170a",x"2a180a",x"2f1b0c",x"321c0d",x"2f1a0c",x"301b0c",x"2e190b",x"291609",x"2a170a",x"28170a",x"251509",x"271609",x"2a180a",x"261609",x"261609",x"26150a",x"231409",x"221409",x"26160a",x"27160a",x"251509",x"281609",x"2a190c",x"2e1a0c",x"2e1a0c",x"2e1a0c",x"301b0d",x"331c0d",x"351d0e",x"341d0e",x"301b0d",x"311c0d",x"331c0e",x"321c0d",x"2d190b",x"2c190b",x"2c180a",x"2d190b",x"29170a",x"2a180a",x"492a15",x"492a15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231c15",x"231c15",x"231c15",x"211a14",x"201a13",x"211b15",x"201a13",x"1f1912",x"1e1710",x"1c160f",x"1b140d",x"17110a",x"150e07",x"564b40",x"574b41",x"544a3f",x"52473c",x"54473c",x"4f4338",x"514338",x"524439",x"514136",x"58493c",x"564639",x"574638",x"58473a",x"534133",x"4d3d31",x"503e31",x"523f31",x"544133",x"544234",x"524135",x"544335",x"544234",x"584536",x"594536",x"594435",x"544133",x"513d2e",x"533e2d",x"553f2f",x"554031",x"533d2d",x"533e2e",x"4c3829",x"4f3b2b",x"503b2b",x"4b3625",x"4e3a2a",x"4c3726",x"4e3a29",x"503c2c",x"4c3725",x"4e3927",x"4d3826",x"4b3524",x"4a3727",x"443222",x"453223",x"483423",x"453326",x"453223",x"453324",x"453324",x"463325",x"463424",x"443121",x"463325",x"463325",x"463425",x"473525",x"4b3929",x"4a3727",x"4a392c",x"4e3b2b",x"4b3829",x"4c3a2a",x"4d3a2b",x"493829",x"49382b",x"473628",x"4a382a",x"463629",x"4a382b",x"493728",x"473528",x"4d3a2b",x"4d3929",x"4a3829",x"4b3628",x"4c3828",x"4c382a",x"4c392b",x"483426",x"4a3526",x"48362a",x"48372a",x"4c382b",x"4f3b2d",x"533f30",x"533d2c",x"584130",x"584230",x"594331",x"56402f",x"5b4534",x"594433",x"5c4737",x"5a4636",x"5b4637",x"5a4536",x"5a4536",x"574335",x"584639",x"574539",x"574538",x"57473a",x"584739",x"54463b",x"58483c",x"54463a",x"57493c",x"55473c",x"56483c",x"504237",x"54473c",x"54473c",x"53473d",x"4c4136",x"473c31",x"4a3e33",x"4c4138",x"4f453b",x"554b41",x"53493f",x"50311c",x"4c2f1b",x"492914",x"4e301b",x"492a14",x"4a2a14",x"4c2e1a",x"4a3120",x"4d3424",x"482913",x"4c311f",x"483121",x"412511",x"4e311e",x"4d321f",x"4a301f",x"4b3222",x"452712",x"4b301e",x"4d311f",x"402410",x"452b18",x"452812",x"452712",x"482d1b",x"442712",x"422511",x"472c1b",x"432611",x"5f4c3f",x"614c3f",x"614c3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3f2310",x"3f2310",x"402511",x"331d0d",x"39210f",x"3c210f",x"29180a",x"301b0c",x"2f1a0c",x"2f1a0b",x"231409",x"2e1a0c",x"2e1a0c",x"301b0c",x"2b180b",x"26160a",x"221409",x"150e07",x"150e07",x"482712",x"2c190b",x"27170a",x"2c190b",x"2c190b",x"25160a",x"1d1108",x"150e07",x"150e07",x"4d2c14",x"150e07",x"432712",x"1c1108",x"150e07",x"3a210f",x"311c0c",x"2f1b0c",x"2f1a0b",x"301b0c",x"2e1a0b",x"2d190b",x"2a170a",x"251509",x"1e1208",x"150e07",x"150e07",x"150e07",x"351d0c",x"150e07",x"150e07",x"150e07",x"3d210e",x"3a200d",x"3f2310",x"3c210f",x"3f230f",x"3f2310",x"311c0d",x"150e07",x"2e1a0b",x"231409",x"391f0d",x"170f07",x"28170a",x"2c190b",x"2b180b",x"231409",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"150e07",x"150e07",x"311d0e",x"2e1a0b",x"1c1108",x"1a1008",x"1c1108",x"1d1108",x"201208",x"241509",x"241509",x"28170a",x"2c180b",x"311b0b",x"361e0d",x"361e0d",x"341d0c",x"321c0c",x"311b0c",x"301a0b",x"341d0c",x"351d0c",x"341c0c",x"341c0c",x"351c0c",x"371e0d",x"381f0d",x"371e0d",x"381e0d",x"3c210e",x"3f230f",x"3a200e",x"341c0c",x"301a0b",x"2f1a0b",x"2e1a0b",x"2e1a0c",x"2c190b",x"2b180b",x"2c190b",x"2c190b",x"2a180b",x"27160a",x"27160a",x"25150a",x"26160a",x"251509",x"27160a",x"251509",x"241409",x"231409",x"241509",x"241509",x"241509",x"231509",x"231409",x"231409",x"26160a",x"2a180b",x"2e1b0c",x"301c0d",x"2d1a0c",x"28170b",x"25150a",x"221409",x"1d1108",x"1f1208",x"432611",x"241509",x"26160a",x"28160a",x"29170a",x"2c180b",x"2b180a",x"2b180a",x"2b180a",x"2b180a",x"301b0c",x"321c0c",x"301b0c",x"2d190b",x"2b180b",x"28170a",x"25150a",x"28170b",x"2a180b",x"2b190b",x"2a180b",x"261509",x"27160a",x"251509",x"251509",x"251509",x"241509",x"26160a",x"29180b",x"2b180b",x"2b180b",x"29170a",x"251509",x"27160a",x"231409",x"1e1108",x"1e1208",x"221409",x"231409",x"201208",x"1f130a",x"1c120a",x"1f140d",x"21170f",x"241910",x"281b12",x"2c1f16",x"2e2015",x"312117",x"362418",x"362418",x"372519",x"362418",x"352417",x"352318",x"352418",x"352419",x"332217",x"2f2016",x"2d1f16",x"2c1f16",x"2a1d13",x"271b12",x"251b13",x"2a1c11",x"4e2e18",x"4e2e18",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221c15",x"221c15",x"201912",x"211a14",x"201a13",x"201a13",x"201a13",x"1f1811",x"1f1812",x"1d160f",x"1b150e",x"171009",x"150e07",x"53483e",x"53483d",x"51453a",x"55493f",x"55493e",x"52453a",x"54473c",x"39200e",x"3d200d",x"3b210d",x"3c210e",x"3e2310",x"3f2310",x"3f230f",x"3c210e",x"3f2310",x"3e220f",x"422511",x"432611",x"432611",x"482912",x"3f230f",x"40220f",x"40230f",x"331b0b",x"412410",x"452611",x"442611",x"442611",x"462711",x"432511",x"3f230f",x"391e0c",x"42240f",x"442711",x"422510",x"40230f",x"40230f",x"3e230f",x"3a200d",x"381d0c",x"361d0c",x"3d210f",x"3b200d",x"3c200e",x"432510",x"3b200d",x"3d210e",x"3e220e",x"3f230f",x"422510",x"3e220f",x"3c210e",x"402310",x"3b200e",x"381e0c",x"3c210e",x"3d210e",x"3c210e",x"3b200d",x"3b200d",x"3d220e",x"3e220f",x"3d210e",x"3a1f0d",x"3d220e",x"3f2310",x"3d220f",x"3c200e",x"3a1f0d",x"3d210f",x"422511",x"452711",x"462711",x"442611",x"4a2a13",x"492912",x"4c3a2d",x"4c3a2c",x"4a392d",x"422b1c",x"665143",x"614d3f",x"634f42",x"634f42",x"614e41",x"624e41",x"634f41",x"5e4a3c",x"614c3e",x"604a3b",x"614d3f",x"604d40",x"614e40",x"605043",x"655041",x"614d3f",x"654f40",x"655142",x"624e3f",x"655143",x"5d4b3d",x"5d4a3d",x"5f4d3f",x"5e4c40",x"5c4b3d",x"5e4d41",x"5e4e41",x"5c4b3f",x"5d4d40",x"5c4c40",x"5a4b3f",x"5b4b3f",x"5b4b3e",x"5e4d3f",x"604f42",x"59483a",x"604c3f",x"604f43",x"5c4b3d",x"604c3e",x"604d3f",x"624f41",x"5d4b3d",x"58473a",x"5b493b",x"5e4d40",x"5f4e42",x"5d4b3d",x"5b483a",x"615043",x"625043",x"624f41",x"5e4b3e",x"5c4c40",x"5c4d41",x"5e4c3f",x"5b493c",x"5a4b3e",x"5a4a3d",x"5b4a3c",x"5c4a3d",x"59483c",x"5a4b40",x"5c4b3e",x"59493c",x"5a483c",x"5e4d40",x"5c4b3f",x"5a4a3e",x"5d4d40",x"5b4b3f",x"5f4e41",x"543624",x"543624",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"452914",x"452914",x"432612",x"311c0d",x"361e0d",x"3b200e",x"1c1008",x"27160a",x"29170a",x"2d1a0b",x"231409",x"1e1208",x"28170a",x"28170a",x"25150a",x"231509",x"150e07",x"150e07",x"412410",x"150e07",x"3c220f",x"150e07",x"150e07",x"1b1108",x"150e07",x"150e07",x"150e07",x"462712",x"150e07",x"150e07",x"150e07",x"4b2b14",x"150e07",x"150e07",x"29170a",x"28160a",x"2f1a0b",x"2d190b",x"2e1a0b",x"2f1a0c",x"2f1b0c",x"2b180b",x"2b180a",x"261509",x"1d1108",x"150e07",x"351d0d",x"27160a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3c210e",x"351e0d",x"341d0d",x"402410",x"29170a",x"2a180b",x"29170a",x"25150a",x"191008",x"150e07",x"3e2310",x"301c0d",x"150e07",x"2d190b",x"1f1309",x"150e07",x"150e07",x"150e07",x"351e0d",x"25150a",x"1e1108",x"1a1008",x"180f08",x"191008",x"1c1108",x"1c1108",x"1d1108",x"211309",x"231409",x"281609",x"2d190b",x"301b0b",x"301a0b",x"2e1a0b",x"2d190b",x"2e190b",x"331c0c",x"341d0d",x"341d0c",x"331c0c",x"331c0c",x"351d0d",x"361e0d",x"39200e",x"3a200e",x"3c210e",x"381e0d",x"39200e",x"361e0d",x"351d0d",x"301a0b",x"281609",x"28160a",x"2b180b",x"2a180b",x"29180b",x"28170a",x"26160a",x"241509",x"221409",x"231409",x"231409",x"221409",x"1f1208",x"1c1108",x"1c1108",x"1d1108",x"1c1108",x"1b1108",x"1b1108",x"1b1008",x"1a1008",x"1a1008",x"1c1108",x"1f1208",x"1f1208",x"1d1108",x"1d1208",x"1f1208",x"1d1108",x"1b1108",x"191008",x"170f07",x"150e07",x"1e1208",x"221409",x"27160a",x"27160a",x"251509",x"27160a",x"2a180a",x"2d1a0b",x"2d1a0b",x"2b180a",x"2b180a",x"2d190b",x"2d190b",x"2c190b",x"27160a",x"211309",x"1f1309",x"221409",x"251509",x"241509",x"251509",x"26160a",x"27160a",x"26160a",x"231509",x"1e1208",x"1a1008",x"1a1008",x"1c1108",x"1c1108",x"1a1008",x"180f08",x"160e07",x"150e07",x"160e07",x"191008",x"1e1208",x"1f1208",x"21140c",x"1d120b",x"1a140c",x"1c150e",x"1f170f",x"221a13",x"211a12",x"241c15",x"261d16",x"281e16",x"2c2118",x"2e2219",x"302219",x"30231a",x"2f2218",x"2f2218",x"312219",x"312319",x"312319",x"2f2219",x"302319",x"2d2117",x"2d2118",x"2a1e16",x"261c14",x"3a2416",x"4d2e17",x"301d12",x"2f1d11",x"321f12",x"352113",x"342114",x"362214",x"301e13",x"332013",x"312013",x"2f1f12",x"2c1c10",x"281a0f",x"26180e",x"25170d",x"21150c",x"1c130b",x"462814",x"462814",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"231c16",x"211a13",x"201912",x"201a13",x"201913",x"1e1710",x"1f1912",x"1d1710",x"1b150e",x"171009",x"150e07",x"150e07",x"53483d",x"51453a",x"55493f",x"55493e",x"3c230f",x"3f2411",x"301b0d",x"2f1a0b",x"38200d",x"311b0c",x"29170a",x"2f1a0b",x"2d190b",x"311b0c",x"301a0b",x"311c0c",x"2f1b0c",x"301b0c",x"2e1a0b",x"311b0c",x"2e1a0b",x"2e1a0b",x"321c0c",x"2f1b0c",x"28170a",x"311b0c",x"311c0c",x"311c0c",x"301b0c",x"27160a",x"311c0d",x"321c0d",x"331e0e",x"301c0d",x"2f1c0c",x"301c0c",x"311c0c",x"28160a",x"2d190b",x"2f1b0c",x"37200f",x"321c0d",x"301b0c",x"311c0d",x"2f1a0b",x"2a170a",x"29170a",x"251509",x"251509",x"2b180b",x"2b180a",x"29170a",x"2d190b",x"2b180a",x"2b180a",x"2f1a0b",x"2f1a0b",x"2d190b",x"2f1a0b",x"2c180b",x"2e190b",x"2e1a0b",x"2f1a0b",x"2d190b",x"2b180a",x"2c180a",x"301a0b",x"311b0c",x"331c0d",x"311b0c",x"281609",x"2d190b",x"361e0d",x"341d0d",x"341d0d",x"3b200e",x"2b190c",x"321d0d",x"38271b",x"38271b",x"634f41",x"584a3e",x"5b4b3f",x"5d4d41",x"5b4b3f",x"5e4f43",x"55483d",x"54463a",x"58493d",x"57483b",x"57483c",x"58483d",x"57493e",x"57493e",x"594a3e",x"584a3f",x"5a4c40",x"5b4c40",x"56483e",x"594a3f",x"574a3e",x"584a3f",x"5a4c41",x"5a4c40",x"5d4e42",x"584a3e",x"57493e",x"53463b",x"55483d",x"594c41",x"54473c",x"584a40",x"55493f",x"574b41",x"524439",x"594d42",x"57493e",x"584a3e",x"5a4c40",x"57483c",x"5a4c41",x"584a3f",x"584b40",x"57483c",x"56463a",x"584a3e",x"55473a",x"584a3e",x"5d4e42",x"57473b",x"594a3e",x"594b3f",x"5a4a3e",x"5b4b3e",x"5b4b3f",x"5c4c40",x"56473a",x"56483c",x"5b4c41",x"594b3f",x"56483c",x"55483d",x"594b3f",x"58493d",x"5a4c40",x"57473c",x"5b4e42",x"54473c",x"54463b",x"4e4338",x"5c4b3e",x"5c4c3f",x"533929",x"533929",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"442813",x"442813",x"3f2411",x"341d0d",x"351d0d",x"351d0d",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"351d0d",x"311b0b",x"150e07",x"251509",x"2e1a0b",x"150e07",x"150e07",x"1a1008",x"4a2913",x"2d190b",x"150e07",x"26160a",x"201309",x"150e07",x"28170a",x"3f2310",x"2c190b",x"39200e",x"231409",x"2b190b",x"2b180b",x"2c190b",x"2f1b0c",x"331c0d",x"2d190b",x"301b0c",x"28170a",x"27160a",x"150e07",x"150e07",x"442712",x"27160a",x"26160a",x"221409",x"201309",x"150e07",x"150e07",x"150e07",x"4d2c15",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"462813",x"150e07",x"150e07",x"231509",x"150e07",x"150e07",x"2d1a0c",x"150e07",x"361e0d",x"150e07",x"2a180b",x"1e1208",x"150e07",x"150e07",x"150e07",x"321c0c",x"38200e",x"321d0d",x"29170a",x"28160a",x"2d190b",x"2b180b",x"2c180b",x"301b0c",x"311c0c",x"311b0c",x"351e0d",x"361d0d",x"381f0d",x"3c210e",x"3b210e",x"3c210e",x"3d210f",x"3c210f",x"3c220f",x"3b200e",x"3b210e",x"3b200e",x"3a200e",x"381f0d",x"371e0c",x"371d0c",x"351d0c",x"3b210e",x"3f230f",x"412410",x"422510",x"3f2310",x"402410",x"381f0d",x"39200e",x"361e0d",x"341e0d",x"331d0d",x"321c0d",x"321c0d",x"311c0d",x"301b0c",x"301c0c",x"311c0c",x"2d190b",x"29170a",x"2c180b",x"2d190b",x"2f1a0b",x"301b0c",x"301b0c",x"2e1a0c",x"26160a",x"26160a",x"27160a",x"29170b",x"2a180b",x"29170a",x"2a170b",x"2a180b",x"2a180b",x"2a170b",x"29170a",x"2a170a",x"2a180a",x"361d0d",x"321c0c",x"2a180a",x"2a170a",x"27160a",x"26190f",x"26190e",x"231409",x"3c2d24",x"3c2e24",x"2b190b",x"2b190b",x"2a180b",x"2b190b",x"2b180b",x"2a180b",x"2b190b",x"2c190b",x"2e1a0c",x"2f1b0c",x"301c0c",x"301b0d",x"2f1b0b",x"2d190b",x"2b180b",x"25150a",x"22140a",x"211409",x"23150a",x"23150a",x"24150a",x"24150a",x"24150a",x"231409",x"211309",x"211309",x"211309",x"221409",x"221409",x"221409",x"22140a",x"24160b",x"25170d",x"24170d",x"25180e",x"251910",x"23180f",x"231910",x"241a11",x"251911",x"271b11",x"281b11",x"281b11",x"261a11",x"261b12",x"271a11",x"271a11",x"271a12",x"271b11",x"271a12",x"251910",x"24190f",x"251a11",x"251910",x"422714",x"301d12",x"2f1d11",x"321f12",x"352113",x"342114",x"362214",x"301e13",x"332013",x"312013",x"2f1f12",x"2c1c10",x"281a0f",x"26180e",x"25170d",x"21150c",x"1c130b",x"462814",x"462814",x"000000",x"000000",x"000000",x"000000",x"000000",x"221c15",x"221c15",x"231c16",x"201912",x"201912",x"201a13",x"201a13",x"1f1912",x"1d1610",x"1d1610",x"1b150e",x"17110a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"3f230f",x"39210e",x"381f0e",x"442810",x"402510",x"3e230f",x"3b210f",x"3b220f",x"371f0e",x"351e0d",x"3f2410",x"39200e",x"361d0d",x"3e230f",x"3d2210",x"3c220f",x"3e2410",x"3b220f",x"3a210f",x"3a210f",x"3e2310",x"3e2310",x"3b220f",x"402512",x"361f0f",x"3e2411",x"341d0d",x"371e0d",x"38200e",x"3a200e",x"38200e",x"37200f",x"351e0d",x"361e0d",x"3c2310",x"3e2411",x"38200e",x"351d0d",x"371f0d",x"3b210e",x"381e0d",x"361e0d",x"3b210f",x"39200e",x"331d0d",x"311c0c",x"2d190b",x"2e1a0b",x"2f1b0b",x"331c0c",x"351d0c",x"351d0d",x"3a200e",x"341d0d",x"341d0d",x"351d0d",x"391f0e",x"381f0d",x"341c0c",x"321b0b",x"321b0b",x"331c0b",x"351d0d",x"361e0d",x"39200e",x"361f0d",x"371f0d",x"361e0e",x"361e0d",x"3b210f",x"3b210f",x"3d2310",x"3e2310",x"422713",x"412612",x"3d291c",x"3d291c",x"635042",x"5a4e44",x"3c2c20",x"2e231a",x"31261d",x"2e241c",x"31271f",x"3b2e25",x"382e26",x"342a22",x"32281e",x"332921",x"2c2118",x"32281f",x"342921",x"382d24",x"362a21",x"382b21",x"352b23",x"32271e",x"2c231b",x"31261d",x"2d221a",x"31271f",x"2f241c",x"382b22",x"3a2e24",x"3d3229",x"3d322a",x"3e3229",x"362b22",x"372c22",x"342d25",x"3e342b",x"362d25",x"2e251d",x"382d24",x"3b2e24",x"3a2d23",x"392d23",x"372a21",x"413328",x"41362d",x"41362d",x"41342a",x"403227",x"403329",x"3f3127",x"392a1f",x"433328",x"423328",x"3b2b20",x"37291f",x"3a2b21",x"3c2f25",x"33251b",x"38281c",x"372519",x"332217",x"2e2015",x"3a2a1f",x"3e2f24",x"372d25",x"403228",x"3e3026",x"3a2b20",x"2f251d",x"38291f",x"3a291d",x"3b2c22",x"3a2c22",x"4b2e1a",x"4b2e1a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"432712",x"432712",x"3f2410",x"311c0d",x"321c0d",x"2e1a0b",x"2b180a",x"341d0d",x"38200e",x"361e0e",x"321c0c",x"2d190b",x"341d0d",x"351f0e",x"311b0c",x"2f1a0b",x"3f230f",x"432611",x"331c0d",x"2d190b",x"321c0c",x"412511",x"422611",x"452712",x"432611",x"462812",x"150e07",x"1d1208",x"27170a",x"1e1208",x"150e07",x"150e07",x"442813",x"2e1b0c",x"442712",x"28170a",x"2f1b0c",x"341d0d",x"2f1a0b",x"2e190b",x"2c180a",x"2b180a",x"261509",x"28160a",x"1e1208",x"150e07",x"150e07",x"442510",x"25150a",x"27170a",x"29170b",x"170f07",x"150e07",x"231409",x"462712",x"1f1309",x"231409",x"29170a",x"2b190b",x"1d1208",x"150e07",x"170f07",x"422510",x"1f1209",x"150e07",x"331c0d",x"201208",x"3c210f",x"341e0d",x"150e07",x"28170a",x"211409",x"150e07",x"150e07",x"150e07",x"331c0c",x"311c0d",x"301b0b",x"29170a",x"221409",x"241409",x"29170a",x"271609",x"2c190b",x"2d190b",x"301b0c",x"351e0e",x"331c0c",x"39200e",x"3a200e",x"3d220f",x"3f2410",x"3e2310",x"3c210f",x"3b210f",x"3b210f",x"3b210e",x"371f0d",x"391f0e",x"381f0d",x"391f0d",x"3a200e",x"3c210f",x"371d0c",x"361d0c",x"3b200e",x"3f230f",x"3f230f",x"3f2310",x"391f0d",x"3a210f",x"371f0e",x"331d0d",x"301b0c",x"2f1a0c",x"311c0c",x"301b0d",x"2a170a",x"2c190b",x"2e1a0c",x"2e1a0b",x"2c190b",x"2f1a0c",x"2f1b0c",x"2f1b0c",x"301b0c",x"2f1b0c",x"2f1b0c",x"311c0d",x"311c0d",x"331d0d",x"341e0e",x"331d0d",x"341e0e",x"331d0d",x"341e0e",x"351e0e",x"361f0e",x"361f0e",x"361e0d",x"351d0d",x"321b0c",x"301b0b",x"2f1a0b",x"2a170a",x"27160a",x"241509",x"1f1208",x"1a1008",x"422612",x"311c0c",x"301b0c",x"311b0c",x"2f1b0c",x"301b0c",x"2f1a0b",x"341d0d",x"371f0e",x"371f0d",x"371e0d",x"38200e",x"3b220f",x"39210f",x"38200f",x"341d0d",x"301b0c",x"2b180b",x"28170a",x"27160a",x"29170a",x"2e1a0c",x"2f1b0c",x"2f1b0c",x"2d1a0c",x"2c1a0b",x"2c190b",x"2b190b",x"2a190b",x"261609",x"27160a",x"251509",x"29170a",x"271609",x"2b180a",x"281709",x"2c190b",x"251509",x"231409",x"211309",x"201309",x"221409",x"241409",x"241509",x"231409",x"201309",x"1c1108",x"1c1108",x"1d1208",x"1f1208",x"20140a",x"23150b",x"25160c",x"28190e",x"2d1b0f",x"321e11",x"301c11",x"2e1c0f",x"311e12",x"332013",x"352013",x"352013",x"301e13",x"352114",x"342011",x"321e11",x"2e1d11",x"2b1a0f",x"291a0f",x"291a0f",x"23150b",x"20140b",x"1a1008",x"422613",x"422613",x"000000",x"000000",x"000000",x"000000",x"000000",x"221c15",x"221c15",x"211a14",x"211a14",x"201913",x"201a13",x"211a14",x"1f1811",x"1d1710",x"1d1710",x"1b150e",x"17110a",x"150e07",x"150e07",x"000000",x"000000",x"4b2d14",x"3f240e",x"3f230f",x"42250f",x"3e230e",x"3f240f",x"3a210e",x"331c0c",x"402510",x"432611",x"3b210f",x"3a210f",x"3c210f",x"3b200e",x"3c220f",x"39200e",x"3a200e",x"381f0e",x"3d2310",x"3a210f",x"3a210f",x"3b200f",x"361e0e",x"3d230f",x"38200e",x"371e0d",x"351d0d",x"381f0e",x"3d2310",x"3e2310",x"38200e",x"38200e",x"38200e",x"3b220f",x"3b210f",x"341d0d",x"39200e",x"331c0b",x"391f0d",x"311b0b",x"351d0c",x"3c210e",x"3a1f0d",x"351d0c",x"361d0d",x"331d0c",x"361f0e",x"301b0c",x"351e0d",x"321c0c",x"361e0d",x"361e0d",x"361f0d",x"321c0d",x"371f0e",x"2f1a0b",x"331c0c",x"321c0c",x"341d0d",x"301a0b",x"351d0d",x"391f0e",x"331c0c",x"321b0b",x"321b0b",x"331c0c",x"39200e",x"361e0d",x"341c0c",x"391f0e",x"3d220f",x"3e2310",x"3d220f",x"422410",x"422511",x"3c210f",x"37261c",x"37261c",x"5d5045",x"5c4c3f",x"614f41",x"5a4c41",x"170f07",x"180f08",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1d1208",x"1d1208",x"1e1209",x"1e1209",x"1e1208",x"1e1209",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"201309",x"211409",x"231409",x"231509",x"231509",x"25160a",x"25150a",x"26160a",x"251509",x"25150a",x"26160a",x"27160a",x"27160a",x"29170b",x"2a180b",x"2a190b",x"341d0d",x"2e1a0b",x"2f1a0b",x"2c190b",x"2c190b",x"2a1a0d",x"291a0d",x"2a1a0d",x"2b1b0d",x"311d0f",x"3d2311",x"3a2211",x"5a4a3e",x"5c4b3e",x"5a4a3d",x"57493d",x"584a3f",x"58473a",x"5a493c",x"58483b",x"58493d",x"57483b",x"55473c",x"58493c",x"57483d",x"54453a",x"56493e",x"574a3e",x"54463b",x"4b3b2f",x"4a3d33",x"4f4035",x"4a3c32",x"473a2f",x"5c4535",x"57351f",x"57351f",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3e2310",x"3e2310",x"412511",x"311c0d",x"39210f",x"39200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"432712",x"150e07",x"3f2511",x"201409",x"150e07",x"150e07",x"150e07",x"150e07",x"4f2d15",x"2a180b",x"150e07",x"150e07",x"150e07",x"442611",x"39200e",x"2f1b0c",x"2b180a",x"271609",x"2f1a0b",x"301a0b",x"2e190b",x"2e1a0b",x"2e190b",x"2d190b",x"2e190b",x"201308",x"1e1208",x"150e07",x"150e07",x"3a200e",x"231409",x"1e1208",x"150e07",x"150e07",x"381f0e",x"3c2310",x"1b1108",x"2e1b0c",x"2f1a0b",x"2e1a0b",x"2a180a",x"2d1a0b",x"1d1208",x"150e07",x"29170a",x"150e07",x"27160a",x"2a180a",x"2e1b0c",x"321c0d",x"2f1b0c",x"150e07",x"2d1a0c",x"211409",x"150e07",x"150e07",x"150e07",x"301b0d",x"321c0e",x"341e0f",x"27170c",x"24160c",x"22150b",x"25170b",x"25160b",x"29170c",x"29190c",x"2d1a0d",x"2e1b0d",x"351e0d",x"371e0d",x"3c220f",x"3f2410",x"3f2410",x"3c210f",x"39200e",x"361e0d",x"351d0c",x"341c0b",x"361d0c",x"39200f",x"3a200f",x"39200f",x"3b210e",x"3c210f",x"3d220f",x"3b210e",x"3f230f",x"422511",x"432611",x"3f230f",x"3d210f",x"39200e",x"311b0b",x"301b0c",x"311c0c",x"2b180a",x"2d190b",x"311d0d",x"311d0d",x"301c0d",x"2f1c0d",x"2e1b0c",x"2c190b",x"2d1c0d",x"2f1d0f",x"301c0e",x"2f1c0e",x"2f1c0e",x"301e10",x"2f1d0f",x"2d1b0f",x"2d1c0f",x"2d1b0f",x"2e1c0f",x"2d1c0e",x"2c1b0f",x"2a190e",x"2c1b0e",x"2c1a0e",x"2e1b0f",x"301d0f",x"2f1a0d",x"2e1b0c",x"2e1a0d",x"2b180c",x"2a190c",x"27180c",x"23150b",x"1c1108",x"180f07",x"402513",x"2e1a0b",x"2d190b",x"2f1a0b",x"321c0d",x"331c0d",x"361f0e",x"3a220f",x"3b2210",x"3a200f",x"381f0e",x"381f0e",x"381f0e",x"3a210f",x"381f0e",x"341d0d",x"2e1a0b",x"29170a",x"29170a",x"2c190b",x"2f1b0c",x"301c0c",x"311c0c",x"301c0c",x"2f1b0c",x"2f1b0c",x"2e1a0b",x"2d190b",x"2a180b",x"29170a",x"29170a",x"2a180a",x"2d190b",x"2c180a",x"2c190a",x"2e1a0b",x"2c180a",x"2a170a",x"251509",x"231409",x"24150a",x"26160a",x"27160a",x"28170b",x"26160a",x"221409",x"1e1208",x"1d1108",x"1c1108",x"1d1108",x"1e1208",x"221409",x"25170b",x"29190c",x"2e1b0d",x"321c0e",x"331d0e",x"311d0d",x"321c0d",x"331d0f",x"351e0f",x"331d0e",x"331d0e",x"321c0e",x"2f1c0d",x"2c1a0c",x"2d1a0d",x"29190d",x"26170b",x"2a1a0d",x"27170b",x"221509",x"1d1108",x"2d1a0c",x"2d1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"211b14",x"211b14",x"201a13",x"201913",x"1f1811",x"201a13",x"211a14",x"1f1912",x"1d160f",x"1d1610",x"1b140d",x"171009",x"150e07",x"150e07",x"000000",x"000000",x"513215",x"4b2d14",x"4d2c12",x"4b2b10",x"43270f",x"3c210e",x"3c220e",x"42260f",x"3c220e",x"391f0d",x"3f2310",x"3e220f",x"3c210f",x"3f2411",x"3e2411",x"3d2310",x"371f0e",x"361e0d",x"361e0d",x"38200e",x"3c210f",x"371f0e",x"331d0d",x"381f0d",x"341d0d",x"39200e",x"38200e",x"361f0e",x"301b0c",x"311c0c",x"351e0d",x"321d0d",x"361f0e",x"371f0e",x"38200e",x"351d0d",x"351e0d",x"351d0c",x"311b0b",x"351d0c",x"351d0c",x"3a200d",x"311a0a",x"331c0b",x"381f0d",x"321c0c",x"351d0d",x"3a210f",x"371f0e",x"38200e",x"3a210f",x"38200e",x"371f0d",x"351e0d",x"2c180a",x"2e190b",x"2e190b",x"321c0c",x"341d0c",x"381f0d",x"321c0c",x"381f0e",x"361e0d",x"321c0c",x"361d0d",x"381f0d",x"3b210f",x"3a200e",x"3a200e",x"3a200e",x"3b210f",x"371d0d",x"3a200e",x"3d220f",x"3a1f0d",x"4b2b14",x"3b210e",x"35281f",x"5c4e42",x"615145",x"5b4c40",x"544a40",x"170f07",x"180f07",x"180f07",x"190f08",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1c1108",x"1b1008",x"1c1108",x"1d1108",x"1e1208",x"1f1208",x"201308",x"211309",x"221409",x"221409",x"221409",x"221409",x"221309",x"241409",x"241509",x"231409",x"25150a",x"27160a",x"27160a",x"29180b",x"2a180b",x"2a180b",x"28170a",x"28170a",x"27160a",x"27160a",x"27160a",x"241509",x"221409",x"201309",x"1f1208",x"1f1208",x"201309",x"211409",x"211309",x"211409",x"211409",x"211409",x"231509",x"25150a",x"27160a",x"27160a",x"28170a",x"261509",x"261509",x"28170a",x"241509",x"221409",x"1e1208",x"1a1008",x"160e07",x"150e07",x"1a1008",x"191008",x"180f07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"402511",x"402511",x"412511",x"2d1a0c",x"351f0e",x"351c0c",x"190f07",x"221409",x"251509",x"261609",x"251509",x"27160a",x"2f1a0c",x"26150a",x"231409",x"201208",x"170f07",x"150e07",x"150e07",x"1c1108",x"271609",x"170f07",x"1e1108",x"211309",x"1d1108",x"150e07",x"150e07",x"150e07",x"3a220f",x"150e07",x"150e07",x"422611",x"150e07",x"422611",x"2d1a0b",x"331d0d",x"331d0d",x"301b0c",x"321c0c",x"2e190b",x"2e190b",x"2c180b",x"29180b",x"1e1208",x"191008",x"150e07",x"371f0e",x"26160a",x"150e07",x"150e07",x"150e07",x"462611",x"26150a",x"221409",x"331d0d",x"311c0c",x"2f1a0b",x"331d0d",x"2e1b0c",x"2a190b",x"150e07",x"150e07",x"412511",x"1d1108",x"3b210f",x"150e07",x"39200e",x"27170a",x"321d0d",x"150e07",x"2b190b",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1c0d",x"2e1c0d",x"28180b",x"21140b",x"1d130a",x"1f130a",x"24160b",x"21150a",x"23160a",x"27170b",x"2e1c0d",x"2d1b0d",x"321c0e",x"381f0f",x"3a2110",x"381f0f",x"361e0f",x"37200f",x"301b0d",x"321c0d",x"331d0e",x"351e0e",x"361e0e",x"371e0e",x"371e0e",x"361e0e",x"351d0d",x"361e0e",x"391f0f",x"371e0e",x"391e0d",x"3a1f0d",x"391e0d",x"39200e",x"351d0c",x"311b0b",x"2f1a0b",x"2f1a0b",x"2d1a0b",x"2c180b",x"2b180a",x"28160a",x"261509",x"29170a",x"29190c",x"26170b",x"26170b",x"25160b",x"26170d",x"29190d",x"29190f",x"29190d",x"2a1a0f",x"2b1b10",x"2d1c11",x"2d1d11",x"2d1d11",x"2d1d11",x"2b1b0f",x"2b1b10",x"2b1b0f",x"2d1d10",x"301e11",x"301d0f",x"311d0f",x"2d1b0f",x"2b1a0e",x"27170b",x"29190c",x"27180c",x"23160b",x"1f130a",x"1a110a",x"2b180b",x"2d190b",x"2e190b",x"311b0c",x"331c0c",x"311b0b",x"341d0d",x"39200f",x"3b210f",x"341c0c",x"39200e",x"3e2411",x"3d2310",x"3c220f",x"3a210f",x"361f0e",x"311c0c",x"2d1a0b",x"2d1a0b",x"301c0c",x"311c0d",x"341e0e",x"331d0d",x"331d0d",x"321c0d",x"2f1b0b",x"2c190b",x"2a180a",x"2c190b",x"29170a",x"2c190b",x"2c190b",x"2c190a",x"2d190a",x"281609",x"2c190a",x"2d190a",x"2c180a",x"27160a",x"27160a",x"251509",x"261509",x"28170a",x"28170a",x"26160a",x"211309",x"1e1208",x"1c1108",x"1c1108",x"1d1108",x"1f1208",x"221409",x"241409",x"27160a",x"2b180a",x"2c180a",x"2d190a",x"2f1a0b",x"2d190a",x"2d180a",x"2d190a",x"2d190a",x"2e190b",x"2f1a0b",x"2d180a",x"2c190b",x"2b180b",x"29180a",x"28170a",x"26160a",x"231409",x"1e1208",x"1b1108",x"372010",x"372010",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"1f1912",x"211a14",x"201a13",x"1f1811",x"1f1812",x"1f1912",x"1d160f",x"1d1710",x"1b150e",x"17110a",x"150e07",x"150e07",x"000000",x"563416",x"59361a",x"523215",x"4f3015",x"533314",x"4b2e14",x"472b12",x"412711",x"412710",x"3e2410",x"3d220f",x"3f2411",x"3c2110",x"39200f",x"3b2111",x"3a2111",x"341d0e",x"351d0e",x"3a2110",x"3b2211",x"3b2311",x"3f2412",x"3b2211",x"382110",x"3e2312",x"361f0f",x"351f0f",x"351f0f",x"372010",x"372010",x"382110",x"38200f",x"382010",x"351e0f",x"311c0d",x"361e0f",x"392010",x"371f0f",x"321c0d",x"301b0d",x"351e0e",x"2d1a0c",x"301b0c",x"3a200f",x"341d0b",x"381f0c",x"301a0b",x"371f0d",x"321c0c",x"351d0d",x"361e0d",x"371f0d",x"351e0d",x"331d0c",x"341d0c",x"2a170a",x"2e190a",x"301a0b",x"331c0c",x"2e190b",x"321c0c",x"311b0b",x"341c0c",x"301a0b",x"311b0b",x"361d0c",x"321b0b",x"341c0c",x"351d0c",x"351d0c",x"361e0d",x"381e0d",x"351d0c",x"3a200e",x"3d220f",x"3e230f",x"3f230f",x"472813",x"644e3e",x"655041",x"150e07",x"4d4339",x"554b41",x"160e07",x"160e07",x"160e07",x"2b1a0a",x"231609",x"1d1108",x"1f1308",x"1d1208",x"1f1209",x"221409",x"24160a",x"26160a",x"27170a",x"28170a",x"28170a",x"27170a",x"25160a",x"241509",x"231409",x"201308",x"1f1208",x"201208",x"221409",x"221409",x"211409",x"201309",x"1e1208",x"1b1008",x"190f08",x"180f07",x"191008",x"1a1008",x"1a1008",x"1c1108",x"1d1208",x"1d1208",x"1d1108",x"201309",x"23150a",x"241509",x"25160a",x"25160a",x"25160a",x"25150a",x"241509",x"24150a",x"25160a",x"25150a",x"25160a",x"25150a",x"24150a",x"231409",x"201309",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1e1208",x"1f1208",x"1f1208",x"1e1108",x"1c1108",x"1e1208",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"180f07",x"170f07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"432612",x"432612",x"412511",x"301b0c",x"3a220f",x"3c210e",x"1d1108",x"2d190b",x"2b180b",x"251509",x"27160a",x"27160a",x"2b180b",x"29170a",x"27160a",x"211309",x"251509",x"190f07",x"150e07",x"150e07",x"201208",x"211208",x"241409",x"211309",x"261509",x"221409",x"150e07",x"150e07",x"150e07",x"26160a",x"472712",x"2c190b",x"150e07",x"40230f",x"2c180b",x"26160a",x"2e1a0c",x"2f1a0b",x"2c190b",x"341d0d",x"29170a",x"251509",x"1c1108",x"150e07",x"150e07",x"201309",x"3f2310",x"150e07",x"150e07",x"25150a",x"412511",x"180f07",x"29170a",x"361f0e",x"321d0d",x"311b0c",x"2d190b",x"2c190b",x"2a170a",x"1f1208",x"150e07",x"150e07",x"3a210f",x"2c1a0b",x"150e07",x"3a200e",x"2b180a",x"1e1208",x"2c190b",x"150e07",x"26160a",x"211309",x"150e07",x"150e07",x"150e07",x"150e07",x"29190d",x"29190d",x"28170b",x"20150c",x"20140c",x"20140b",x"24170d",x"23160d",x"26170d",x"28170c",x"29180c",x"301d0e",x"331d0e",x"371f0f",x"392010",x"392010",x"371f0f",x"361f0f",x"341d0e",x"331d0e",x"351d0e",x"341d0e",x"371f0f",x"381f0f",x"371e0f",x"3a2010",x"361e0e",x"361e0e",x"3b2110",x"381f0e",x"381f0e",x"381d0c",x"341b0b",x"331a0b",x"321a0b",x"2e190a",x"2a1709",x"261409",x"261509",x"251409",x"271509",x"29170a",x"28170a",x"27170b",x"23150b",x"201309",x"201209",x"20120a",x"21140c",x"28190e",x"2a1a0f",x"2b1b10",x"2a1b10",x"291a0f",x"2b1c12",x"2c1c12",x"2a1c11",x"2b1c12",x"2a1c12",x"27190f",x"27190f",x"2a1a0f",x"2b1b10",x"2d1d10",x"301d0f",x"2f1c0f",x"2c1b0e",x"2b1a0f",x"28180c",x"23160b",x"1f130a",x"1c120a",x"191109",x"2f1c0c",x"341e0e",x"331d0d",x"311b0c",x"351d0d",x"38200f",x"3c2310",x"39200e",x"371f0d",x"371e0d",x"3b210e",x"3c220f",x"3f2411",x"3d2310",x"3b2210",x"361f0e",x"321c0d",x"2f1b0c",x"2f1b0c",x"321d0d",x"351e0e",x"361f0e",x"351f0e",x"351e0e",x"331d0d",x"301b0c",x"2f1a0b",x"2b180a",x"28170a",x"2b180b",x"2d1a0b",x"2a170a",x"2b180a",x"311b0b",x"2e1a0b",x"2f1a0b",x"2d190a",x"2c180a",x"28170a",x"27160a",x"231309",x"27160a",x"29170a",x"29170a",x"261509",x"231409",x"201309",x"1e1208",x"1e1208",x"1f1208",x"211409",x"241509",x"27160a",x"2a180a",x"2e190b",x"321c0c",x"311b0c",x"301a0b",x"2f1a0b",x"2c180a",x"2d190b",x"2d190b",x"2b170a",x"2a160a",x"281509",x"271509",x"271609",x"271609",x"261509",x"251509",x"231409",x"1e1108",x"1a1008",x"452914",x"452914",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"211a14",x"211a14",x"211a14",x"201a13",x"1f1812",x"1f1811",x"1d160f",x"1b150e",x"19130c",x"17110a",x"150e07",x"150e07",x"543114",x"5b3616",x"5b3818",x"543315",x"503115",x"5e3b17",x"543416",x"472b13",x"432812",x"482c13",x"492c15",x"3e2512",x"3f2612",x"382111",x"3d2312",x"3e2513",x"3f2513",x"3c2311",x"3a2112",x"382011",x"351f10",x"362010",x"392112",x"3b2312",x"3c2413",x"3a2212",x"372011",x"331e10",x"301d0f",x"352010",x"351f10",x"362011",x"382111",x"3b2312",x"3a2212",x"3a2312",x"321e0f",x"3a2111",x"362010",x"3a2111",x"311d0f",x"3a2111",x"3b2111",x"3f2412",x"351f0f",x"392110",x"341f0f",x"3a2111",x"362011",x"382010",x"382111",x"382110",x"3c2211",x"3a2112",x"382011",x"382011",x"341f10",x"341f10",x"3d2412",x"382110",x"382111",x"351e0e",x"341d0e",x"371e0f",x"371f0f",x"3c2211",x"432713",x"432713",x"3e2311",x"3b2110",x"3b2110",x"3f2311",x"3d2311",x"3d2210",x"422411",x"3f2411",x"412411",x"402411",x"462713",x"502f16",x"502e16",x"5f4f43",x"554b41",x"52483e",x"150e07",x"160e07",x"160e07",x"231509",x"201308",x"231509",x"1f1308",x"1d1108",x"1d1208",x"201309",x"221409",x"241509",x"25150a",x"241509",x"241509",x"241509",x"25160a",x"241509",x"221409",x"1f1208",x"1e1108",x"1e1108",x"1f1208",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1c1108",x"1a1008",x"180f07",x"180f07",x"191008",x"1a1008",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"201309",x"221409",x"231509",x"231509",x"24150a",x"25160a",x"25160a",x"24150a",x"25160a",x"24150a",x"221409",x"211309",x"201309",x"1f1208",x"201208",x"1f1208",x"1d1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"1e1208",x"1a1008",x"1b1008",x"1a1008",x"191008",x"180f07",x"170f07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"3f2410",x"3f2410",x"3b210f",x"2b180b",x"341e0d",x"432611",x"25150a",x"2d1a0b",x"27160a",x"29170a",x"2a180b",x"27160a",x"29170a",x"2a180b",x"27170a",x"2b190b",x"1f1309",x"150e07",x"150e07",x"361f0e",x"2c1a0b",x"28170a",x"27160a",x"221409",x"27160a",x"231409",x"1b1108",x"150e07",x"150e07",x"442511",x"39200e",x"2a180b",x"150e07",x"29180b",x"38200e",x"211409",x"2c1a0b",x"2b190b",x"2c190b",x"29170a",x"241509",x"150e07",x"231509",x"341e0e",x"341d0d",x"351e0d",x"150e07",x"150e07",x"472912",x"27170a",x"1b1108",x"26160a",x"29170a",x"27160a",x"2c180b",x"28160a",x"28170a",x"27160a",x"231409",x"150e07",x"150e07",x"4f2d15",x"150e07",x"2e1a0b",x"3a200e",x"2e1a0b",x"3a200e",x"311b0b",x"241409",x"150e07",x"29170a",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"29190d",x"28170b",x"20150c",x"20140c",x"20140b",x"24170d",x"23160d",x"26170d",x"28170c",x"29180c",x"301d0e",x"331d0e",x"371f0f",x"392010",x"392010",x"371f0f",x"361f0f",x"341d0e",x"331d0e",x"351d0e",x"341d0e",x"371f0f",x"381f0f",x"371e0f",x"3a2010",x"361e0e",x"361e0e",x"3b2110",x"381f0e",x"381f0e",x"381d0c",x"341b0b",x"331a0b",x"321a0b",x"2e190a",x"2a1709",x"261409",x"261509",x"251409",x"271509",x"29170a",x"28170a",x"27170b",x"23150b",x"201309",x"201209",x"20120a",x"21140c",x"28190e",x"2a1a0f",x"2b1b10",x"2a1b10",x"291a0f",x"2b1c12",x"2c1c12",x"2a1c11",x"2b1c12",x"2a1c12",x"27190f",x"27190f",x"2a1a0f",x"2b1b10",x"2d1d10",x"301d0f",x"2f1c0f",x"2c1b0e",x"2b1a0f",x"28180c",x"23160b",x"1f130a",x"1c120a",x"191109",x"2f1c0c",x"341e0e",x"331d0d",x"311b0c",x"351d0d",x"38200f",x"3c2310",x"39200e",x"371f0d",x"371e0d",x"3b210e",x"3c220f",x"3f2411",x"3d2310",x"3b2210",x"361f0e",x"321c0d",x"2f1b0c",x"2f1b0c",x"321d0d",x"351e0e",x"361f0e",x"351f0e",x"351e0e",x"331d0d",x"301b0c",x"2f1a0b",x"2b180a",x"28170a",x"2b180b",x"2d1a0b",x"2a170a",x"2b180a",x"311b0b",x"2e1a0b",x"2f1a0b",x"2d190a",x"2c180a",x"28170a",x"27160a",x"231309",x"27160a",x"29170a",x"29170a",x"261509",x"231409",x"201309",x"1e1208",x"1e1208",x"1f1208",x"211409",x"241509",x"27160a",x"2a180a",x"2e190b",x"321c0c",x"311b0c",x"301a0b",x"2f1a0b",x"2c180a",x"2d190b",x"2d190b",x"2b170a",x"2a160a",x"281509",x"271509",x"271609",x"271609",x"261509",x"251509",x"231409",x"1e1108",x"1a1008",x"452914",x"452914",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"1f1811",x"211a14",x"201a13",x"211a14",x"1f1912",x"1f1912",x"1d1710",x"1c150e",x"1a130c",x"171009",x"150e07",x"150e07",x"573216",x"543114",x"5c3717",x"5f3a18",x"593517",x"573515",x"533113",x"4d2e13",x"482a11",x"4d2d14",x"442812",x"422611",x"402410",x"3f2411",x"3c2110",x"351e0e",x"351e0e",x"371f0f",x"3f2410",x"3d2211",x"3e2211",x"392010",x"3e2412",x"3f2512",x"3c2110",x"3a2010",x"371f0f",x"371e0f",x"38200f",x"331c0e",x"321c0d",x"38200f",x"38200f",x"3d2211",x"3d2311",x"3b2110",x"38200f",x"39200f",x"3c2110",x"3a2010",x"3c2211",x"3a2110",x"3e2210",x"341d0d",x"321c0d",x"3a200f",x"331d0e",x"351e0f",x"351d0e",x"3d2311",x"3d2311",x"392110",x"3e2412",x"382010",x"3d2311",x"3b2211",x"402412",x"3d2210",x"3c2211",x"3b2211",x"3c2211",x"341e0f",x"3b2110",x"3d2311",x"331d0e",x"361e0e",x"3d2211",x"3b2110",x"3b2111",x"3d2311",x"3d2311",x"3d2311",x"3f2311",x"442712",x"452713",x"3f2410",x"3e2210",x"462813",x"4b2d15",x"533218",x"4f2c14",x"4d2d15",x"554b41",x"160e07",x"160e07",x"160e07",x"160e07",x"201309",x"211409",x"231509",x"241609",x"1d1108",x"1d1208",x"201309",x"221409",x"241509",x"25150a",x"241509",x"241509",x"241509",x"25160a",x"241509",x"221409",x"1f1208",x"1e1108",x"1e1108",x"1f1208",x"1f1208",x"422511",x"371f0d",x"361e0d",x"2f1a0b",x"341d0d",x"2f1a0c",x"38200f",x"351e0e",x"311b0b",x"2f1a0b",x"321c0c",x"311b0c",x"301c0d",x"351e0d",x"361e0d",x"351e0d",x"341d0d",x"361f0e",x"2f1a0b",x"2f1a0b",x"351d0d",x"321c0c",x"301b0c",x"341d0d",x"351d0d",x"341d0d",x"39200e",x"341d0d",x"371f0e",x"341d0d",x"2f1a0b",x"331c0c",x"361e0d",x"331c0c",x"351e0d",x"321b0c",x"341d0d",x"341d0c",x"1c1108",x"1a1008",x"1b1008",x"1a1008",x"191008",x"180f07",x"170f07",x"341d0c",x"311b0b",x"301b0c",x"321c0c",x"351e0d",x"351d0d",x"331d0c",x"351d0d",x"351e0d",x"2e190b",x"341d0d",x"371f0d",x"341d0d",x"371f0e",x"341d0d",x"331c0c",x"301a0b",x"311b0c",x"351e0d",x"351d0d",x"321c0c",x"2f1b0b",x"2e1a0b",x"2f1a0b",x"281609",x"2d180a",x"2e1a0b",x"2f1a0b",x"2f1a0b",x"301a0b",x"311c0c",x"361e0d",x"361e0d",x"341d0d",x"321c0c",x"2d190b",x"341d0d",x"321c0c",x"351e0d",x"371f0e",x"301b0c",x"311c0c",x"331c0d",x"301b0c",x"361e0d",x"361e0d",x"341e0d",x"331d0d",x"341d0d",x"2d190b",x"2c190b",x"311c0c",x"331d0d",x"321c0c",x"371f0e",x"351e0d",x"361e0e",x"38200e",x"361e0d",x"351d0d",x"341d0d",x"381f0e",x"38200e",x"39210f",x"38200e",x"331c0d",x"311b0c",x"311c0c",x"321c0c",x"361e0e",x"361e0d",x"38200e",x"3a210f",x"361f0e",x"38200e",x"351e0d",x"341d0d",x"371f0d",x"381f0e",x"371f0e",x"38200e",x"321c0d",x"371f0e",x"371f0e",x"3a210f",x"39200f",x"341e0d",x"351d0d",x"311b0b",x"2e1a0b",x"351d0d",x"371f0e",x"351d0d",x"361e0d",x"311b0c",x"311b0c",x"311c0c",x"341d0d",x"361e0d",x"321c0c",x"361e0d",x"341d0d",x"331c0c",x"341d0c",x"321c0c",x"361e0d",x"361e0d",x"361e0d",x"351e0d",x"351e0d",x"341c0d",x"321c0c",x"321c0c",x"442611",x"341d0c",x"341d0c"),
(x"432611",x"432611",x"422511",x"2e1a0b",x"341d0d",x"3c200d",x"221309",x"2a180a",x"28170a",x"261509",x"281609",x"281609",x"261509",x"27160a",x"241409",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"381f0e",x"150e07",x"1e1208",x"201208",x"1b1008",x"150e07",x"150e07",x"150e07",x"432611",x"2c180b",x"27170a",x"24150a",x"150e07",x"150e07",x"2e1a0b",x"3a200e",x"201208",x"1d1108",x"27160a",x"26160a",x"150e07",x"150e07",x"381f0e",x"2e1a0b",x"381f0d",x"150e07",x"25160a",x"331d0d",x"150e07",x"201309",x"26160a",x"2a180b",x"29180b",x"2c190b",x"2d1a0b",x"251509",x"180f07",x"150e07",x"150e07",x"170f07",x"422511",x"150e07",x"412510",x"371f0e",x"351f0d",x"311c0c",x"150e07",x"27160a",x"28170a",x"150e07",x"27160a",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"201a13",x"211a14",x"211a13",x"201a13",x"1f1811",x"1f1811",x"1d160f",x"1b140d",x"19130c",x"171009",x"150e07",x"150e07",x"4d2c12",x"533115",x"513014",x"543215",x"533112",x"533113",x"4f2d12",x"472911",x"472912",x"41250f",x"452711",x"39200e",x"412410",x"452711",x"492a13",x"482913",x"412511",x"3e220f",x"3c200d",x"3d210e",x"3c210e",x"3f230f",x"412410",x"422611",x"442611",x"422510",x"432612",x"422611",x"3c220f",x"3e240f",x"412511",x"3f2411",x"402510",x"3a200e",x"391f0d",x"391f0e",x"3f2310",x"3d220f",x"3f230f",x"3e220f",x"3f220f",x"3d210e",x"361e0d",x"3d220f",x"3b200e",x"3a200e",x"39200e",x"39200e",x"391e0d",x"3f2310",x"3a210e",x"3a200e",x"3d220e",x"3b200e",x"3a210e",x"3d220f",x"3d220f",x"3c210e",x"371f0d",x"3f230f",x"39200e",x"3a200e",x"3e220f",x"3e220f",x"3f2410",x"3e2310",x"3e230f",x"3d220f",x"381f0d",x"381e0d",x"391f0d",x"3f230f",x"3f230f",x"3f220f",x"40230f",x"3e220e",x"42240f",x"442510",x"442510",x"482811",x"4b2a14",x"442611",x"512d15",x"26150a",x"331c0d",x"150e07",x"150e07",x"201208",x"201208",x"201208",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"564336",x"422511",x"371f0d",x"361e0d",x"2f1a0b",x"341d0d",x"2f1a0c",x"38200f",x"351e0e",x"311b0b",x"2f1a0b",x"321c0c",x"311b0c",x"301c0d",x"351e0d",x"361e0d",x"351e0d",x"341d0d",x"361f0e",x"2f1a0b",x"2f1a0b",x"351d0d",x"321c0c",x"301b0c",x"341d0d",x"351d0d",x"341d0d",x"39200e",x"341d0d",x"371f0e",x"341d0d",x"2f1a0b",x"331c0c",x"361e0d",x"331c0c",x"351e0d",x"321b0c",x"341d0d",x"341d0c",x"371e0d",x"381f0d",x"321c0c",x"381f0e",x"351d0c",x"331c0c",x"331c0c",x"341d0c",x"311b0b",x"301b0c",x"321c0c",x"351e0d",x"351d0d",x"331d0c",x"351d0d",x"351e0d",x"2e190b",x"341d0d",x"371f0d",x"341d0d",x"371f0e",x"341d0d",x"331c0c",x"301a0b",x"311b0c",x"351e0d",x"351d0d",x"321c0c",x"2f1b0b",x"2e1a0b",x"2f1a0b",x"281609",x"2d180a",x"2e1a0b",x"2f1a0b",x"2f1a0b",x"301a0b",x"311c0c",x"361e0d",x"361e0d",x"341d0d",x"321c0c",x"2d190b",x"341d0d",x"321c0c",x"351e0d",x"371f0e",x"301b0c",x"311c0c",x"331c0d",x"301b0c",x"361e0d",x"361e0d",x"341e0d",x"331d0d",x"341d0d",x"2d190b",x"2c190b",x"311c0c",x"331d0d",x"321c0c",x"371f0e",x"351e0d",x"361e0e",x"38200e",x"361e0d",x"351d0d",x"341d0d",x"381f0e",x"38200e",x"39210f",x"38200e",x"331c0d",x"311b0c",x"311c0c",x"321c0c",x"361e0e",x"361e0d",x"38200e",x"3a210f",x"361f0e",x"38200e",x"351e0d",x"341d0d",x"371f0d",x"381f0e",x"371f0e",x"38200e",x"321c0d",x"371f0e",x"371f0e",x"3a210f",x"39200f",x"341e0d",x"351d0d",x"311b0b",x"2e1a0b",x"351d0d",x"371f0e",x"351d0d",x"361e0d",x"311b0c",x"311b0c",x"311c0c",x"341d0d",x"361e0d",x"321c0c",x"361e0d",x"341d0d",x"331c0c",x"341d0c",x"321c0c",x"361e0d",x"361e0d",x"361e0d",x"351e0d",x"351e0d",x"341c0d",x"321c0c",x"321c0c",x"442611",x"341d0c",x"341d0c"),
(x"402411",x"402411",x"311b0c",x"2d190b",x"38200e",x"371f0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"391f0c",x"1a1008",x"251509",x"311b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"422510",x"331d0d",x"211409",x"27160a",x"241509",x"231409",x"241509",x"1e1208",x"150e07",x"150e07",x"3c220f",x"241509",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"2e1b0c",x"311c0c",x"1f1209",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1209",x"3c2210",x"402511",x"150e07",x"361e0d",x"3a200e",x"351d0d",x"311b0c",x"2f1b0c",x"371f0d",x"3b210e",x"311b0b",x"381f0d",x"150e07",x"29170a",x"190f08",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"211a14",x"201a13",x"201912",x"211a14",x"1f1912",x"1f1912",x"1d160f",x"1b140d",x"19130c",x"17110a",x"150e07",x"4d2c13",x"472910",x"4a2b11",x"502e14",x"523214",x"533115",x"523114",x"4c2d12",x"492a12",x"4a2c11",x"42270f",x"442711",x"3f2310",x"422511",x"462812",x"3f230f",x"3d230f",x"3e220f",x"482912",x"492a14",x"492a14",x"482a13",x"442711",x"412410",x"3f230f",x"3e230f",x"422511",x"422510",x"3f230f",x"412410",x"371e0d",x"3b210e",x"3e230f",x"3e2410",x"3e2310",x"3f2411",x"412411",x"3e220f",x"3e2310",x"3d230f",x"391e0d",x"3a200d",x"3a200e",x"402310",x"3d210e",x"3b200d",x"3d210e",x"3b1f0d",x"40230f",x"422410",x"3f230f",x"40230f",x"462711",x"3e220f",x"412410",x"3c210e",x"422510",x"3c210f",x"402410",x"462812",x"402410",x"442712",x"432611",x"3d220f",x"391f0d",x"432611",x"3f2410",x"3e220f",x"3d220f",x"40240f",x"40240f",x"3f230f",x"3f230f",x"3f230f",x"40230f",x"40230e",x"432510",x"40230f",x"41230e",x"41230e",x"3f210e",x"41230e",x"4c2a13",x"4c2a13",x"2d190b",x"2d190b",x"150e07",x"150e07",x"231409",x"221409",x"231509",x"231509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"59483b",x"59483b",x"462712",x"2d1a0b",x"2b190b",x"1c1108",x"201309",x"1a1008",x"150e07",x"1d1208",x"150e07",x"150e07",x"180f07",x"1d1208",x"1d1208",x"150e07",x"1d1208",x"191008",x"1d1108",x"170f07",x"1a1008",x"150e07",x"150e07",x"150e07",x"170f07",x"1b1108",x"150e07",x"170f07",x"180f07",x"1d1108",x"1e1209",x"150e07",x"1c1108",x"201309",x"1c1108",x"170f07",x"150e07",x"150e07",x"1a1008",x"180f07",x"150e07",x"170f07",x"191007",x"1d1108",x"1a1008",x"1a1008",x"180f07",x"150e07",x"150e07",x"201309",x"1a1008",x"1d1108",x"1d1108",x"190f08",x"150e07",x"1c1108",x"1d1208",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"1f1309",x"1d1108",x"1c1108",x"150e07",x"1a1008",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"190f07",x"1a1008",x"180f07",x"180f07",x"1f1208",x"231409",x"1c1108",x"150e07",x"1a1008",x"180f07",x"1d1108",x"170f07",x"1a1008",x"170f07",x"150e07",x"191008",x"1a1008",x"1c1108",x"1f1208",x"180f07",x"150e07",x"180f07",x"1a1008",x"1c1108",x"170f07",x"150e07",x"150e07",x"1e1208",x"191008",x"180f07",x"190f08",x"201309",x"1f1208",x"1c1108",x"201309",x"1e1208",x"1d1208",x"1d1208",x"211409",x"1b1108",x"180f08",x"1b1108",x"211309",x"1b1108",x"191008",x"1b1108",x"180f08",x"1c1108",x"1a1008",x"1a1008",x"211409",x"1f1208",x"1d1108",x"1c1108",x"221409",x"150e07",x"150e07",x"1d1208",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"1b1108",x"170f07",x"1c1108",x"1a1008",x"1f1208",x"150e07",x"1e1108",x"150e07",x"1a1008",x"1e1208",x"1c1108",x"170f07",x"170f07",x"170f07",x"180f08",x"150e07",x"1c1108",x"1a1008",x"170f07",x"170f07",x"150e07",x"150e07",x"2f1b0c",x"28170a",x"28170a"),
(x"3f230f",x"3f230f",x"3a200e",x"2a170a",x"331d0d",x"3b200e",x"492812",x"4d2b14",x"43240f",x"452510",x"492812",x"4a2913",x"462611",x"452611",x"43240f",x"42240e",x"42240f",x"371e0c",x"3c200d",x"3e220e",x"3b200d",x"381e0d",x"3d210d",x"3d210e",x"321b0b",x"271509",x"271509",x"3d210e",x"381f0d",x"321b0b",x"3d220f",x"402410",x"2e1a0b",x"3a210f",x"402511",x"3f2310",x"3a200e",x"3b210e",x"3b200e",x"4b2913",x"4a2a13",x"472812",x"452712",x"442711",x"3d2310",x"4f2d15",x"512e15",x"492812",x"422410",x"42240f",x"482812",x"4e2d14",x"543117",x"523017",x"543118",x"573319",x"4a2b14",x"492b14",x"4f2d15",x"3f230f",x"321c0b",x"2c180b",x"331c0c",x"3e220f",x"2a180b",x"432611",x"351d0d",x"2f1a0b",x"331c0c",x"351d0d",x"1a1008",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"484745",x"565555",x"494747",x"525251",x"4c4b4b",x"4d4d4d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494949",x"525252",x"000000",x"000000",x"000000",x"000000",x"353535",x"333333",x"333333",x"323232",x"323232",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"201a13",x"1f1912",x"201912",x"211a13",x"1f1811",x"1f1812",x"1d1610",x"1b150e",x"19120b",x"171009",x"150e07",x"523013",x"4e2d12",x"41260f",x"492c12",x"4b2c12",x"573514",x"4c2d12",x"4a2d12",x"4b2d12",x"422611",x"452910",x"41250f",x"371e0d",x"39200e",x"452812",x"472913",x"442813",x"472914",x"452813",x"492a14",x"4b2b15",x"482913",x"432510",x"41230f",x"40230f",x"40230f",x"3e220f",x"432611",x"432511",x"412510",x"3e220f",x"3b200e",x"3e220f",x"3f230f",x"3c210e",x"361e0c",x"371e0d",x"3e230f",x"3d220f",x"3b210e",x"3d210e",x"402410",x"3e220e",x"40240f",x"422410",x"422510",x"3f220f",x"422410",x"40230f",x"422410",x"41240f",x"442611",x"432510",x"472812",x"412410",x"402310",x"3f2310",x"3f2310",x"381f0e",x"40230f",x"412410",x"402410",x"3b200e",x"3b200e",x"3e230f",x"33190a",x"341b0b",x"361c0c",x"391f0d",x"3c210e",x"3b200e",x"3e220f",x"442611",x"3e220e",x"3b200e",x"422510",x"432511",x"40230f",x"3f230f",x"3b200d",x"3c200d",x"40220f",x"522e15",x"4c2a13",x"2d190b",x"2d190b",x"150e07",x"150e07",x"221409",x"221409",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5b4738",x"5b4738",x"492a13",x"321d0d",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"5d4d36",x"907659",x"967b5d",x"967d5d",x"8f7558",x"8c7459",x"967c5e",x"967c5d",x"957b5c",x"91795c",x"987b5f",x"93795d",x"957a5e",x"8c6f57",x"997e60",x"f8cea0",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331c0c",x"2b180b",x"2b180b"),
(x"3f2310",x"3f2310",x"3c210f",x"301b0c",x"351e0d",x"3f2310",x"241509",x"2d190b",x"2d1a0b",x"2e1a0b",x"301b0c",x"2a180a",x"2e1a0b",x"2d1a0b",x"2d190b",x"2c190b",x"2c190b",x"231509",x"251509",x"251509",x"1d1108",x"211409",x"150e07",x"150e07",x"3e220f",x"150e07",x"40230f",x"211309",x"150e07",x"150e07",x"150e07",x"150e07",x"482812",x"2f1a0b",x"1d1108",x"150e07",x"150e07",x"241409",x"311b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331c0b",x"150e07",x"211107",x"1b0f07",x"150e07",x"150e07",x"150e07",x"150e07",x"3d210d",x"1d1108",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e4c4a",x"454443",x"4a4847",x"484745",x"565555",x"5a5a5a",x"525251",x"4c4b4b",x"4d4d4d",x"404040",x"3f3f3f",x"444444",x"404040",x"383838",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5f5f5e",x"616161",x"494949",x"565656",x"4c4c4c",x"000000",x"000000",x"3c3c3c",x"3c3c3c",x"353535",x"333333",x"2f2f2f",x"2f2f2f",x"323232",x"323232",x"353535",x"434343",x"404040",x"322f2c",x"333333",x"3b3837",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201912",x"201912",x"211a14",x"211a14",x"201a13",x"201a13",x"201912",x"1f1811",x"1c160f",x"1c150f",x"19130c",x"17100a",x"150e07",x"513013",x"513013",x"3a230c",x"3b240c",x"39230c",x"36210b",x"331e0b",x"38220c",x"37210c",x"2a190a",x"2f1d0a",x"1f1208",x"1a1008",x"211308",x"221308",x"231409",x"211308",x"261509",x"231309",x"231309",x"241409",x"29170a",x"271509",x"221208",x"1e1007",x"1c1007",x"231308",x"251509",x"261509",x"271509",x"261509",x"251409",x"261509",x"261609",x"241509",x"29170a",x"29170a",x"2a180a",x"29170a",x"271509",x"271509",x"271509",x"29160a",x"27160a",x"28170a",x"2c190b",x"2b180b",x"29170a",x"2b180b",x"2b180b",x"29170a",x"2c180b",x"2a180a",x"2d190b",x"2b180b",x"2d190b",x"25160a",x"241509",x"251509",x"2a180b",x"2b190b",x"2f1b0c",x"321d0d",x"2e1b0c",x"2f1c0d",x"2c190b",x"301b0c",x"2e1a0b",x"311c0c",x"341e0d",x"321d0d",x"301b0c",x"2b180a",x"2d1a0b",x"2d1a0c",x"2c190b",x"2a180a",x"2d190b",x"2e1a0b",x"2c190b",x"29170a",x"311b0c",x"422511",x"472812",x"472812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c4536",x"5c4536",x"422410",x"29170a",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"574633",x"997e5f",x"947a5d",x"997e60",x"997e60",x"947a5c",x"806950",x"8a7156",x"846e52",x"806950",x"997e60",x"997e60",x"9a7e60",x"93785b",x"92775d",x"95785b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2b190b",x"2a180b",x"2a180b"),
(x"412511",x"412511",x"422511",x"331d0d",x"331c0c",x"3c210f",x"26160a",x"341d0d",x"321c0c",x"351e0d",x"351e0d",x"2e1a0b",x"2d190b",x"2c190b",x"2d190b",x"2e1a0b",x"2e1a0b",x"2a180a",x"2c190b",x"2c190b",x"2d190b",x"27160a",x"1b1008",x"150e07",x"150e07",x"341d0c",x"2b180a",x"1e1208",x"2b180a",x"231409",x"231509",x"150e07",x"150e07",x"2a180b",x"3d220f",x"180f08",x"402410",x"1e1208",x"150e07",x"211409",x"2b190b",x"2d1a0b",x"27170a",x"1d1208",x"231409",x"261609",x"241509",x"241409",x"261509",x"211309",x"28170a",x"2b180b",x"27160a",x"2c190b",x"2e1a0b",x"2a180a",x"251509",x"211409",x"150e07",x"150e07",x"2c190b",x"301a0b",x"170f07",x"251509",x"27160a",x"211409",x"150e07",x"150e07",x"201309",x"150e07",x"251509",x"1d1208",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"585656",x"565554",x"555452",x"464443",x"5d5b5b",x"696868",x"656464",x"626262",x"5d5d5d",x"575656",x"4b4b4b",x"414141",x"3f3f3f",x"444444",x"404040",x"363636",x"383838",x"464646",x"3e3e3e",x"000000",x"000000",x"606060",x"606060",x"5f5f5e",x"505050",x"545454",x"454545",x"3b3b3b",x"000000",x"5d5c5c",x"454545",x"414141",x"545454",x"535353",x"464646",x"303030",x"353535",x"323232",x"434343",x"404040",x"322f2c",x"393939",x"363535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"211a14",x"211b14",x"211a14",x"201913",x"1f1912",x"1f1912",x"1d1610",x"1c150e",x"19130c",x"17110a",x"150e07",x"150e07",x"432810",x"2c1c09",x"2d1c09",x"3b250b",x"33200b",x"2e1d0a",x"2f1d0a",x"301e0b",x"29190a",x"2a1a0a",x"1f1208",x"201308",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1e1208",x"1f1208",x"201309",x"221409",x"231409",x"231409",x"241509",x"251509",x"26160a",x"27170a",x"28170a",x"29180b",x"29180b",x"28170a",x"26160a",x"251509",x"241509",x"24150a",x"231409",x"221409",x"211309",x"201309",x"1f1209",x"1d1208",x"1c1108",x"1b1108",x"1b1108",x"1b1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1308",x"201309",x"211409",x"221409",x"231409",x"25160a",x"26160a",x"27160a",x"27160a",x"26160a",x"27160a",x"241509",x"241509",x"221409",x"201309",x"1c1108",x"180f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301c0c",x"412410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e4635",x"5e4635",x"422511",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"63533e",x"715b44",x"7b664d",x"997e60",x"997e60",x"92775b",x"997e60",x"987d5e",x"977f61",x"997e60",x"997e60",x"997e60",x"997d5e",x"9c7f62",x"93795c",x"8d7358",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0b",x"301b0c",x"301b0c"),
(x"402410",x"402410",x"402410",x"331d0d",x"331c0c",x"432611",x"2d190b",x"301b0c",x"301b0c",x"331c0c",x"301b0c",x"341d0d",x"341d0d",x"2f1b0c",x"29170a",x"29170a",x"2b180b",x"321c0c",x"2d190b",x"2c190b",x"241509",x"2d190b",x"241509",x"150e07",x"150e07",x"150e07",x"211308",x"251509",x"2c190b",x"2b180b",x"27160a",x"221409",x"150e07",x"150e07",x"191008",x"331b0b",x"170f07",x"1e1208",x"27160a",x"29170a",x"2a180a",x"2f1a0b",x"29170a",x"29180a",x"25160a",x"321c0d",x"28170a",x"2c190b",x"27160a",x"25160a",x"2d1a0b",x"2d1a0b",x"2e1a0b",x"2e1a0b",x"29170a",x"2c190b",x"29170a",x"27160a",x"1f1208",x"150e07",x"150e07",x"271609",x"221409",x"29170a",x"29170a",x"28160a",x"1d1108",x"150e07",x"150e07",x"371f0d",x"211409",x"211409",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5f5d5d",x"585656",x"646363",x"666565",x"343332",x"353433",x"353434",x"333333",x"393838",x"353433",x"555555",x"616161",x"555555",x"4a413e",x"404040",x"3d3d3d",x"3c3c3c",x"424242",x"373736",x"383838",x"3a3a3a",x"4c4c4c",x"585858",x"626262",x"545454",x"5d5d5d",x"343434",x"343434",x"5e5d5d",x"5e5d5d",x"5d5d5d",x"6a6a6a",x"585858",x"4b4b4b",x"4a4a4a",x"4f4f4f",x"494949",x"2e2e2e",x"383838",x"616161",x"505050",x"2b2b2b",x"2f2e2e",x"2f2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a14",x"201a14",x"201912",x"201a13",x"201a13",x"201a13",x"1f1811",x"1f1811",x"1c160f",x"1b140d",x"19120b",x"150e07",x"150e07",x"150e07",x"2f1d0a",x"301e0a",x"33200a",x"301f0a",x"3a240b",x"2c1b0a",x"291a0a",x"2c1b0a",x"271809",x"261709",x"231509",x"291a09",x"1f1308",x"1e1208",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1e1108",x"1f1208",x"201208",x"211409",x"231409",x"231409",x"231409",x"241509",x"251509",x"27160a",x"28160a",x"27160a",x"26160a",x"26160a",x"27160a",x"27160a",x"26160a",x"241509",x"25160a",x"25160a",x"25160a",x"25160a",x"24150a",x"211409",x"1f1309",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1e1208",x"201309",x"201409",x"201309",x"211409",x"23150a",x"24150a",x"241509",x"26160a",x"26160a",x"27170a",x"29180b",x"2b190b",x"2b190b",x"2a180b",x"28170a",x"26160a",x"231409",x"201309",x"1c1108",x"191008",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583e2d",x"583e2d",x"482912",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"705b46",x"997e60",x"9a7f60",x"997e60",x"997e60",x"997e60",x"997e60",x"997e60",x"997e60",x"94795c",x"987c5e",x"997e60",x"997e60",x"987c60",x"987d5e",x"6e5b43",x"180f07",x"170f07",x"160e07",x"150e07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"160f07",x"160f07",x"150e07",x"150e07",x"160e07",x"150e07",x"160f07",x"160f07",x"150e07",x"160f07",x"160e07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"160f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1a0b",x"341e0e",x"341e0e"),
(x"3d220f",x"3d220f",x"3f2410",x"331d0d",x"341c0c",x"361d0c",x"1e1108",x"271509",x"261409",x"291609",x"2d190b",x"2f1a0b",x"2c190a",x"2f1a0b",x"29170a",x"29170a",x"281509",x"271509",x"2b180a",x"29170a",x"28160a",x"221409",x"211409",x"170f07",x"150e07",x"432611",x"28170a",x"251609",x"29170a",x"241509",x"28160a",x"1b1108",x"150e07",x"150e07",x"371d0c",x"160f07",x"1d1108",x"261409",x"261509",x"2c190b",x"29170a",x"28160a",x"281609",x"241409",x"221409",x"2b180a",x"231409",x"29170a",x"261609",x"2b180b",x"2a170a",x"27160a",x"2b180b",x"311b0c",x"2c190b",x"2d1a0c",x"2b190b",x"27170a",x"201309",x"150e07",x"482912",x"331c0c",x"251509",x"29170a",x"251509",x"241509",x"1d1108",x"150e07",x"150e07",x"3d230f",x"231509",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"606060",x"606060",x"646464",x"595858",x"333232",x"363432",x"343332",x"4d4d4d",x"434343",x"3a3a3a",x"333333",x"424242",x"3c3c3c",x"3b3b3b",x"5d5d5d",x"4a4a4a",x"3f3f3f",x"3b3b3b",x"343434",x"353535",x"404040",x"383838",x"373737",x"474747",x"515151",x"555555",x"5a5a5a",x"313131",x"313131",x"000000",x"5a5959",x"545454",x"3e3e3e",x"303030",x"362e28",x"2e2e2e",x"4b4b4b",x"464747",x"343434",x"3a3a3a",x"4f4f4f",x"3d3d3d",x"303030",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b3b3a",x"3d3d3d",x"3e3e3e",x"3e3e3e",x"404040",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a14",x"201a14",x"1f1811",x"211a14",x"211a14",x"201912",x"1f1811",x"1d160f",x"1d1710",x"1c150e",x"19120b",x"150e07",x"150e07",x"150e07",x"34210b",x"33200b",x"311f0a",x"2e1d0a",x"33200a",x"311f0a",x"251708",x"1f1309",x"281909",x"271809",x"241609",x"211408",x"1c1108",x"1d1108",x"1e1208",x"1f1209",x"1f1309",x"201309",x"1f1309",x"201309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"221409",x"211409",x"211309",x"231409",x"241509",x"25150a",x"27170a",x"29180b",x"28170a",x"2b190b",x"2c1a0c",x"2d1a0c",x"2c1a0c",x"2d1a0c",x"2c190b",x"2b190b",x"2b190c",x"2b190b",x"2a180b",x"27160a",x"25150a",x"25150a",x"241509",x"221409",x"221409",x"201309",x"1e1208",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1f1309",x"201309",x"1f1208",x"211409",x"211409",x"221409",x"25150a",x"241509",x"27160a",x"28170a",x"261509",x"241409",x"241409",x"241409",x"231309",x"201208",x"1f1108",x"1c1108",x"1a1008",x"180f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563f31",x"563f31",x"351c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"554333",x"8a7158",x"907559",x"735d47",x"856c53",x"836d52",x"846c52",x"8c7558",x"988062",x"917a5c",x"8b7357",x"897055",x"7e684f",x"836c51",x"8d7359",x"4f3f2e",x"1d1308",x"1b1108",x"181007",x"180f07",x"1c1208",x"1c1208",x"191007",x"1b1108",x"1a1107",x"160f07",x"181007",x"170f07",x"160f07",x"170f07",x"150e07",x"181007",x"181007",x"160f07",x"191007",x"170f07",x"191007",x"170f07",x"170f07",x"170f07",x"150e07",x"191007",x"191107",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"361f0e",x"361f0e"),
(x"391f0e",x"391f0e",x"3e2310",x"331d0d",x"321c0c",x"432511",x"241509",x"28170a",x"2c190b",x"2a180b",x"301c0c",x"2e1a0c",x"301b0c",x"2e190b",x"311c0c",x"2f1b0b",x"2d190b",x"2c190b",x"2d190b",x"2d190b",x"28170a",x"241509",x"150e07",x"150e07",x"150e07",x"150e07",x"2d190b",x"150e07",x"251509",x"231409",x"201308",x"150e07",x"150e07",x"4a2912",x"1c1108",x"1f1208",x"261609",x"2a170a",x"2d190b",x"29180a",x"27160a",x"26160a",x"221409",x"241509",x"241509",x"251509",x"28160a",x"28170a",x"29170b",x"27170a",x"27170a",x"2d1a0b",x"2b190b",x"2d1a0c",x"2e1b0c",x"2c190b",x"211309",x"23150a",x"150e07",x"150e07",x"341d0d",x"432611",x"150e07",x"241409",x"26160a",x"1d1208",x"150e07",x"150e07",x"432510",x"1f1208",x"201309",x"1a1108",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"676665",x"676665",x"5d5d5d",x"323232",x"333232",x"333232",x"565454",x"565454",x"4b4a4a",x"474747",x"333333",x"323232",x"333333",x"353535",x"3f3f3f",x"4c4c4c",x"4c4c4c",x"414141",x"3f3f3f",x"343434",x"383838",x"373737",x"353535",x"474747",x"454545",x"444444",x"353535",x"313131",x"323232",x"000000",x"545454",x"474646",x"383838",x"323232",x"323231",x"343332",x"3f3f3f",x"4f4f4f",x"525252",x"575757",x"474747",x"303030",x"313131",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"323232",x"343434",x"3d3d3d",x"3b3b3b",x"3b3b3a",x"3d3d3d",x"3e3e3e",x"3e3e3e",x"404040",x"353535",x"343434",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1912",x"1f1912",x"211a13",x"1f1912",x"201a13",x"1f1811",x"1f1912",x"1d1710",x"1d1711",x"1b140e",x"19120c",x"150e07",x"150e07",x"150e07",x"000000",x"301f0a",x"2d1d09",x"2b1b09",x"301e0a",x"34210b",x"2b1b0a",x"211409",x"261709",x"1d1208",x"201409",x"1f1309",x"1f1309",x"1f1309",x"201309",x"201309",x"201309",x"201309",x"201309",x"211409",x"201309",x"201309",x"201309",x"211409",x"211309",x"221409",x"25160a",x"25160a",x"25150a",x"221409",x"241509",x"261509",x"26160a",x"27160a",x"29170a",x"2a180b",x"2d1a0c",x"2e1b0c",x"2d1a0c",x"2c1a0b",x"2c190b",x"2a190b",x"2a180b",x"28170a",x"2a180b",x"28170a",x"27160a",x"27170a",x"25160a",x"24150a",x"221409",x"211409",x"201309",x"1f1309",x"201309",x"211409",x"211409",x"221409",x"211309",x"211409",x"211309",x"24160a",x"25160a",x"26160a",x"27160a",x"28170a",x"29170a",x"2a170a",x"2b180b",x"2b190b",x"2a180a",x"26160a",x"241509",x"221409",x"1d1208",x"190f08",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"49392e",x"49392e",x"40230f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"170f07",x"191007",x"1c1208",x"1a1107",x"1b1108",x"191007",x"1f1408",x"1b1108",x"1b1108",x"1b1108",x"201508",x"211508",x"1f1408",x"191007",x"180f07",x"1e1308",x"1d1208",x"1b1108",x"1d1308",x"1d1208",x"170f07",x"191007",x"180f07",x"170f07",x"191007",x"160e07",x"1a1107",x"1a1107",x"170f07",x"1b1108",x"181007",x"1b1108",x"181007",x"191007",x"191007",x"150e07",x"1b1108",x"1c1208",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"38200e",x"38200e"),
(x"3c210e",x"3c210e",x"432511",x"311c0c",x"301a0b",x"3a200e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3b200e",x"170f07",x"371e0d",x"321c0c",x"150e07",x"150e07",x"150e07",x"1a1008",x"422510",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"30190a",x"1e1208",x"150e07",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"29170a",x"170f07",x"150e07",x"201309",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"656463",x"656463",x"5f5f5f",x"323232",x"323232",x"000000",x"5f5d5d",x"5f5d5d",x"5d5d5d",x"505050",x"404040",x"3b3b3b",x"323232",x"3f3e3e",x"4b4b4b",x"5b5b5b",x"515151",x"4a4a4a",x"464646",x"434343",x"484848",x"474747",x"525252",x"434343",x"4e4e4e",x"323232",x"323232",x"353535",x"000000",x"000000",x"000000",x"383838",x"383838",x"323232",x"323232",x"474747",x"4a4a4a",x"4a4a4a",x"292929",x"2f2f2f",x"454545",x"3f3f3f",x"2f2f2f",x"323232",x"333333",x"343434",x"353535",x"333333",x"333333",x"323232",x"343434",x"3d3d3d",x"3e3e3e",x"3e3e3e",x"4f4f4f",x"4d4d4d",x"474747",x"4a4a4a",x"3a3a3a",x"373737",x"3a3a3a",x"454545",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"211a14",x"201912",x"201a13",x"1f1811",x"1f1812",x"1d1710",x"1d160f",x"1b140d",x"17110a",x"150e07",x"150e07",x"150e07",x"000000",x"2d1d0a",x"2b1b0a",x"1f1308",x"241708",x"281909",x"231609",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1f1208",x"1f1309",x"201309",x"201309",x"201309",x"201309",x"201309",x"1c1108",x"221409",x"201309",x"201208",x"241509",x"26160a",x"26160a",x"25150a",x"25150a",x"28170a",x"2b190c",x"2c1a0c",x"2a180b",x"2a180b",x"2c190b",x"2c190b",x"2d1a0c",x"2c1a0b",x"2a180b",x"2a180b",x"2a180b",x"28170a",x"28160a",x"2a190b",x"29180b",x"27160a",x"251509",x"211308",x"201208",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"1f1208",x"201309",x"211409",x"221409",x"221409",x"23150a",x"23150a",x"24150a",x"25150a",x"251509",x"29170a",x"2a180b",x"2b180b",x"2c190b",x"2c190b",x"2b180b",x"29180a",x"28170a",x"26160a",x"231509",x"1d1208",x"180f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463528",x"40230f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"170f07",x"1a1107",x"1d1208",x"1b1208",x"1c1208",x"191007",x"201508",x"1c1208",x"1d1208",x"1c1208",x"221508",x"221608",x"1f1408",x"1b1108",x"170f07",x"1e1308",x"1d1308",x"1c1208",x"1f1408",x"1e1308",x"170f07",x"1b1108",x"181007",x"180f07",x"191107",x"160e07",x"1b1108",x"1b1108",x"180f07",x"1b1108",x"191007",x"1b1108",x"181007",x"1a1107",x"191007",x"160e07",x"1c1208",x"1c1208",x"1a1107",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"150e07",x"150e07",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1f1309",x"150e07",x"1f1209",x"150e07",x"1e1208",x"150e07",x"1a1008",x"150e07",x"150e07",x"27170b",x"452813",x"452813"),
(x"311b0c",x"311b0c",x"3b210e",x"2e1a0b",x"341c0c",x"39200e",x"3c210e",x"422410",x"402310",x"422510",x"452712",x"462711",x"442611",x"462712",x"432510",x"40230f",x"3d220f",x"412511",x"472912",x"3f2310",x"462711",x"3f230f",x"371e0d",x"381f0d",x"3a210f",x"3c220f",x"3a210f",x"3e2310",x"3f2410",x"412410",x"3c210e",x"2f1a0b",x"321c0b",x"41230f",x"3c200d",x"391e0c",x"3c200d",x"40240f",x"452611",x"432510",x"3f220f",x"432510",x"3e220f",x"3c220f",x"40230f",x"3e220f",x"3c220f",x"422611",x"3e230f",x"3f2410",x"432611",x"3e220f",x"3b200e",x"412511",x"3e220f",x"3d220f",x"402410",x"3f2410",x"3a200f",x"2f1a0b",x"341c0c",x"361e0d",x"36200e",x"402410",x"402410",x"3a210f",x"2b180b",x"311b0c",x"39200f",x"301c0c",x"211409",x"1d1209",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5857",x"565655",x"5f5f5f",x"333333",x"393939",x"343433",x"4f4f4f",x"4f4f4f",x"595959",x"515151",x"4b4b4b",x"585858",x"565656",x"505050",x"323232",x"393939",x"565656",x"555555",x"535353",x"505050",x"4b4b4b",x"4f4f4f",x"434343",x"545454",x"494949",x"3b3b3b",x"383838",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"2b2b2b",x"242323",x"393939",x"5c5c5c",x"323232",x"353535",x"4d4d4d",x"585858",x"484848",x"313131",x"313131",x"353535",x"353535",x"3c3c3c",x"343434",x"343434",x"373737",x"4f4f4f",x"575757",x"4b4b4b",x"454545",x"393939",x"454545",x"424242",x"494949",x"4f4f4f",x"424242",x"4e4e4e",x"484848",x"484848",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a14",x"201a14",x"201912",x"1f1812",x"201a13",x"1e1811",x"1e1711",x"1d1610",x"1b140d",x"1a130c",x"171009",x"150e07",x"150e07",x"150e07",x"1e150a",x"1f150a",x"1a1107",x"171007",x"191007",x"1b1107",x"221509",x"1b1108",x"1c1108",x"1e1208",x"1d1208",x"1e1208",x"1f1209",x"1e1208",x"1e1208",x"1f1309",x"1f1208",x"1f1208",x"1f1309",x"1f1208",x"201309",x"1f1208",x"201309",x"221409",x"24150a",x"24150a",x"241509",x"27160a",x"241509",x"27160a",x"29180b",x"27170a",x"251509",x"251509",x"29180b",x"29180b",x"261509",x"241409",x"251509",x"29170a",x"27160a",x"261509",x"26160a",x"27160a",x"26160a",x"26160a",x"261509",x"26160a",x"251509",x"231409",x"221409",x"211409",x"201309",x"1f1208",x"1f1208",x"211309",x"201309",x"201309",x"201309",x"201309",x"211309",x"211309",x"231409",x"26160a",x"28170a",x"29180b",x"2a180b",x"2b180b",x"2b180b",x"2a180a",x"27160a",x"25150a",x"231409",x"1f1309",x"1b1108",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"342619",x"322518",x"2f2318",x"2f2317",x"32251a",x"302318",x"2f2318",x"2e2318",x"2f2318",x"302418",x"312419",x"2d2116",x"2f2217",x"332518",x"2f2316",x"2f2317",x"2f2216",x"302417",x"2c2115",x"291f15",x"2c2116",x"291f15",x"2a1f15",x"2a1e14",x"281d13",x"2a1f14",x"2d2014",x"463528",x"40230f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"170f07",x"1a1107",x"1d1208",x"1b1208",x"1c1208",x"191007",x"201508",x"1c1208",x"1d1208",x"1c1208",x"221508",x"221608",x"1f1408",x"1b1108",x"170f07",x"1e1308",x"1d1308",x"1c1208",x"1f1408",x"1e1308",x"170f07",x"1b1108",x"181007",x"180f07",x"191107",x"160e07",x"1b1108",x"1b1108",x"180f07",x"1b1108",x"191007",x"1b1108",x"181007",x"1a1107",x"191007",x"160e07",x"1c1208",x"1c1208",x"1a1107",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"150e07",x"150e07",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1e1208",x"150e07",x"1f1309",x"150e07",x"1f1209",x"150e07",x"1e1208",x"150e07",x"1a1008",x"150e07",x"150e07",x"27170b",x"452813",x"000000"),
(x"331b0b",x"331b0b",x"321a0b",x"291609",x"291609",x"271509",x"241208",x"2a1609",x"2a1609",x"2d180a",x"291509",x"2b1609",x"2e190b",x"321c0c",x"331c0c",x"351d0d",x"311b0c",x"2d190b",x"2d190b",x"301b0c",x"351d0d",x"331c0c",x"321c0c",x"2d180a",x"2d180a",x"371f0d",x"371e0d",x"301b0b",x"341d0d",x"331c0c",x"371f0d",x"2c170a",x"351e0d",x"331c0c",x"331c0c",x"351d0d",x"331c0c",x"321c0c",x"311b0b",x"321c0c",x"29170a",x"2c180a",x"311b0c",x"2e1a0b",x"301b0c",x"301b0c",x"321c0c",x"28160a",x"2e190b",x"221208",x"231308",x"271509",x"291609",x"2a170a",x"2a170a",x"2f1b0c",x"2c190b",x"2d1a0b",x"2e1a0b",x"2e1a0b",x"2e1a0b",x"2f1b0c",x"311c0c",x"311c0c",x"341d0d",x"301b0c",x"2a180a",x"2f1b0c",x"2d190b",x"2d190b",x"2b190c",x"27170b",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"515151",x"575757",x"5a5a5a",x"545454",x"343433",x"323232",x"373737",x"474442",x"505050",x"4f4f4f",x"4f4f4f",x"272727",x"303030",x"4a4a4a",x"333333",x"3d3d3d",x"565656",x"5e5e5e",x"404040",x"515151",x"4f4f4f",x"5e5e5e",x"333333",x"474747",x"5b5b5b",x"4d4d4d",x"343434",x"323232",x"363636",x"414141",x"555555",x"474747",x"494949",x"454545",x"303030",x"1f1f1f",x"616161",x"313131",x"313131",x"4d4d4d",x"535353",x"4d4d4d",x"565656",x"636363",x"5b5b5b",x"545454",x"4e4e4e",x"595959",x"5e5e5e",x"5e5754",x"555555",x"4c4c4c",x"464646",x"404040",x"3c3c3c",x"414141",x"424242",x"424242",x"474747",x"4b4b4b",x"535353",x"464646",x"3b3b3b",x"3b3b3b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a13",x"201a13",x"201a13",x"211a14",x"1f1811",x"1f1811",x"1d160f",x"1d1710",x"1b140d",x"19130c",x"17100a",x"150e07",x"150e07",x"150e07",x"1e150a",x"1f150a",x"1c130a",x"1f1408",x"170f07",x"170f07",x"190f08",x"1a1008",x"1b1008",x"1b1108",x"1a1008",x"190f07",x"1a0f07",x"1b1008",x"1b1008",x"1b1008",x"1c1108",x"1e1208",x"1e1208",x"1f1208",x"1d1108",x"1e1208",x"201309",x"211409",x"221409",x"24150a",x"221409",x"231409",x"241409",x"26160a",x"231409",x"27170a",x"28180b",x"28180b",x"29180b",x"2a190b",x"2a190b",x"2b190b",x"2b190b",x"2b190b",x"29170a",x"27160a",x"27160a",x"27160a",x"26150a",x"251509",x"241409",x"251509",x"251509",x"241409",x"211309",x"201309",x"201309",x"1f1208",x"1f1208",x"201208",x"201308",x"201309",x"201309",x"201309",x"201309",x"211309",x"221409",x"241509",x"231309",x"241409",x"241409",x"241409",x"231408",x"221208",x"1f1108",x"1d1108",x"1d1108",x"1b1008",x"180f07",x"160e07",x"150e07",x"150e07",x"2f2216",x"332518",x"342619",x"322518",x"2f2318",x"2f2317",x"32251a",x"302318",x"2f2318",x"2e2318",x"2f2318",x"302418",x"312419",x"2d2116",x"2f2217",x"332518",x"2f2316",x"2f2317",x"2f2216",x"302417",x"2c2115",x"291f15",x"2c2116",x"291f15",x"2a1f15",x"2a1e14",x"281d13",x"2a1f14",x"2d2014",x"241b13",x"271d13",x"211911",x"241b12",x"241b12",x"251c12",x"261c10",x"2d1f11",x"2e2011",x"312111",x"322211",x"2f2011",x"302111",x"2b1d11",x"2a1c0f",x"2b1d0f",x"2a1c0f",x"2d1e0f",x"2d1e0f",x"2b1d10",x"2a1d0f",x"291c0e",x"26190c",x"26190c",x"22180d",x"1f160d",x"1b140c",x"1d150c",x"1c140c",x"291b0b",x"17110a",x"18110a",x"1b1209",x"1a1107",x"1b1108",x"160f07",x"170f07",x"1f150b",x"1a1109",x"1a110a",x"1c130a",x"23170b",x"1b120a",x"1d140b",x"1b130a",x"22170d",x"23190f",x"1f160c",x"19120c",x"17110a",x"17110a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"381f0e",x"381f0e",x"381f0e",x"2c190b",x"2f1b0c",x"321c0c",x"351e0d",x"321c0c",x"371f0e",x"361f0e",x"361f0e",x"38210f",x"38200f",x"2e190b",x"2d180a",x"2f1a0c",x"361f0e",x"301c0d",x"2e1a0c",x"311c0c",x"301b0c",x"331d0d",x"341d0d",x"311b0c",x"301a0b",x"2a170a",x"331c0c",x"361f0d",x"301a0b",x"301b0b",x"2f1a0b",x"2f1a0b",x"331c0d",x"331d0d",x"311c0c",x"2e1a0b",x"2f1b0b",x"2b180b",x"2e1a0b",x"2d190b",x"2b180a",x"2a170a",x"281609",x"261509",x"291609",x"29170a",x"2a180a",x"301b0c",x"29180b",x"27170a",x"2b180b",x"2e1a0c",x"251509",x"29170a",x"261509",x"2b180a",x"221309",x"221309",x"271509",x"271509",x"281509",x"261509",x"2b180a",x"29170a",x"2c180b",x"28170a",x"2a170a",x"2c190b",x"2d1a0b",x"2a180b",x"27170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"515151",x"545454",x"676767",x"4e4e4e",x"323232",x"363636",x"464646",x"5c5c5c",x"454545",x"1a1a1a",x"2d2d2d",x"313131",x"4a4a4a",x"333333",x"565656",x"626262",x"5b5b5b",x"3c3c3c",x"4d4d4d",x"646464",x"3a3a3a",x"373737",x"5c5c5c",x"4c4c4c",x"555555",x"5f5f5f",x"2e2e2e",x"3e3e3e",x"414141",x"555555",x"515151",x"494949",x"4f4f4f",x"5e5e5e",x"4b4b4b",x"292929",x"2d2d2d",x"363535",x"000000",x"4d4d4d",x"484848",x"414141",x"363636",x"393939",x"4c4c4c",x"606060",x"5c5c5c",x"545454",x"464646",x"444444",x"4a4a4a",x"484848",x"383838",x"3a3a3a",x"3f3f3f",x"575757",x"4b4b4b",x"4b4b4b",x"434343",x"313131",x"323232",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"201a14",x"201a14",x"201a13",x"1e1710",x"1f1811",x"1f1812",x"1d160f",x"1d1610",x"1b150e",x"1a130c",x"17110a",x"150e07",x"150e07",x"1c130a",x"1d140a",x"1e150a",x"1b120a",x"1f1408",x"241708",x"201408",x"1f150b",x"21160a",x"20160b",x"24180b",x"21160b",x"271a0c",x"281a0e",x"22180d",x"2c1d10",x"2b1e0f",x"251a0e",x"2c1e11",x"271c11",x"2a1d10",x"332311",x"3a2712",x"2a1d11",x"2d1f11",x"2c1e11",x"2a1c0f",x"2d1f11",x"261b10",x"2b1d0f",x"2f1f10",x"332210",x"34220f",x"342312",x"332312",x"372512",x"2f1f11",x"302011",x"332212",x"302112",x"2e2013",x"312213",x"322214",x"322316",x"352515",x"342415",x"362617",x"382717",x"382819",x"3a2716",x"372716",x"392818",x"382818",x"372618",x"372718",x"3a2818",x"372618",x"342518",x"342517",x"392718",x"362618",x"372719",x"362619",x"322316",x"322419",x"35261a",x"322418",x"35271a",x"362619",x"39281a",x"362619",x"342619",x"352619",x"372719",x"362719",x"332416",x"302316",x"332519",x"342617",x"2d2216",x"332519",x"322619",x"312519",x"2e2317",x"302418",x"33261a",x"2f2317",x"2e2318",x"2d2318",x"2f2318",x"312519",x"31251a",x"2b2014",x"2f2216",x"322518",x"312316",x"2e2317",x"2e2116",x"322518",x"2c2115",x"2a2016",x"2e2216",x"291e14",x"2b1f15",x"2b1f14",x"2a1e14",x"2a1f14",x"281d13",x"231b12",x"251c13",x"211a12",x"241b13",x"251c13",x"261c12",x"251b10",x"2e1f11",x"2e2011",x"2e2011",x"352412",x"2f2011",x"312212",x"2a1d11",x"261a0e",x"2d1f0f",x"261a0e",x"2f200f",x"2b1d0f",x"2d1e10",x"271b0f",x"2a1c0e",x"25190c",x"26190d",x"22180d",x"20160d",x"1a140c",x"1f160d",x"1b130b",x"3a250d",x"17100a",x"18110a",x"1b1309",x"191007",x"1b1108",x"160f07",x"170f07",x"21170b",x"1a1109",x"181009",x"18110a",x"23170a",x"1d130a",x"23170b",x"1c1309",x"1c140c",x"23190f",x"1f160c",x"19120c",x"171009",x"17110a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"2a180a",x"351d0d",x"39200e",x"39200f",x"2f1b0c",x"2f1b0c",x"241509",x"231509",x"2a190b",x"2f1c0c",x"301c0c",x"2f1b0c",x"180f08",x"211409",x"341d0d",x"2f1b0c",x"301b0c",x"2c190b",x"2f1b0c",x"2e1a0b",x"2d190b",x"2c190b",x"2a180a",x"2c190b",x"2b180a",x"2b180a",x"2d190b",x"2c180b",x"26160a",x"2a180a",x"2d1a0b",x"2f1b0c",x"2d1a0b",x"29170a",x"2f1b0c",x"2d1a0b",x"341d0d",x"311b0c",x"2d190b",x"2c190b",x"2e1a0b",x"301b0b",x"331c0c",x"2f1b0c",x"311c0c",x"29160a",x"301a0b",x"311b0b",x"321c0c",x"2d180a",x"2b170a",x"2a170a",x"2d190b",x"29170a",x"221409",x"2b180a",x"301a0b",x"2e190b",x"301b0c",x"341d0d",x"351e0d",x"301b0b",x"2d190b",x"301b0c",x"321c0c",x"29170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"5a5a5a",x"535353",x"575757",x"626262",x"616161",x"5e5e5e",x"5b5b5b",x"515151",x"303030",x"212121",x"2c2c2c",x"000000",x"000000",x"000000",x"5d5c5c",x"5b5b5b",x"5b5b5b",x"4d4d4d",x"3e3e3e",x"3a3a3a",x"313232",x"5e5e5e",x"474747",x"444444",x"3f3f3f",x"565656",x"646464",x"646464",x"686868",x"5f5f5f",x"5e5e5e",x"525252",x"202020",x"2f2f2f",x"2f2f2f",x"202020",x"000000",x"000000",x"000000",x"000000",x"373737",x"363636",x"353535",x"343434",x"393939",x"3f3f3f",x"3a3a3a",x"3f3f3f",x"444444",x"444444",x"525252",x"424242",x"303030",x"323232",x"3b3b3b",x"313131",x"313131",x"333333",x"313131",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1811",x"1f1811",x"201912",x"211a14",x"1f1811",x"1f1811",x"1e1711",x"1d1710",x"1b140e",x"19130c",x"17110a",x"150e07",x"150e07",x"1a1108",x"1c1208",x"1f1408",x"1b1108",x"231608",x"201408",x"1f1408",x"221508",x"231608",x"201408",x"26190b",x"23170a",x"23170a",x"23170b",x"26190d",x"2f1f0f",x"23190f",x"271b0e",x"2a1c0f",x"271a0e",x"2d1f11",x"322212",x"3a2712",x"302111",x"2f2011",x"322211",x"2b1e0f",x"2f200f",x"291c0f",x"2d1f0f",x"312010",x"2f200f",x"382511",x"382510",x"372310",x"3c2711",x"36230f",x"3a2713",x"392712",x"322212",x"312010",x"302111",x"352413",x"342314",x"342313",x"322213",x"352515",x"382616",x"352516",x"392716",x"362616",x"3b2916",x"362617",x"372615",x"362516",x"362617",x"382719",x"332519",x"342416",x"362719",x"332517",x"2f2115",x"302318",x"2e2218",x"2b2015",x"312417",x"302318",x"302318",x"372719",x"362719",x"312318",x"322417",x"332519",x"322418",x"342517",x"302215",x"2f2317",x"2e2217",x"312417",x"2d2117",x"302417",x"2f2317",x"2d2216",x"302318",x"2e2216",x"302317",x"2f2318",x"2d2116",x"2b2016",x"2c2015",x"2e2115",x"2f2317",x"2c2117",x"2e2216",x"332416",x"302214",x"2e2115",x"2d2115",x"2d2115",x"2c2116",x"291d12",x"2c2014",x"271d13",x"291e14",x"261c13",x"2a1e11",x"2a1e12",x"2d2013",x"251b12",x"251b11",x"211910",x"21180f",x"231a11",x"241a10",x"241a10",x"2d1e10",x"2c1d10",x"2b1d0f",x"31200f",x"2e1f0f",x"2f1f10",x"281c0f",x"25180d",x"2b1d0d",x"23190d",x"2c1d0d",x"2a1c0d",x"291c0d",x"24180c",x"271a0d",x"24180c",x"24190d",x"22180d",x"1f150d",x"171009",x"1d130a",x"1b120a",x"1b120a",x"171009",x"1b1209",x"1f1408",x"1c1208",x"191007",x"180f07",x"201408",x"201508",x"19110a",x"1b1209",x"1b130a",x"21160b",x"181007",x"211508",x"1c130a",x"1b1209",x"24180d",x"1b130b",x"18110a",x"17110a",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"331d0d",x"2b180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"180f07",x"150e07",x"150e07",x"1e1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"27170a",x"2d1a0c",x"2b190b",x"2a180b",x"27160a",x"251509",x"211309",x"221309",x"281609",x"221308",x"201208",x"231409",x"201309",x"1b1108",x"201309",x"27160a",x"251509",x"231509",x"29170a",x"251509",x"241409",x"25150a",x"27160a",x"2a180b",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"535353",x"545454",x"575757",x"515151",x"424242",x"3e3e3e",x"3c3c3c",x"363636",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d4d4d",x"3e3e3e",x"3a3a3a",x"363635",x"000000",x"000000",x"3e3e3e",x"404040",x"3f3f3f",x"404040",x"393939",x"323232",x"333333",x"2c2c2c",x"313131",x"322f2d",x"303030",x"2f2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"343434",x"393939",x"3f3f3f",x"3a3a3a",x"343434",x"353535",x"3b3b3b",x"323232",x"323232",x"2f2f2f",x"373737",x"3c3c3c",x"323232",x"333333",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211a14",x"211a14",x"1e1811",x"1e1811",x"1f1912",x"1f1811",x"1d160f",x"1c160f",x"1b150e",x"19130c",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1408",x"160f07",x"1c1208",x"1f1408",x"241708",x"1d1208",x"241608",x"261809",x"291a09",x"27190c",x"26190b",x"25170a",x"25190a",x"20160d",x"21170d",x"291b0e",x"291b0f",x"2c1e10",x"302010",x"382411",x"3b2711",x"291c0f",x"2b1d0f",x"342311",x"2e1f10",x"332210",x"2d1f0f",x"39250f",x"3a250f",x"34220e",x"412a10",x"3e2910",x"38250f",x"32210e",x"302011",x"312110",x"3b2711",x"352310",x"2f2010",x"2b1e11",x"362412",x"312213",x"332313",x"312214",x"342413",x"342415",x"322313",x"382614",x"362617",x"382817",x"312315",x"352616",x"332417",x"332517",x"332415",x"2d2015",x"2f2216",x"2e2217",x"2e2217",x"2b2017",x"2b2016",x"292017",x"291f16",x"2d1f15",x"2a2017",x"292016",x"2f2318",x"2f2318",x"2e2116",x"302317",x"2f2216",x"2f2317",x"302316",x"2f2317",x"2a2016",x"2e2217",x"302418",x"2a2016",x"2e2217",x"2e2318",x"291f15",x"2a1f15",x"2c2116",x"2d2115",x"2d2216",x"2a2015",x"292016",x"2b1f13",x"2e2014",x"2c2015",x"2a2015",x"2b2116",x"2f2317",x"302216",x"2e2216",x"2c2115",x"2a1e13",x"2c1f13",x"2c2014",x"2c2014",x"251b11",x"261c12",x"241b11",x"2b1f12",x"281d12",x"261b10",x"241a10",x"241a10",x"211810",x"221911",x"231910",x"1f170e",x"21180f",x"281c0f",x"2b1d0f",x"281b0d",x"2e1f0e",x"291c0d",x"2a1d0d",x"25180d",x"22170c",x"2a1c0d",x"22170c",x"2a1c0d",x"271a0c",x"281b0d",x"22160b",x"24180b",x"21160a",x"21170a",x"1e150a",x"1c130a",x"19110a",x"1d130b",x"171009",x"25190b",x"1b1209",x"181007",x"1c1208",x"1c1208",x"1a1107",x"1c1208",x"221608",x"1b1108",x"170f07",x"181007",x"231608",x"160e07",x"150e07",x"1d1308",x"1a1107",x"1a1107",x"1f150b",x"1c130a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"150e07",x"150e07",x"150e07",x"4e4133",x"4d4032",x"493d2f",x"504335",x"46392d",x"534235",x"5c4d3f",x"4f4134",x"4d4034",x"534234",x"4b3c2f",x"4c3d2f",x"180f07",x"150e07",x"150e07",x"1e1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"27170a",x"2d1a0c",x"2b190b",x"2a180b",x"27160a",x"251509",x"211309",x"221309",x"281609",x"221308",x"201208",x"231409",x"201309",x"1b1108",x"201309",x"27160a",x"251509",x"231509",x"29170a",x"251509",x"241409",x"25150a",x"27160a",x"2a180b",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"515151",x"4a4a4a",x"424242",x"3e3e3e",x"373737",x"333333",x"41230f",x"3c200e",x"3e210e",x"40220e",x"40220e",x"41240f",x"41230f",x"41240f",x"3f220e",x"41240f",x"412410",x"432510",x"40230f",x"40230f",x"000000",x"000000",x"000000",x"3f3f3f",x"404040",x"393939",x"323232",x"333333",x"303030",x"313131",x"322f2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"353535",x"383838",x"3b3b3b",x"323232",x"323232",x"323232",x"000000",x"3c3c3c",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1811",x"1e1811",x"1f1912",x"1f1912",x"201912",x"1e1711",x"1d1610",x"1d1710",x"1c150e",x"19130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"231608",x"180f07",x"1b1108",x"160f07",x"181007",x"170f07",x"1d1308",x"1e1308",x"231608",x"26190b",x"20150a",x"1a120a",x"24170a",x"26190c",x"25190d",x"2d1d0e",x"291b0e",x"31200e",x"35220e",x"362310",x"2f1f0e",x"2b1c0e",x"33210e",x"34220e",x"31210f",x"32200e",x"33210e",x"33210e",x"3b270f",x"412b11",x"3b260f",x"34220e",x"2f1f0e",x"38250f",x"2b1d0e",x"312110",x"342310",x"312110",x"24190f",x"302112",x"382613",x"322212",x"2f2013",x"362513",x"2f2113",x"302214",x"2e2115",x"342415",x"322314",x"382614",x"2c2015",x"2f2316",x"312316",x"2e2217",x"2a2016",x"2b2016",x"281e15",x"271d15",x"261d15",x"261d14",x"241c13",x"251d15",x"281e16",x"251d14",x"261d15",x"271d13",x"2c2016",x"281e14",x"281d14",x"291f15",x"291e15",x"2a1f16",x"2a1f15",x"2a1f16",x"291f15",x"2d2115",x"281e16",x"291f15",x"2a1f14",x"281e14",x"271e15",x"271e15",x"2b2016",x"291f15",x"291f15",x"261d14",x"2a2015",x"2c2014",x"2b2016",x"291f15",x"281e14",x"2a1e13",x"2b1f14",x"2b1e13",x"2b1f13",x"291e14",x"291d12",x"281d12",x"2a1e13",x"261c13",x"241b12",x"241b12",x"241a0f",x"231a11",x"23180f",x"20180f",x"211911",x"1f170f",x"1e160e",x"1e160d",x"1d150e",x"20170e",x"23180d",x"26190d",x"271a0d",x"291c0d",x"26190d",x"291b0d",x"20150a",x"20150b",x"25180a",x"1e140b",x"281a0b",x"23170a",x"26190b",x"20160b",x"24180a",x"20160b",x"20150a",x"1e140a",x"1c130a",x"17100a",x"18110a",x"150e07",x"170f07",x"160f07",x"170f07",x"181007",x"170f07",x"191007",x"1b1108",x"160e07",x"170f07",x"160f07",x"1b1108",x"170f07",x"150e07",x"150e07",x"160f07",x"160f07",x"160f07",x"1a1107",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"4e4133",x"4e4133",x"4d4032",x"493d2f",x"504335",x"46392d",x"534235",x"5c4d3f",x"4f4134",x"48392d",x"534234",x"4b3c2f",x"4c3d2f",x"403429",x"4d3d30",x"493d2f",x"47392d",x"44392b",x"423628",x"45392c",x"473a2c",x"614a3b",x"5e4738",x"554234",x"5d483a",x"5c4738",x"5b483a",x"544637",x"403329",x"544738",x"5a493a",x"58493a",x"57493a",x"574a3a",x"504335",x"493f32",x"493c30",x"5d4a3b",x"544335",x"4a3c2f",x"5a4a3a",x"574537",x"564537",x"5b4a3b",x"5c4f3e",x"615444",x"5d4f3f",x"5b4d3e",x"604e3e",x"594b3b",x"594c3c",x"584a3a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381e0d",x"381e0d",x"3e220e",x"3e220e",x"41230f",x"3c200e",x"3e210e",x"40220e",x"41230f",x"41240f",x"41230f",x"41240f",x"3f220e",x"41240f",x"412410",x"432510",x"40230f",x"40230f",x"412410",x"41240f",x"412410",x"432511",x"462812",x"472812",x"472812",x"442611",x"482812",x"482912",x"4c2b14",x"472813",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1912",x"1f1912",x"1f1812",x"1f1912",x"1f1912",x"1d1710",x"1c150e",x"1b140d",x"1c150e",x"19130c",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"271809",x"150e07",x"17110a",x"17100a",x"1c1309",x"2b1b0b",x"20150a",x"19130c",x"1e150c",x"20160d",x"32200e",x"291c0d",x"24180c",x"26190d",x"22180d",x"2a1c0d",x"33210e",x"23180c",x"37230f",x"271a0d",x"2e1f0e",x"30200e",x"24180c",x"30200e",x"2f1f0e",x"2b1d0e",x"25180d",x"1d150b",x"281a0d",x"2a1d0f",x"1d160e",x"2c1d0f",x"2d1f11",x"2e2011",x"2d2011",x"302113",x"2b1e12",x"2a1f12",x"261c12",x"251c12",x"362515",x"2e2115",x"231b14",x"281e15",x"251c15",x"261d15",x"261d15",x"271e15",x"231b13",x"261e15",x"241d15",x"251d15",x"241c14",x"241c15",x"231c13",x"231c15",x"221c15",x"261c15",x"241c13",x"251d15",x"241d15",x"241c13",x"241b12",x"281f16",x"271d15",x"251d15",x"251c14",x"2a2016",x"251c14",x"271f15",x"271e15",x"271e15",x"241c14",x"281d13",x"271d13",x"261d15",x"271d13",x"241b13",x"261c13",x"281d13",x"281d14",x"251b12",x"261d14",x"291e15",x"281d13",x"281e14",x"2a1f14",x"271d13",x"251c12",x"231a12",x"271d12",x"241b12",x"231a12",x"21180f",x"211910",x"20180f",x"221911",x"1f1710",x"1c150e",x"1c150f",x"1c150e",x"1c150e",x"1c150e",x"1a130c",x"1e150c",x"1e160c",x"23170c",x"23170a",x"23170b",x"25190b",x"1c1309",x"1d130a",x"23170b",x"1b120a",x"25190a",x"20150b",x"25180b",x"20150b",x"23170b",x"20150a",x"1d130a",x"1c1309",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"594a3b",x"594a3b",x"483d30",x"44392d",x"524637",x"524638",x"534737",x"514134",x"42362a",x"483d30",x"4d3f31",x"45392c",x"43372b",x"403529",x"4a3e30",x"463b2d",x"473b2e",x"44392b",x"413528",x"45392c",x"463a2c",x"614a3b",x"5e4738",x"554234",x"5d483a",x"5c4738",x"5b483a",x"544637",x"403329",x"544738",x"5a493a",x"58493a",x"57493a",x"574a3a",x"504335",x"493f32",x"5d4b3d",x"5d4a3b",x"544335",x"4a3c2f",x"5a4a3a",x"574537",x"564537",x"5b4a3b",x"5c4f3e",x"615444",x"5d4f3f",x"5b4d3e",x"604e3e",x"594b3b",x"594c3c",x"584a3a",x"5c4b3b",x"504233",x"574838",x"5f4c3c",x"564838",x"534536",x"554838",x"564838",x"504335",x"584a3a",x"554838",x"514537",x"534637",x"574939",x"584839",x"564838",x"514335",x"514536",x"544738",x"4d4133",x"504335",x"514537",x"544538",x"5f4c3c",x"6c5242",x"6c5242",x"5f4e3e",x"664f3f",x"5e4d3c",x"604e3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1108",x"1d1108",x"261509",x"27160a",x"341d0d",x"381f0e",x"3a210e",x"3c220f",x"3b210e",x"3c210f",x"3e230f",x"3f230f",x"3e220f",x"432511",x"432510",x"452711",x"422410",x"3f220f",x"412410",x"41240f",x"412410",x"432511",x"462812",x"472812",x"452711",x"442611",x"482812",x"482912",x"4c2b14",x"472813",x"472813",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1912",x"1f1912",x"1f1811",x"1f1812",x"1f1812",x"1d160f",x"1d160f",x"1b140d",x"19130c",x"19120b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"17110a",x"17110a",x"171009",x"171009",x"19110a",x"1a120a",x"1b130b",x"1c140c",x"1a140c",x"271a0c",x"20170d",x"26190d",x"1f150d",x"1b1209",x"1d140a",x"1c1309",x"20150a",x"1f140a",x"1d130a",x"1d130a",x"1d130b",x"1d130a",x"1b140c",x"1c140c",x"1c130b",x"1b140c",x"1d150e",x"1c150e",x"1c150d",x"1d170f",x"1e170f",x"1d170f",x"211a12",x"221911",x"201810",x"211912",x"221b14",x"221b14",x"221b13",x"231b14",x"211913",x"221b13",x"211a12",x"221b13",x"221b14",x"241c14",x"231b14",x"221b14",x"221b14",x"211b13",x"201911",x"201913",x"201912",x"231b13",x"231b14",x"221b13",x"211a13",x"221a12",x"231b14",x"302316",x"241c14",x"211a13",x"211912",x"241b13",x"221a12",x"251c13",x"251c14",x"251c14",x"231b13",x"231b12",x"251b12",x"241b13",x"251c13",x"231b12",x"261d15",x"271d14",x"271d15",x"241b13",x"251c14",x"241a12",x"241a11",x"261c13",x"271c13",x"241b13",x"251b12",x"231b12",x"271d13",x"221911",x"21180f",x"20170f",x"271c11",x"201810",x"20170e",x"1c150d",x"1c150e",x"1c150e",x"1c150e",x"1a130b",x"19120b",x"19130c",x"1c140b",x"1a1209",x"1c130a",x"1e140a",x"1b130a",x"21160a",x"191109",x"1a120a",x"22160b",x"1b120a",x"25180b",x"1e140b",x"23170b",x"1c1208",x"201408",x"1c1208",x"1b1108",x"1a1107",x"181007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"5b4a3b",x"5b4a3b",x"5e4d3d",x"594a3b",x"544738",x"5e513f",x"5c4e3e",x"544738",x"4d4032",x"584a3b",x"504335",x"504234",x"544738",x"4a3e32",x"574838",x"4e4034",x"554637",x"4a3d31",x"4c4033",x"3d3227",x"493d2e",x"493d2f",x"4d4032",x"594838",x"584738",x"5f4c3c",x"5a4a3b",x"594a3b",x"5c4b3b",x"514335",x"534638",x"594c3c",x"5b4d3c",x"604f3f",x"615040",x"4f4133",x"524436",x"5c4f3e",x"564a3b",x"5d4f3f",x"564738",x"5f4f3f",x"56493a",x"594b3c",x"5a4e3d",x"5e5140",x"5f5242",x"5d5040",x"5c503f",x"635140",x"5c4e3e",x"594c3c",x"5a4b3b",x"5c4b3b",x"504233",x"574838",x"5c4b3c",x"564838",x"534536",x"554838",x"564939",x"504335",x"584a3a",x"554838",x"4a3e30",x"534637",x"574939",x"584839",x"564838",x"514335",x"514536",x"544738",x"4d4133",x"504335",x"514537",x"544538",x"5f4c3c",x"6c5242",x"6c5242",x"5f4e3e",x"664f3f",x"5e4d3c",x"604e3f",x"5d4d3c",x"5e4c3d",x"4b3c2f",x"574938",x"5a4a3b",x"5b4839",x"594a3a",x"5c4b3b",x"534536",x"544638",x"5a4a3b",x"5d4b3b",x"594939",x"624d3d",x"534435",x"574939",x"574939",x"584a39",x"574939",x"5d4f3e",x"624d3d",x"594838",x"574335",x"45362a",x"523f32",x"634e3e",x"624d3e",x"614e3e",x"564b3b",x"5b4e3e",x"5e4d3d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1e1208",x"1d1208",x"201309",x"241509",x"29170b",x"2d190b",x"311c0d",x"351e0e",x"37200e",x"37200e",x"371e0d",x"351e0d",x"351d0d",x"3b210f",x"3a200f",x"341c0c",x"351d0d",x"341d0c",x"331c0c",x"321c0c",x"341d0d",x"301b0c",x"321d0d",x"301c0d",x"2d190c",x"2b190b",x"301b0c",x"2f1b0d",x"3b2210",x"351f0e",x"351f0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1811",x"1f1811",x"1f1812",x"1d1710",x"1d160f",x"1e1711",x"1e1711",x"1b140d",x"19120b",x"17100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"171009",x"171009",x"181109",x"191109",x"181109",x"191109",x"181109",x"1b120a",x"181009",x"1a1109",x"1c130a",x"1a1209",x"1b1209",x"1a1209",x"1c1309",x"1d130a",x"1b1209",x"1b120a",x"1b1209",x"1c1309",x"191109",x"1c140c",x"1b130b",x"1b140c",x"1a130b",x"1c150e",x"1c160e",x"1c150e",x"1e1710",x"1e1710",x"1d170f",x"1f1811",x"201911",x"201912",x"201912",x"201912",x"201912",x"211912",x"201912",x"201912",x"211a13",x"221b13",x"221b14",x"231b13",x"211912",x"211a13",x"221b14",x"211a14",x"211b14",x"201912",x"201a13",x"231b14",x"221b14",x"211a13",x"201912",x"221a13",x"211912",x"221a13",x"221a12",x"211a13",x"201a12",x"241c14",x"231b14",x"231b13",x"241b13",x"241c13",x"221b13",x"241c14",x"251c13",x"211911",x"231a12",x"211911",x"211910",x"241b13",x"241b12",x"221911",x"221911",x"231a12",x"231a12",x"241b12",x"251c12",x"231a12",x"231a12",x"201810",x"23180f",x"211910",x"20170f",x"1f1810",x"1e160e",x"1e160e",x"1e160e",x"1c150d",x"1c140d",x"19120b",x"1a130c",x"1a130c",x"19130c",x"17110a",x"19110a",x"1a110a",x"1b1209",x"1c1309",x"19110a",x"1f150a",x"18110a",x"180f07",x"1f1408",x"181007",x"221508",x"1b1108",x"201408",x"1b1108",x"1e1308",x"1c1208",x"1a1107",x"191007",x"181007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"5b4c3d",x"544537",x"453a2d",x"453a2d",x"4a3f31",x"544738",x"5a4b3b",x"58493a",x"56483a",x"604e3e",x"5b4c3c",x"564839",x"584a3b",x"5c4d3d",x"5d4c3d",x"58493a",x"594739",x"554537",x"534336",x"574839",x"5e4d3d",x"5e4d3d",x"5f4d3e",x"5a4b3b",x"58493a",x"4a3e30",x"504536",x"524637",x"544838",x"574839",x"4f4334",x"584a3b",x"554536",x"604e3e",x"5d4d3d",x"514536",x"5b4e3e",x"5d503f",x"5a4c3c",x"574a39",x"514536",x"514335",x"644d3e",x"675040",x"6a5141",x"634f3f",x"65503f",x"614e3e",x"625444",x"5c4e3d",x"5a4a3b",x"5f4d3e",x"594839",x"514134",x"5c4a3c",x"5d4c3c",x"5f4d3e",x"5c4a3b",x"5c4a3a",x"604d3e",x"554638",x"5c4e3d",x"5d4d3d",x"5e4d3d",x"594a3a",x"5a4a3b",x"5c4a3b",x"5d4b3b",x"564738",x"524436",x"554636",x"4f4233",x"564838",x"5a4a3b",x"5b4b3c",x"5e4c3d",x"5f4e3d",x"614f3f",x"644e3f",x"664f3f",x"5e4d3c",x"604e3e",x"5c4c3d",x"5e4c3d",x"4b3c2f",x"574938",x"574435",x"5b4839",x"594a3a",x"5c4b3b",x"534536",x"544638",x"5a4a3b",x"5d4b3b",x"594939",x"624d3d",x"534435",x"574939",x"574939",x"584a39",x"574939",x"5d4f3e",x"624d3d",x"594838",x"574335",x"45362a",x"523f32",x"634e3e",x"624d3e",x"614e3e",x"564b3b",x"5b4e3e",x"5e4d3d",x"5c4d3c",x"594a3a",x"5b4a3b",x"5c493a",x"634e3e",x"534335",x"554738",x"43382c",x"4f3f32",x"5b493a",x"574637",x"4f4030",x"544335",x"544335",x"564334",x"4f4131",x"46382b",x"4a3d2e",x"574a3b",x"4e4031",x"493b2e",x"463a2d",x"534334",x"564536",x"514334",x"4d4032",x"554435",x"534334",x"5d4a3b",x"5d4c3c",x"604e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1209",x"1f1209",x"1f1309",x"221409",x"27160a",x"2d190b",x"311b0c",x"351f0e",x"371f0e",x"371f0d",x"371f0d",x"371e0d",x"381f0d",x"3c210f",x"3b210f",x"3c210f",x"3e230f",x"3d220f",x"3c220f",x"3b210f",x"3d2310",x"38200e",x"341d0d",x"351f0e",x"321c0d",x"311c0d",x"2b180b",x"29180b",x"27170b",x"24150a",x"221409",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1d1610",x"1d1610",x"1d1610",x"1d1610",x"1c150e",x"1b150e",x"1a130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"171009",x"18110a",x"181109",x"181009",x"18110a",x"181009",x"19110a",x"17110a",x"18110a",x"19110a",x"191109",x"19110a",x"19110a",x"1a120a",x"1a1209",x"1a1109",x"1a110a",x"1a110a",x"1b1209",x"19110a",x"191109",x"18110a",x"1a140c",x"1a130c",x"19130c",x"1c150e",x"1c150e",x"1c150e",x"1d160f",x"1e1610",x"1d170f",x"201912",x"201811",x"1f1811",x"1f1911",x"1f1811",x"201912",x"1e1711",x"1f1811",x"201912",x"201911",x"201912",x"211911",x"211912",x"201912",x"1f1911",x"1f1811",x"1f1811",x"201912",x"201a13",x"231b14",x"211b13",x"211a13",x"1f1811",x"201811",x"1f1911",x"1f1811",x"201911",x"201912",x"201812",x"211a12",x"201911",x"211911",x"221a12",x"221a12",x"201912",x"211912",x"231b12",x"221a12",x"221911",x"211a12",x"211810",x"221911",x"231b12",x"211911",x"211911",x"211911",x"221911",x"221a12",x"221911",x"201811",x"201810",x"1f1710",x"211910",x"201810",x"1f170f",x"1d150e",x"1d160e",x"1d150e",x"1d150e",x"1a130c",x"1a130c",x"1a130c",x"1a120b",x"18110a",x"171009",x"171009",x"191109",x"191109",x"1a1209",x"191007",x"170f07",x"1c1208",x"160e07",x"170f07",x"1e1308",x"181007",x"201508",x"1a1107",x"1f1408",x"1a1107",x"1d1308",x"1b1108",x"191007",x"191007",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"43372a",x"453a2d",x"453a2d",x"4a3f31",x"574a3a",x"5a4b3b",x"58493a",x"56483a",x"5b4c3d",x"5b4c3c",x"564839",x"584a3b",x"5c4d3d",x"5d4c3d",x"58493a",x"594739",x"554537",x"534336",x"574839",x"5e4d3d",x"5e4d3d",x"5f4d3e",x"5a4b3b",x"58493a",x"504134",x"58493a",x"514436",x"544838",x"564838",x"584a3b",x"5e4c3d",x"604b3b",x"624e3f",x"5f4c3d",x"614d3e",x"5e4e3d",x"5e4d3e",x"5e4e3e",x"594c3d",x"5b4e3d",x"57493a",x"594c3d",x"5a493a",x"605242",x"635443",x"625242",x"5f4f3f",x"665646",x"675645",x"685645",x"635442",x"605342",x"645343",x"625141",x"635141",x"5f4e3e",x"5f4f3e",x"5c4e3d",x"594b3c",x"4f4435",x"5a4d3d",x"594d3c",x"584b3b",x"604f40",x"5c4b3c",x"674f40",x"614f3e",x"604e3e",x"5b4a3b",x"534637",x"584a3a",x"5b4c3d",x"5f4f3f",x"5c4f3f",x"514134",x"4f4033",x"584b3c",x"584b3b",x"5b4c3c",x"5a493a",x"574838",x"5c4b3b",x"59493a",x"4f3e32",x"5e4a3b",x"5e4b3b",x"5c4939",x"5b4838",x"604b3c",x"5a4a3a",x"5b4b3b",x"5d4b3b",x"5e4c3b",x"5a4a3a",x"5c4c3b",x"594a39",x"59493a",x"5a4b3a",x"5b4c3b",x"645443",x"5c4e3d",x"5b4b3b",x"514435",x"4a3c2f",x"513f32",x"4f3d31",x"5c4c3c",x"5d4d3c",x"5c4d3d",x"54493a",x"594c3d",x"5e4d3d",x"5c4d3c",x"594a3a",x"5b4a3b",x"5c493a",x"634e3e",x"534335",x"554738",x"43382c",x"4f3f32",x"5b493a",x"574637",x"4f4030",x"544335",x"544335",x"564334",x"4f4131",x"46382b",x"4a3d2e",x"574a3b",x"4e4031",x"493b2e",x"463a2d",x"534334",x"564536",x"514334",x"4d4032",x"554435",x"594838",x"5d4a3b",x"5d4c3c",x"604e3e",x"624f3f",x"645040",x"614e3f",x"514437",x"554739",x"5a4738",x"5f4a3b",x"5a4739",x"5e4a3a",x"6b5040",x"6c5141",x"684f3f",x"1e1208",x"1f1208",x"231409",x"271509",x"29170a",x"2d190a",x"2f1a0b",x"311a0b",x"321b0b",x"331b0b",x"351d0c",x"381f0d",x"3b210f",x"3e220f",x"3e230f",x"3c210f",x"3b210e",x"39200e",x"381f0d",x"351d0c",x"371e0d",x"3c220f",x"371f0e",x"37200e",x"341e0d",x"2f1b0c",x"2d1a0c",x"28170a",x"27170b",x"231509",x"231509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1d1710",x"1d1710",x"1c150f",x"1b150e",x"1b140d",x"19130c",x"1a130c",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"171009",x"17100a",x"171009",x"171009",x"17110a",x"17110a",x"17100a",x"17110a",x"171009",x"17110a",x"17110a",x"17110a",x"181109",x"181109",x"18110a",x"18110a",x"181109",x"19110a",x"181109",x"181109",x"18110a",x"18110a",x"1a130c",x"19120b",x"1a130c",x"1c150e",x"1c140d",x"1c150e",x"1e1711",x"1d160f",x"1e1810",x"1d160f",x"1f1711",x"201912",x"1f1911",x"1e1710",x"1e1711",x"1f1912",x"1f1711",x"201912",x"1f1911",x"201911",x"1f1911",x"201812",x"201912",x"1e1711",x"1f1811",x"1f1811",x"1f1811",x"201811",x"1e1811",x"1f1811",x"1e1710",x"201912",x"1f1912",x"1f1812",x"1f1812",x"1f1912",x"1f1811",x"1f1911",x"1f1811",x"1f1911",x"1f1811",x"1f1810",x"201912",x"201811",x"201911",x"211912",x"211912",x"211911",x"1f1811",x"1e170f",x"201810",x"1e170f",x"1f1710",x"1e1710",x"1e1710",x"1e1710",x"201810",x"1f1710",x"1f1710",x"1e1711",x"1e170f",x"1d150e",x"1c150e",x"1c150e",x"1c150e",x"1c150e",x"1a130c",x"1a140c",x"1a130c",x"19130c",x"17110a",x"171009",x"171009",x"171009",x"170f07",x"170f07",x"180f07",x"191007",x"160f07",x"1b1108",x"160e07",x"170f07",x"1c1208",x"180f07",x"1f1408",x"1a1107",x"1d1308",x"191007",x"1c1208",x"1a1107",x"181007",x"181007",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"504134",x"58493a",x"514436",x"554638",x"564838",x"584a3b",x"5e4c3d",x"5f4c3d",x"624e3f",x"5f4c3d",x"614d3e",x"5e4e3d",x"5e4d3e",x"5e4e3e",x"594c3d",x"5b4e3d",x"57493a",x"594c3d",x"5a493a",x"605242",x"635443",x"625242",x"5f4f3f",x"665646",x"675645",x"685645",x"635442",x"605342",x"645343",x"625141",x"635141",x"5e4f3f",x"635443",x"5e503f",x"615142",x"5e5041",x"625644",x"625443",x"625242",x"605342",x"5e5140",x"5d5040",x"56493b",x"56483a",x"5b4c3d",x"5a4d3d",x"594b3c",x"5b4f3e",x"605242",x"5a4d3d",x"5d5040",x"615443",x"645443",x"5e5241",x"615242",x"5d5040",x"605343",x"5d4e3e",x"5c4e3d",x"5c4f3e",x"5d4e3e",x"5c4d3d",x"5b4839",x"5a4939",x"544637",x"564838",x"564839",x"574a3a",x"624e3e",x"624f3f",x"5b4c3c",x"5a4c3b",x"5d4d3c",x"574a3b",x"5e4d3d",x"614e3e",x"5d4e3d",x"5e4d3d",x"5f4d3d",x"4c3d30",x"5e4c3d",x"5a4c3b",x"5b4c3b",x"5b4b3a",x"524334",x"514234",x"5e4f3e",x"5c4d3d",x"584a3a",x"5c4c3c",x"5c4c3c",x"5e4d3d",x"594a3a",x"574939",x"5b4b3a",x"4c3f31",x"4c3f31",x"594a3a",x"584737",x"524334",x"574536",x"5a4636",x"4c3f30",x"4c3e2f",x"564434",x"504334",x"473a2d",x"423528",x"4b3e30",x"4c3f31",x"4d4031",x"504334",x"514232",x"5d493a",x"5b4839",x"584838",x"5d4a3b",x"5d4b3b",x"604e3e",x"624f3f",x"645040",x"614e3f",x"514437",x"554739",x"5a4738",x"5f4a3b",x"5a4739",x"5e4a3a",x"6b5040",x"6c5141",x"684f3f",x"4e4234",x"211309",x"26150a",x"29170a",x"2f1a0b",x"301b0b",x"2f190b",x"301a0b",x"321a0b",x"361d0c",x"371e0d",x"3a1f0e",x"3b200e",x"3d210f",x"3e220f",x"3e230f",x"3e230f",x"3e220f",x"412511",x"3f2310",x"3c210e",x"351d0b",x"381f0d",x"341d0c",x"331c0c",x"291709",x"2d1a0b",x"2b190b",x"27170b",x"27170b",x"27170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1e1711",x"1d1610",x"1b150e",x"1b150e",x"1b150e",x"19120c",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"17110a",x"171009",x"171009",x"17110a",x"18110a",x"17110a",x"17110a",x"171009",x"17100a",x"171009",x"171009",x"160f07",x"160e07",x"160e07",x"150e07",x"160e07",x"160f07",x"181009",x"181009",x"181009",x"18100a",x"1a130c",x"1a130c",x"19120c",x"19130c",x"1c150f",x"1b140e",x"1b140d",x"1d160f",x"1d160f",x"1e1710",x"1e1710",x"1d160f",x"1d160f",x"1e1610",x"1f1811",x"1f1811",x"1f1811",x"1f1710",x"1f1710",x"1f1911",x"201812",x"201912",x"1f1912",x"201912",x"1f1912",x"201913",x"1f1811",x"201913",x"1f1812",x"1f1811",x"1f1912",x"1f1811",x"1f1811",x"1d1710",x"1d1610",x"1d1610",x"1d1710",x"1e1710",x"1c150e",x"1e1810",x"1d160f",x"1f1710",x"1e1710",x"1d170f",x"1e1710",x"1d170f",x"1f1811",x"1e1710",x"1e1710",x"1d160f",x"1e170f",x"1d170f",x"1e170f",x"1e1711",x"1d170f",x"1e1811",x"1f1710",x"1e1811",x"1c150d",x"1c150e",x"1c160e",x"1c160e",x"1c150d",x"1c150e",x"19120b",x"1a130c",x"19120c",x"1a130c",x"19120c",x"171009",x"17110a",x"18110a",x"17110a",x"150e07",x"160f07",x"160f07",x"170f07",x"180f07",x"160f07",x"1a1107",x"150e07",x"160f07",x"1b1108",x"170f07",x"1d1308",x"191007",x"1c1208",x"181007",x"1b1108",x"191007",x"180f07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e4f3f",x"635443",x"5e503f",x"615142",x"5e5041",x"625644",x"625443",x"625242",x"605342",x"5e5140",x"5d5040",x"56493b",x"56483a",x"5b4c3d",x"5a4d3d",x"594b3c",x"5b4f3e",x"605242",x"5a4d3d",x"5d5040",x"615443",x"645443",x"5e5241",x"615242",x"5d5040",x"605343",x"625141",x"5c4e3d",x"5c4f3e",x"5d4e3e",x"605140",x"5c4d3e",x"5a4d3d",x"5f4d3e",x"5b4b3c",x"5d4c3d",x"5f4d3d",x"5d4c3d",x"5b4c3d",x"5b4d3d",x"5b4c3d",x"635142",x"625443",x"645242",x"665343",x"605242",x"635444",x"605041",x"655545",x"635343",x"655343",x"615040",x"5f5040",x"605242",x"605040",x"574839",x"5e4f3f",x"61503f",x"5f503f",x"615141",x"635141",x"635141",x"614c3c",x"654f3f",x"614b3c",x"5a4b3a",x"594c3c",x"594b3b",x"594d3c",x"594c3c",x"5b4f3f",x"57493a",x"57493a",x"564839",x"574839",x"614c3d",x"5f4c3c",x"604b3c",x"5f4b3b",x"604c3c",x"5b4a3a",x"614c3c",x"59483a",x"5a4838",x"624c3c",x"614c3d",x"594b3c",x"594c3c",x"5f4d3d",x"5c4c3c",x"604e3e",x"594a3b",x"5d4a3c",x"594638",x"514436",x"514436",x"534738",x"554737",x"5f4a3b",x"5e493a",x"4f4234",x"26160a",x"2c190b",x"321d0d",x"37200f",x"3b2210",x"3f2511",x"402511",x"3e2310",x"3d210f",x"3d210f",x"3c210e",x"3c210e",x"3c210e",x"402410",x"422511",x"412410",x"3f2410",x"402411",x"3f2410",x"331c0b",x"351d0c",x"381f0d",x"361e0c",x"331c0c",x"2f1a0b",x"2c180a",x"261609",x"28180b",x"28180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1c160f",x"1b150e",x"1b150e",x"1b140d",x"1a130c",x"19120c",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"261809",x"1c1007",x"1e1308",x"1a1008",x"1d1108",x"201309",x"231509",x"24150a",x"26160a",x"25150a",x"25150a",x"241509",x"231409",x"241509",x"251509",x"241409",x"221409",x"221409",x"221409",x"231409",x"221409",x"211409",x"211409",x"1e1208",x"1d1108",x"1c1108",x"1a1008",x"190f07",x"190f07",x"1a1008",x"1c1108",x"1d1208",x"1d1208",x"1e1208",x"1f1209",x"201309",x"211309",x"231409",x"25150a",x"24150a",x"26160a",x"26160a",x"25160a",x"25150a",x"25160a",x"24150a",x"24150a",x"24150a",x"241509",x"231509",x"231409",x"211309",x"1f1208",x"1f1208",x"1e1108",x"1e1208",x"1c1108",x"1e1208",x"1d1108",x"1c1108",x"1f1208",x"1c1108",x"1c1108",x"1e1208",x"1c1108",x"1b1108",x"1b1008",x"1a1008",x"190f08",x"180f07",x"150e07",x"17100a",x"171009",x"17100a",x"181009",x"171009",x"181009",x"181009",x"181009",x"181109",x"181009",x"181109",x"18110a",x"181109",x"181109",x"181109",x"181009",x"181109",x"181009",x"170f09",x"28170b",x"28170b",x"22140a",x"231509",x"271809",x"2b1b0a",x"171009",x"181009",x"161009",x"160f08",x"160f08",x"160f08",x"170f08",x"150e08",x"150e08",x"150e08",x"150e08",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"181007",x"170f07",x"191007",x"180f07",x"180f07",x"170f07",x"180f07",x"170f07",x"160f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c4d3e",x"5a4d3d",x"5f4d3e",x"5b4b3c",x"5d4c3d",x"5f4d3d",x"5d4c3d",x"5b4c3d",x"5b4d3d",x"5b4c3d",x"635142",x"625443",x"645242",x"665343",x"605242",x"635444",x"605041",x"655545",x"665645",x"655343",x"615040",x"5f5040",x"615141",x"605040",x"574839",x"5e4f3f",x"625141",x"5f503f",x"615141",x"635141",x"635444",x"645141",x"675343",x"645141",x"645242",x"655443",x"645242",x"655342",x"615040",x"5d4e3e",x"5a4b3c",x"5e4d3d",x"5f4e3f",x"5a4a3b",x"5a4b3c",x"635242",x"605141",x"635342",x"645543",x"5e503f",x"605040",x"5f5141",x"534436",x"605040",x"635040",x"635041",x"5d4e3e",x"5e5041",x"645343",x"665343",x"665243",x"59493a",x"5c493a",x"624d3c",x"654e3e",x"5e4a3b",x"614b3c",x"624c3d",x"5e4b3b",x"5d4a3a",x"241509",x"2a180b",x"2e1a0c",x"321c0d",x"39200f",x"3d2310",x"3c220f",x"3d220f",x"3f230f",x"3e220f",x"412410",x"3c200e",x"412410",x"40230f",x"3d210e",x"3e220f",x"412410",x"402410",x"422611",x"371e0c",x"371e0c",x"391f0d",x"2f1a0b",x"2b180a",x"2c180a",x"2d190b",x"29170a",x"231408",x"28170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1c150e",x"1c150e",x"1b150e",x"1a130c",x"19120b",x"171009",x"17100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"321f0a",x"311e0a",x"251708",x"241609",x"1d1208",x"1c1108",x"1d1208",x"211409",x"24150a",x"26170a",x"28170b",x"29180b",x"2a180b",x"29180b",x"29180b",x"29180b",x"27160a",x"26160a",x"25150a",x"241509",x"25160a",x"26160a",x"25160a",x"24150a",x"231509",x"221409",x"201208",x"1f1208",x"201308",x"201309",x"1f1208",x"201208",x"211309",x"211309",x"231409",x"241509",x"231409",x"231409",x"231409",x"201308",x"211308",x"271609",x"221308",x"221408",x"28170a",x"29180b",x"28170a",x"28170a",x"27170a",x"27160a",x"27170a",x"27160a",x"26160a",x"241509",x"221409",x"211309",x"201309",x"201309",x"1f1208",x"1f1309",x"1f1208",x"201309",x"1f1208",x"1f1208",x"211309",x"201309",x"201309",x"1e1208",x"1d1208",x"1c1108",x"1b1008",x"191008",x"180f07",x"150e07",x"150e07",x"17100a",x"181009",x"171009",x"181009",x"181009",x"181009",x"170f07",x"170f07",x"170f07",x"150e07",x"160e07",x"2b180b",x"28170a",x"181009",x"181109",x"512f16",x"3e2f24",x"482a13",x"28170b",x"27180b",x"26160a",x"2c1b0a",x"311e0b",x"2e1c09",x"2f1d0a",x"161009",x"160f08",x"160f08",x"533c2d",x"4c3b2e",x"5a473a",x"4e2c14",x"150e08",x"150e08",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"181007",x"170f07",x"191007",x"180f07",x"180f07",x"170f07",x"180f07",x"170f07",x"160f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"645141",x"675343",x"645141",x"645242",x"655443",x"645242",x"655342",x"615040",x"5d4e3e",x"5a4b3c",x"5e4d3d",x"5f4e3f",x"5a4a3b",x"5a4b3c",x"615342",x"605141",x"635342",x"645543",x"645545",x"605040",x"5f5141",x"534436",x"605040",x"635040",x"635041",x"5d4e3e",x"5e5041",x"645343",x"665343",x"665243",x"594a3c",x"604f3f",x"614f3f",x"644d3d",x"634e3e",x"604e3e",x"674e3f",x"604c3c",x"5f4e3e",x"201309",x"251509",x"2a180b",x"2d190b",x"311c0c",x"321c0c",x"361d0d",x"39200e",x"3a200e",x"3a200e",x"3a200e",x"3b210e",x"3d220f",x"3d220e",x"3f230f",x"3b210e",x"3d220f",x"3c210f",x"3d220f",x"3e2310",x"311a0a",x"321b0b",x"341d0c",x"311b0b",x"2e1a0b",x"2e190b",x"2e1a0b",x"2d190a",x"2d190a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"1b150e",x"1b140e",x"1a130c",x"1a130c",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"32200a",x"33200a",x"32200a",x"311f0a",x"261808",x"231609",x"1c1108",x"1b1108",x"1f1309",x"201309",x"26160a",x"28180b",x"29190c",x"2b1a0c",x"2b190c",x"2b190c",x"2b190b",x"2b190c",x"2a180b",x"28180b",x"26160a",x"251509",x"231409",x"25150a",x"26160a",x"25150a",x"25150a",x"241509",x"241509",x"231509",x"24150a",x"24150a",x"24150a",x"24150a",x"241509",x"241509",x"26160a",x"27170b",x"261509",x"261609",x"251509",x"27160a",x"271609",x"28170a",x"231408",x"271609",x"2c1a0c",x"2b190b",x"29180b",x"2a180b",x"29170a",x"29170b",x"29170b",x"29180b",x"29180b",x"27170a",x"241509",x"231409",x"211309",x"201309",x"201309",x"201309",x"201309",x"201309",x"201208",x"1f1208",x"211409",x"23150a",x"221409",x"211409",x"1e1208",x"1c1108",x"1c1108",x"1b1108",x"191008",x"170f07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"170f07",x"170f07",x"160e07",x"150e07",x"160e07",x"160e07",x"160e07",x"391e0d",x"4a2913",x"150e07",x"482a15",x"4c2d16",x"26170b",x"231509",x"311e0a",x"301e0b",x"301e0a",x"301f0a",x"2f1d0a",x"000000",x"2e1a0b",x"2e1a0b",x"150e07",x"3d220f",x"432611",x"432712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"625443",x"695443",x"615343",x"625141",x"615040",x"605141",x"5d4e3e",x"615443",x"605141",x"625140",x"614e3f",x"615443",x"635443",x"605343",x"605140",x"645443",x"615141",x"615242",x"554637",x"58493a",x"5b4d3d",x"5b4c3d",x"5c4d3d",x"605140",x"655544",x"625243",x"624f40",x"635141",x"685443",x"645141",x"5f4d3d",x"614f3f",x"5e503f",x"5e4d3d",x"615342",x"5e5141",x"5e5040",x"5d4f3f",x"5f5241",x"564a3b",x"605142",x"625141",x"635543",x"615242",x"615342",x"1b1108",x"624f3f",x"544738",x"27160a",x"2a180b",x"321c0d",x"321c0d",x"301c0c",x"321c0c",x"311b0c",x"311c0c",x"311c0c",x"321c0c",x"331d0d",x"351e0d",x"3b2210",x"3e2411",x"3c2310",x"3a200f",x"3b220f",x"3f2512",x"3f2511",x"3a200f",x"3a210e",x"341d0c",x"361f0d",x"321c0b",x"2e1a0b",x"2d1a0b",x"28170a",x"231509",x"211409",x"241609",x"241609",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150d",x"1b150d",x"1b150e",x"1c150e",x"19130c",x"19120b",x"1a130c",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"311f0a",x"32200a",x"32200a",x"301e0a",x"281909",x"211508",x"170f07",x"191008",x"1c1108",x"1e1208",x"221409",x"25160a",x"26160a",x"27170a",x"29180b",x"2a190b",x"2a190b",x"29190b",x"28170b",x"27170a",x"26160a",x"25150a",x"241509",x"25150a",x"26160a",x"25160a",x"26160a",x"26170a",x"26160a",x"27170b",x"26160a",x"25160a",x"25160a",x"28170b",x"2a190b",x"28170b",x"2a190b",x"26160a",x"29180b",x"28170b",x"231408",x"28170a",x"271609",x"28160a",x"28160a",x"271609",x"2a190b",x"29180b",x"29170b",x"27160a",x"27160a",x"271609",x"251509",x"251509",x"261509",x"251509",x"241509",x"231409",x"211309",x"201309",x"1e1208",x"1e1208",x"201309",x"201309",x"221409",x"211409",x"221509",x"221509",x"211409",x"201309",x"1d1208",x"1d1108",x"1c1108",x"1b1108",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"1a1107",x"191007",x"170f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"311d0d",x"482812",x"442611",x"492b14",x"150e07",x"452610",x"3b1f0d",x"1f1208",x"1c1008",x"241609",x"301d0b",x"33200a",x"301e0a",x"311f0a",x"32200a",x"1e1108",x"1e1108",x"150e07",x"331c0c",x"40220e",x"4a2b15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"655241",x"655242",x"675242",x"615342",x"615343",x"605443",x"5e5141",x"635242",x"634f40",x"665040",x"634e3f",x"655141",x"645040",x"5f4d3e",x"5b4a3b",x"584a3b",x"584a3a",x"534637",x"524637",x"5c4e3e",x"574b3c",x"5b4f3f",x"5c4f3f",x"615544",x"605142",x"615444",x"5c5041",x"5e5041",x"615343",x"5f5344",x"5c4e3f",x"625443",x"695443",x"615343",x"604f3f",x"615040",x"605141",x"5d4e3e",x"615443",x"605141",x"625140",x"614e3f",x"615443",x"635443",x"605343",x"605140",x"645443",x"615141",x"615242",x"554637",x"58493a",x"5b4d3d",x"5b4c3d",x"5c4d3d",x"605140",x"655544",x"625243",x"624f40",x"635141",x"685443",x"645141",x"5f4d3d",x"4f4234",x"514435",x"5b493a",x"624c3c",x"504234",x"231c16",x"241d17",x"261f19",x"241d17",x"201a13",x"1d1710",x"17110a",x"150e07",x"170f07",x"1a1108",x"1e1209",x"26160a",x"2b1a0c",x"2e1b0d",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"311c0c",x"311c0d",x"331d0d",x"351e0d",x"38200e",x"3a210f",x"3b210f",x"3a210f",x"3c210f",x"3c210f",x"3c220f",x"3c220f",x"3b210f",x"3b220f",x"3f2511",x"3a220f",x"38200e",x"331d0c",x"331d0d",x"301c0c",x"2b1a0b",x"25160a",x"221509",x"201308",x"201308",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b140d",x"19120b",x"19130c",x"1a130c",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1e0a",x"321f0a",x"32200a",x"2f1e0a",x"291a09",x"261809",x"211608",x"180f08",x"1a1008",x"1b1108",x"1e1209",x"22150a",x"27170b",x"27180b",x"28180b",x"27170a",x"27170a",x"29180b",x"29190b",x"28180b",x"27170b",x"25160a",x"25160a",x"25150a",x"25160a",x"25150a",x"251509",x"25160a",x"25160a",x"24150a",x"231509",x"241509",x"241509",x"25150a",x"26160a",x"27160a",x"27160a",x"29180b",x"29180b",x"29170b",x"28170a",x"28170a",x"2a180b",x"29180b",x"2b190b",x"29170b",x"2a180b",x"28170a",x"28160a",x"261509",x"261509",x"241409",x"241409",x"251509",x"251509",x"261609",x"261509",x"241509",x"231409",x"211309",x"1f1208",x"1f1208",x"1e1208",x"1f1208",x"201309",x"1f1208",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1d1108",x"1c1108",x"1a1008",x"1a1008",x"190f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"000000",x"1c1208",x"1c1308",x"170f07",x"191007",x"1f1408",x"170f07",x"160f07",x"3c210e",x"422510",x"472812",x"492912",x"2b190c",x"150e07",x"4a2b14",x"4e2e15",x"221409",x"1f1309",x"1b1108",x"2e1d09",x"33200a",x"32200a",x"32200a",x"33200a",x"1d1108",x"1d1108",x"150e07",x"1a1008",x"452610",x"452812",x"4a2c14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b3f32",x"4d3f32",x"524436",x"4b3d31",x"614f40",x"604f40",x"574839",x"5e4e3e",x"675242",x"645342",x"615141",x"645443",x"625443",x"605141",x"645746",x"615444",x"5d5141",x"5f5242",x"605241",x"605141",x"615343",x"554839",x"605241",x"615141",x"625040",x"655142",x"635343",x"615141",x"645242",x"625141",x"655241",x"655242",x"675242",x"615342",x"615343",x"605443",x"5e5141",x"5f5040",x"634f40",x"665040",x"634e3f",x"5f4c3c",x"645040",x"5f4d3e",x"5b4a3b",x"584a3b",x"584a3a",x"534637",x"524637",x"5c4e3e",x"574b3c",x"5b4f3f",x"5c4f3f",x"615544",x"605142",x"615444",x"5c5041",x"5e5041",x"615343",x"5f5344",x"5c4e3f",x"554535",x"584938",x"5b4a3a",x"5b4a3a",x"604c3c",x"5d4b3c",x"604c3c",x"624d3d",x"574839",x"604b3b",x"594838",x"5b493a",x"59493a",x"5b4b3b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"1b150e",x"1f1912",x"221c15",x"241d17",x"241d17",x"211a14",x"201a13",x"1d1710",x"19120b",x"150e07",x"160f07",x"1a1108",x"1e1309",x"24150a",x"29180b",x"2d1a0c",x"2d1a0b",x"2d1a0c",x"311c0d",x"321d0d",x"331d0d",x"341e0d",x"361f0e",x"39210f",x"3b220f",x"3c230f",x"3d220f",x"3c220f",x"3c210f",x"3d220f",x"412511",x"402511",x"3d2310",x"3c220f",x"3a210f",x"3c2310",x"3c2410",x"351e0d",x"321d0c",x"301c0c",x"2b1a0b",x"26160a",x"211308",x"211309",x"1c1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"19120c",x"19130c",x"19130c",x"19120b",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1c09",x"2e1d0a",x"301f0a",x"2f1d0a",x"2b1b09",x"1f1408",x"170f07",x"170f07",x"180f08",x"1a1008",x"1d1208",x"201409",x"23150a",x"24170b",x"24180b",x"26180b",x"27170b",x"26160a",x"26160a",x"25160a",x"231509",x"24150a",x"24150a",x"24150a",x"24150a",x"24150a",x"25160a",x"25160a",x"25160a",x"24150a",x"24150a",x"24150a",x"25150a",x"27160a",x"29180b",x"29180b",x"28170a",x"28170a",x"29170b",x"2a190b",x"28170b",x"26160a",x"2a180b",x"2a190b",x"29170b",x"2a190b",x"29170b",x"27160a",x"27160a",x"251509",x"251509",x"261609",x"261609",x"26160a",x"28170a",x"27170a",x"26160a",x"241509",x"231509",x"201309",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1e1208",x"1f1208",x"201309",x"201309",x"201309",x"201309",x"201208",x"1e1208",x"1d1208",x"1c1108",x"1c1108",x"191007",x"191007",x"160e07",x"150e07",x"150e07",x"150e07",x"32200a",x"231608",x"1f1308",x"1f1308",x"170f07",x"181007",x"180f07",x"150e07",x"472912",x"452811",x"442510",x"3e220f",x"2a190c",x"150e07",x"472a14",x"4a2d16",x"201409",x"1e1209",x"191008",x"301e0a",x"311f0a",x"34210b",x"33200a",x"33200a",x"311f0a",x"190f08",x"150e07",x"231409",x"321d0b",x"4a2a13",x"4b2c14",x"492a13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594b3b",x"574a3a",x"594b3b",x"574537",x"5b4b3b",x"5e4d3e",x"5b4d3d",x"5e4f3f",x"5e4e3f",x"5f503f",x"5d503f",x"665242",x"675241",x"655141",x"655140",x"604f3f",x"5d4d3d",x"5f503f",x"5c4d3e",x"554939",x"5a4c3b",x"584a3a",x"514436",x"544738",x"534537",x"554738",x"4b4032",x"4b3d31",x"4f4033",x"4f4133",x"46382d",x"4b3f32",x"4d3f32",x"524436",x"4b3d31",x"614f40",x"604f40",x"574839",x"5e4e3e",x"675242",x"645342",x"615141",x"645443",x"625443",x"605141",x"645645",x"615444",x"5d5141",x"5f5242",x"5f5242",x"605141",x"615343",x"554839",x"5d5041",x"615141",x"625040",x"655142",x"635343",x"615141",x"645242",x"625141",x"5c4e3e",x"5a4c3b",x"5b4c3c",x"5e4d3d",x"634e3e",x"5d4b3c",x"5a4c3c",x"5c4e3e",x"4c4033",x"5b4a3b",x"544436",x"5e4b3b",x"574838",x"584939",x"5e4a3b",x"564738",x"514336",x"584738",x"4d3e31",x"4a3e2f",x"4c3e31",x"554737",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"1a130c",x"1f1812",x"221b15",x"211a15",x"221c15",x"211b14",x"201913",x"1c160f",x"19120b",x"150e07",x"160e07",x"180f07",x"1d1108",x"231509",x"28170a",x"2b190b",x"2f1b0d",x"301c0d",x"311c0d",x"331d0e",x"331d0d",x"361f0e",x"39210f",x"38200e",x"3b220f",x"3e2511",x"412612",x"412512",x"3e2310",x"3e2410",x"3e2410",x"3d2310",x"3e2410",x"3e2411",x"3c2210",x"38200e",x"37200e",x"361f0e",x"301c0d",x"2d190b",x"28170a",x"231409",x"211409",x"1c1108",x"1c1108",x"1c1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19130c",x"19130c",x"1a130c",x"1a130c",x"19130c",x"1a130c",x"171009",x"17100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"35200c",x"311e0b",x"2c1c09",x"271909",x"211508",x"1d1208",x"150e07",x"160f07",x"170f07",x"191008",x"1b1108",x"1e1309",x"21150a",x"24150a",x"25160a",x"26170b",x"25160a",x"25160a",x"231509",x"23150a",x"23150a",x"231509",x"221509",x"23150a",x"231509",x"24160a",x"24150a",x"25150a",x"26160a",x"27170b",x"28170b",x"26160a",x"27170a",x"27170a",x"28170a",x"29180b",x"2a190b",x"29180b",x"28170b",x"28170b",x"29180b",x"28170a",x"28170b",x"28170a",x"26160a",x"28170b",x"29180b",x"28170b",x"29170b",x"2a190b",x"29180b",x"2a190b",x"2a190b",x"2a180b",x"29180b",x"27160a",x"27160a",x"25150a",x"231509",x"1f1309",x"1e1208",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1f1309",x"1f1309",x"1f1209",x"1f1309",x"201309",x"211409",x"201308",x"201409",x"1b1108",x"1a1008",x"1c1107",x"191007",x"160e07",x"150e07",x"150e07",x"201309",x"37220b",x"32200a",x"211508",x"251708",x"181007",x"170f07",x"1b1108",x"563219",x"583318",x"472813",x"432511",x"3b2210",x"311d0f",x"20140b",x"482812",x"4d2c15",x"1f1309",x"1b1108",x"170f07",x"150e07",x"32200a",x"33200a",x"33200a",x"311f0a",x"301e0a",x"331c0c",x"17110a",x"2e1a0c",x"3a210f",x"422511",x"492a13",x"4f2f16",x"533118",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383431",x"353332",x"353331",x"373332",x"363332",x"363332",x"343231",x"363534",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343332",x"343332",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"584b3b",x"514435",x"4e4133",x"4e4133",x"4e4133",x"4a3e31",x"554939",x"584b3b",x"574a3b",x"564939",x"564939",x"574a3a",x"564939",x"584b3b",x"5e4e3e",x"594b3b",x"574a3a",x"594b3b",x"574537",x"5b4b3b",x"5e4d3e",x"5b4d3d",x"5e4f3f",x"5e4e3f",x"5f503f",x"5d503f",x"665242",x"675241",x"655141",x"655140",x"604f3f",x"5d4d3d",x"5f503f",x"5c4d3e",x"554939",x"5a4c3b",x"584a3a",x"544738",x"544738",x"534537",x"554738",x"524537",x"4b3d31",x"4f4033",x"4f4133",x"544436",x"5e5141",x"615443",x"635241",x"5d4d3e",x"615040",x"5f5040",x"5e5140",x"605140",x"5e5140",x"645141",x"625040",x"615040",x"625141",x"5b4e3e",x"5e5140",x"5d5140",x"5d4f3f",x"5d5140",x"635141",x"655242",x"665242",x"655141",x"5c4f3f",x"5b4d3e",x"614e3e",x"685444",x"5c4d3d",x"584a3b",x"5e4d3e",x"5d4c3c",x"19130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"18110b",x"1f1812",x"221b15",x"211a15",x"221c15",x"211b14",x"201913",x"1c160f",x"19120b",x"150e07",x"160e07",x"180f07",x"1d1108",x"231509",x"28170a",x"2e1b0c",x"2a180b",x"2b180b",x"311d0d",x"331e0e",x"331e0e",x"341e0d",x"331c0d",x"371f0e",x"3a210f",x"3b220f",x"3c2210",x"3f2411",x"3e2411",x"3e2310",x"402511",x"3d2310",x"3b220f",x"381f0e",x"381f0e",x"38200e",x"351e0d",x"321c0c",x"2e1a0b",x"2a180b",x"26160a",x"221409",x"1e1208",x"1e1208",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120c",x"19120c",x"19120c",x"19130c",x"19130c",x"17110a",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2d15",x"4f2f15",x"432811",x"3e260f",x"3b220e",x"361f0d",x"331e0d",x"37200e",x"321d0d",x"36210f",x"331d0d",x"2e1b0d",x"38210f",x"351f0e",x"372110",x"351f0f",x"341e0e",x"341f0f",x"36200f",x"392210",x"331d0d",x"321c0d",x"321d0d",x"36200f",x"3a2210",x"331d0d",x"331d0d",x"301b0c",x"351e0d",x"331d0d",x"351e0e",x"331e0e",x"341e0e",x"331d0d",x"39210f",x"341e0e",x"351e0d",x"321d0d",x"311b0c",x"351e0e",x"331d0d",x"331d0d",x"311b0c",x"311b0c",x"311b0c",x"311b0c",x"331c0c",x"2d1a0b",x"361f0e",x"341e0d",x"361e0e",x"331d0d",x"311b0c",x"331d0d",x"321c0d",x"331d0d",x"321c0d",x"361f0e",x"331d0d",x"341d0d",x"361f0e",x"331c0d",x"331c0c",x"331c0c",x"361e0d",x"321c0d",x"2c180a",x"2b180a",x"301a0b",x"2e190b",x"321b0c",x"321c0c",x"341d0c",x"371e0c",x"341d0c",x"321b0c",x"321c0c",x"341d0c",x"2f1a0b",x"2c180b",x"301a0b",x"43230e",x"33200a",x"34200a",x"3b250c",x"251709",x"1c1208",x"1b1208",x"1b1108",x"4e2d16",x"563218",x"502f16",x"4b2b15",x"462914",x"3e2514",x"24170d",x"4f2d15",x"4d2c15",x"3f2410",x"170f07",x"150e07",x"150e07",x"311f0a",x"321f0a",x"34200a",x"33200a",x"2e1d0a",x"351d0e",x"1d130a",x"331e0f",x"392110",x"3c2310",x"4d2c14",x"533118",x"512e15",x"512d14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"33312f",x"33312f",x"363331",x"383431",x"353332",x"353331",x"373332",x"363332",x"363332",x"343231",x"363534",x"3b3632",x"3a3532",x"353231",x"2f2d2b",x"2f2f2f",x"333333",x"323232",x"333333",x"323232",x"333333",x"313131",x"323131",x"2d2d2d",x"333333",x"333333",x"323232",x"333333",x"333333",x"2b2c2c",x"303030",x"313030",x"343332",x"343332",x"353331",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"584b3b",x"514435",x"4e4133",x"4e4133",x"4e4133",x"4a3e31",x"554939",x"584b3b",x"574a3b",x"564939",x"504334",x"574a3a",x"564939",x"584b3b",x"57493a",x"4d4233",x"4d4234",x"514436",x"56493a",x"5a4a3b",x"5b4c3d",x"5a4b3d",x"5e4e3f",x"604e3e",x"644f3f",x"645141",x"665141",x"594d3d",x"5b4d3e",x"5c4e3e",x"604f3f",x"665141",x"604f3f",x"5d4c3d",x"5a4b3c",x"61503f",x"5f5040",x"615040",x"604e3e",x"574b3b",x"5b4c3c",x"5b4b3b",x"5e4d3d",x"5f503f",x"634f3f",x"604e3e",x"584b3c",x"594d3c",x"5d503f",x"625140",x"5f5140",x"624f3f",x"61503f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"19120b",x"19120c",x"19130c",x"171009",x"160f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"26160a",x"26160a",x"26160a",x"2a180b",x"2a180b",x"301c0d",x"301c0c",x"311c0c",x"321c0c",x"361f0e",x"39200f",x"3b220f",x"3f2511",x"3e2411",x"3e2411",x"3f2511",x"3f2411",x"3e2410",x"3d2310",x"3c2310",x"3b2210",x"39210f",x"351e0d",x"311c0c",x"2c190b",x"27160a",x"241509",x"201309",x"1c1108",x"201309",x"231509",x"2c190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130c",x"1a130c",x"19120c",x"1a130c",x"19130c",x"17110a",x"171009",x"17100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"533116",x"512e15",x"4a2b11",x"4b2d11",x"4c2c13",x"4a2a13",x"482913",x"4a2b14",x"4c2b15",x"452712",x"492913",x"462813",x"462712",x"462813",x"4a2c15",x"482a14",x"482a14",x"472913",x"472913",x"4a2b14",x"4a2a14",x"412410",x"432612",x"4d2e16",x"4b2c15",x"452712",x"412410",x"442711",x"472812",x"462812",x"462914",x"462813",x"452712",x"452813",x"452813",x"432712",x"422611",x"422711",x"452813",x"452813",x"432611",x"402411",x"412410",x"3c220f",x"3c210f",x"412510",x"412510",x"412510",x"422410",x"3f230f",x"412410",x"3e220f",x"3a1f0d",x"3b200e",x"391f0d",x"3d210e",x"3d210f",x"3f220f",x"432511",x"452711",x"4b2b13",x"492a13",x"4c2c14",x"4b2b14",x"4c2c14",x"442611",x"4c2c14",x"442611",x"422410",x"462712",x"482913",x"4f2e16",x"502e15",x"512f16",x"512f17",x"512f16",x"4c2b13",x"482811",x"44240f",x"4c2b13",x"502e16",x"43230e",x"301e0a",x"2f1e0a",x"2c1c09",x"1c1208",x"1d1308",x"1c1208",x"170f07",x"241609",x"4f2e16",x"4a2812",x"502d15",x"512e15",x"4d2d15",x"301c0c",x"502d15",x"512e16",x"2a180b",x"351e0e",x"422510",x"150e07",x"251709",x"291909",x"301e0a",x"2e1d0a",x"2c1c09",x"452911",x"1a1007",x"3d220e",x"41230e",x"3f200d",x"4b2913",x"492710",x"512d14",x"492812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"33302e",x"33302e",x"363331",x"383330",x"343231",x"373533",x"34312f",x"363332",x"353230",x"363433",x"363432",x"393533",x"3a3532",x"353231",x"2f2d2b",x"333333",x"333333",x"323232",x"333333",x"323232",x"323232",x"313131",x"323131",x"2d2d2d",x"333333",x"333333",x"323232",x"323232",x"333333",x"2b2c2c",x"303030",x"313030",x"343332",x"363332",x"353230",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"463a2d",x"463a2d",x"463a2d",x"493b2f",x"4f4134",x"4a3c30",x"4c3f32",x"4d4134",x"4e4235",x"44392d",x"493d31",x"534637",x"4b4033",x"4d4134",x"514537",x"514537",x"514536",x"504335",x"504336",x"554738",x"594739",x"5c4c3d",x"584b3c",x"5d4d3f",x"604d3d",x"605141",x"56493a",x"584b3c",x"5b4e3e",x"605242",x"5c4d3d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"19120b",x"19120c",x"19130c",x"171009",x"160f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"271a0b",x"26190b",x"22170b",x"1c130a",x"20160b",x"24190d",x"22180d",x"20160d",x"1d140c",x"19120c",x"19120b",x"1b130c",x"1c140b",x"1d150c",x"1a140c",x"1d140c",x"1f150c",x"25190c",x"24190d",x"24180d",x"25190d",x"22160a",x"2b1c0b",x"25190b",x"24180a",x"1f150b",x"191109",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"19130c",x"1a130c",x"19130c",x"17110b",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211409",x"211409",x"23150a",x"25160a",x"28170b",x"2d1a0c",x"2f1c0d",x"321d0d",x"331d0d",x"361f0e",x"3a210f",x"3b220f",x"3f2511",x"3d2310",x"3c220f",x"3a210f",x"3b220f",x"3a2210",x"3c2311",x"39210f",x"37200f",x"361f0e",x"351f0e",x"321c0c",x"29170a",x"29170a",x"241409",x"211308",x"341c0c",x"2e190b",x"2e190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120b",x"19120b",x"19120b",x"19130c",x"19120c",x"17110a",x"171009",x"18110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"563318",x"563318",x"5d381a",x"5a3719",x"573419",x"502f16",x"512f16",x"4d2c15",x"492913",x"4e2d15",x"502e16",x"4a2a13",x"4b2a13",x"462711",x"492912",x"4c2b14",x"4c2c15",x"492a13",x"4a2a14",x"4e2d15",x"4c2c14",x"4c2b14",x"4e2d14",x"4a2a13",x"492b14",x"4c2c14",x"4b2b14",x"472812",x"472812",x"4a2b14",x"482913",x"4d2d16",x"4a2b14",x"492a14",x"432711",x"442712",x"432611",x"462914",x"472913",x"482a14",x"482a13",x"452812",x"452812",x"412411",x"3c210e",x"3d210e",x"341c0c",x"3d200e",x"3b1f0d",x"3d210e",x"452812",x"462812",x"412511",x"432610",x"442711",x"432611",x"3e230f",x"3f220f",x"3d220e",x"432510",x"462711",x"482812",x"472913",x"482913",x"472913",x"452711",x"42240f",x"3f230f",x"432510",x"412510",x"472812",x"432410",x"422510",x"4c2b13",x"4a2b12",x"472610",x"4e2e14",x"4e2d15",x"472811",x"4f2d14",x"4a2812",x"42230e",x"503113",x"44280f",x"472a11",x"3f260e",x"1b1108",x"472914",x"38200e",x"2e1a0b",x"402511",x"432611",x"3f2310",x"422511",x"412612",x"211309",x"341e0f",x"2c1a0e",x"371f0f",x"3c2110",x"432511",x"301c0b",x"3e250f",x"492c13",x"513115",x"533316",x"533217",x"4e2c14",x"2f1a0b",x"492911",x"43240f",x"43230e",x"4e2b13",x"44250f",x"512e14",x"512e14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"33312f",x"33312f",x"393330",x"32302f",x"353332",x"373331",x"373433",x"363230",x"383432",x"332e2b",x"383331",x"363230",x"3d3733",x"343231",x"363331",x"313131",x"343434",x"333333",x"313131",x"303030",x"323232",x"323232",x"323232",x"313131",x"313131",x"323232",x"323232",x"313131",x"343434",x"303131",x"323232",x"313030",x"333231",x"353231",x"373331",x"535151",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"493b2f",x"493b2f",x"504234",x"514335",x"524335",x"5a493a",x"634d3d",x"5d483a",x"171009",x"171009",x"514636",x"241c13",x"271f16",x"261d15",x"261e16",x"271f16",x"150e07",x"150e07",x"2a2118",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"9e9e9e",x"150e07",x"150e07",x"150e07",x"171009",x"1a130c",x"1a130c",x"19130c",x"171009",x"17110a",x"17110a",x"1b140d",x"20170f",x"271b0e",x"20160d",x"1c130a",x"1c1108",x"1d140b",x"20170d",x"22170e",x"251a0e",x"1c150e",x"1e170f",x"1e160f",x"201810",x"221910",x"231a10",x"1f170f",x"221911",x"231910",x"261b0f",x"291c10",x"23190f",x"21170c",x"1e150b",x"1e150d",x"1c130c",x"1d130b",x"1a110a",x"180f07",x"191007",x"1d1308",x"1d1308",x"1f1408",x"221508",x"231608",x"1d1308",x"221508",x"231608",x"251809",x"271a0b",x"26190b",x"22170b",x"1c130a",x"20160b",x"24190d",x"22180d",x"20160d",x"1d140c",x"19120c",x"19120b",x"1b130c",x"1c140b",x"1d150c",x"1a140c",x"1d140c",x"1f150c",x"25190c",x"24190d",x"24180d",x"25190d",x"22160a",x"2b1c0b",x"25190b",x"24180a",x"1f150b",x"191109",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"19130c",x"1a130c",x"19130c",x"17110b",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"1d1108",x"311c0c",x"311b0c",x"2d190b",x"2d190b",x"29170a",x"2c190b",x"2f1a0c",x"27160a",x"29160a",x"321c0c",x"2d190b",x"2d190b",x"321c0c",x"2e190b",x"2c180b",x"321c0c",x"2d1a0b",x"2d190b",x"2f1a0b",x"321c0c",x"2d190b",x"321c0c",x"1c1108",x"1c1108",x"29170a",x"321c0d",x"361f0e",x"3a210f",x"3c220f",x"402410",x"3a200e",x"3c210e",x"3e220f",x"402310",x"432510",x"402410",x"422410",x"402310",x"3f230f",x"412410",x"412510",x"442510",x"3c210e",x"422511",x"432511",x"442712",x"432611",x"472813",x"3c220f",x"3f2410",x"472813",x"402510",x"402510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120c",x"19120c",x"1a130c",x"19120b",x"19120c",x"17110a",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"553216",x"593316",x"543114",x"4d2d12",x"4b2a12",x"4b2a12",x"482912",x"472812",x"422510",x"462811",x"472812",x"432611",x"472912",x"4a2a14",x"472913",x"482a13",x"422511",x"442611",x"422410",x"422511",x"3d210e",x"452812",x"472913",x"452712",x"432611",x"422511",x"422511",x"3b200e",x"3b210e",x"3c220f",x"3a200e",x"3b220f",x"412511",x"3f2411",x"3f2411",x"412511",x"3d230f",x"3e2310",x"3c220f",x"3d2310",x"3f2410",x"3f2310",x"3f2410",x"3d2310",x"3f2410",x"422511",x"482a13",x"3f2410",x"3f2410",x"412510",x"3b200e",x"40240f",x"371f0d",x"3b200e",x"3b210e",x"3d220f",x"3c220f",x"3a210f",x"3b220f",x"351e0d",x"3c230f",x"3b210f",x"38200e",x"442712",x"432612",x"422611",x"432611",x"3f2410",x"3b210f",x"3c210f",x"3d220e",x"41230f",x"40230f",x"452610",x"462710",x"452711",x"4a2b12",x"4c2b14",x"4c2c14",x"462711",x"4e2e14",x"583415",x"513012",x"633d16",x"452810",x"2a170a",x"4a2913",x"3f230f",x"2a180c",x"18100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"24160c",x"24170d",x"291a0e",x"26180d",x"422714",x"2e1d0f",x"382210",x"442911",x"492c13",x"4a2c11",x"5c3618",x"1b1108",x"1b1108",x"191007",x"160e07",x"150e07",x"150e07",x"170f07",x"3e2310",x"40230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"474645",x"454242",x"393635",x"343231",x"363433",x"393532",x"35312f",x"363332",x"363331",x"363331",x"34302e",x"3a3431",x"383431",x"3c3531",x"383432",x"363432",x"333232",x"343333",x"333333",x"323232",x"313131",x"313131",x"313131",x"333333",x"313131",x"333333",x"323232",x"313131",x"323232",x"313131",x"313131",x"313131",x"454545",x"4c4b4b",x"4d4b4a",x"434342",x"434342",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"473a2e",x"473a2e",x"352b21",x"4d4135",x"504134",x"2f251c",x"4f3d30",x"5d483a",x"221912",x"291f17",x"4a3f31",x"241c13",x"271f16",x"261d15",x"150e07",x"271f16",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"17110a",x"1a130c",x"19120b",x"19130c",x"171009",x"171009",x"171009",x"19130c",x"21170e",x"261a0d",x"21170d",x"1b1108",x"180f07",x"1d130b",x"1d130b",x"1d150c",x"20160e",x"1d1710",x"1f1810",x"1f160f",x"231a11",x"201810",x"1f170f",x"1e160f",x"20170e",x"20170e",x"22180e",x"281b0e",x"1d150c",x"1d140c",x"1c140c",x"1c130b",x"191109",x"1d130a",x"1a110a",x"180f07",x"191007",x"1d1308",x"1e1308",x"1f1408",x"211508",x"211508",x"1a1107",x"1d1208",x"211508",x"251709",x"281a09",x"26190b",x"20150b",x"18110a",x"1c1309",x"20160a",x"20150a",x"1e140a",x"1b1209",x"171009",x"171009",x"171009",x"191109",x"1b1209",x"18110a",x"1a1109",x"1c130c",x"271a0d",x"24180a",x"20160b",x"23170b",x"20160a",x"2d1d0b",x"271a0c",x"23180a",x"1e140b",x"191109",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"17110a",x"19120b",x"19130c",x"19120b",x"17100a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"717070",x"2f1a0b",x"311c0c",x"311b0c",x"2d190b",x"2d190b",x"29170a",x"2c190b",x"2f1a0c",x"27160a",x"29160a",x"321c0c",x"2d190b",x"2d190b",x"321c0c",x"2e190b",x"2c180b",x"321c0c",x"2d1a0b",x"2d190b",x"2f1a0b",x"321c0c",x"2d190b",x"321c0c",x"311c0c",x"321c0d",x"311c0d",x"2d190b",x"2b180b",x"2d190b",x"2e1a0b",x"2c190b",x"2d1a0b",x"231409",x"27160a",x"241509",x"26160a",x"28170a",x"26160a",x"26160a",x"211409",x"211409",x"221409",x"1e1208",x"1d1108",x"191008",x"1e1209",x"1d1108",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"402510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120b",x"19120b",x"19120c",x"19120b",x"1a130c",x"17100a",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"5a3618",x"533115",x"5e391a",x"5b3719",x"563417",x"513016",x"492b15",x"4e2e17",x"492b16",x"462a15",x"462a14",x"482b16",x"462915",x"442812",x"402512",x"452814",x"422713",x"432713",x"3e2410",x"402513",x"412613",x"3e2412",x"3f2311",x"3d2211",x"402511",x"432814",x"412612",x"3b2211",x"371f10",x"3a2110",x"3c2211",x"351d0e",x"321d0d",x"341d0e",x"371e0f",x"311c0d",x"321c0d",x"331d0e",x"321c0e",x"341d0e",x"301a0d",x"361e0f",x"321d0d",x"301a0c",x"27160b",x"2d190c",x"351e0e",x"38200f",x"3b2211",x"3c2211",x"331d0d",x"301a0c",x"311b0d",x"301b0d",x"2a170b",x"361f0f",x"392110",x"311b0d",x"311c0d",x"321c0e",x"351e0f",x"392110",x"3a2110",x"392110",x"3c2210",x"3c2110",x"3f2411",x"3c2211",x"3d2211",x"351e0f",x"422713",x"432611",x"432813",x"482b15",x"4b2c15",x"4d2e15",x"503017",x"523217",x"553218",x"462510",x"593517",x"593616",x"543415",x"4e3015",x"422913",x"3b2511",x"4a2c18",x"3f2615",x"19120b",x"19120c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"23150a",x"23150a",x"2e1b0d",x"2e1b0e",x"3e2512",x"281a0d",x"392311",x"442b15",x"492e16",x"5a3619",x"5f3a1b",x"160e07",x"180f07",x"191007",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"301b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4847",x"4a4847",x"4c4b49",x"474442",x"474442",x"4d4b4a",x"4e4c4a",x"545251",x"575555",x"54514f",x"595755",x"5d5a57",x"605d5c",x"3d3835",x"373432",x"353331",x"323131",x"323232",x"3b3b3b",x"4d4d4d",x"60605f",x"515151",x"2f2f2f",x"333333",x"2b2b2b",x"313131",x"343434",x"313131",x"333333",x"323232",x"3b3b3b",x"484543",x"4e4e4d",x"504c4b",x"545252",x"4a4847",x"4a4847",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"473a2e",x"352b21",x"4d4135",x"504134",x"2f251c",x"4f3d30",x"5d483a",x"221912",x"291f17",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"17110a",x"171009",x"150e07",x"150e07",x"17110a",x"19130c",x"1f160d",x"24180d",x"1d1308",x"1b1108",x"170f07",x"1a1107",x"1c130a",x"1d140c",x"1e160c",x"1b140d",x"1b150e",x"1b150e",x"1e160d",x"1e160e",x"1d160d",x"1c150f",x"1d150c",x"1d150c",x"20170d",x"271a0b",x"1a1209",x"1a110a",x"19110a",x"19110a",x"170f07",x"1b1108",x"170f07",x"170f07",x"191007",x"1c1208",x"1d1208",x"1f1408",x"201508",x"1f1408",x"181007",x"1c1208",x"1f1408",x"231608",x"211508",x"231608",x"1c1208",x"150e07",x"150e07",x"20150a",x"1f140a",x"1d130a",x"1b1209",x"171009",x"171009",x"171009",x"171009",x"181109",x"171009",x"181009",x"181109",x"191109",x"24180b",x"20150a",x"281b0b",x"23180a",x"25190b",x"26190b",x"231608",x"1c1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"17100a",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"201308",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"160f07",x"180f07",x"160f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130c",x"1a130c",x"19130c",x"1a130c",x"1a130c",x"171009",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"533115",x"543316",x"4e3017",x"583517",x"553318",x"523117",x"4b2d17",x"482c17",x"462a16",x"482c17",x"492c17",x"422815",x"3b2312",x"3f2513",x"3e2513",x"422815",x"3d2312",x"3a2313",x"3b2211",x"3d2412",x"3f2614",x"3d2413",x"3c2212",x"3e2513",x"3d2412",x"3b2312",x"382111",x"3a2212",x"382111",x"341f10",x"382011",x"382111",x"372111",x"392212",x"372111",x"372211",x"372011",x"382111",x"382111",x"382011",x"351d0e",x"331d0e",x"351e0f",x"39200f",x"331d0e",x"361e0f",x"2d1a0d",x"2c1a0c",x"321d0e",x"361e0f",x"341d0e",x"2f1b0d",x"2f1b0c",x"2c180c",x"29170c",x"24130a",x"27170b",x"2e1b0d",x"321c0e",x"301c0e",x"301c0d",x"321c0e",x"351e0e",x"341d0e",x"372010",x"361e0f",x"3b2211",x"3c2211",x"392010",x"381f0f",x"361e0f",x"392010",x"3c2210",x"3c2210",x"3d2310",x"432611",x"432812",x"4d2c15",x"4d2c15",x"4c2b14",x"593616",x"553215",x"563417",x"482b13",x"412711",x"28190b",x"472a14",x"402511",x"17100a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"211409",x"2b190b",x"37200e",x"341e0d",x"1a1107",x"36210d",x"40260f",x"533216",x"593619",x"5b3619",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4847",x"4c4b49",x"474442",x"474442",x"4d4b4a",x"4e4c4a",x"545251",x"575555",x"54514f",x"595755",x"5d5a57",x"605d5c",x"3d3835",x"373432",x"353331",x"323131",x"313131",x"3b3b3b",x"4d4d4d",x"60605f",x"515151",x"494949",x"464646",x"535353",x"3b3b3b",x"3e3e3e",x"454545",x"414141",x"424242",x"4e4e4e",x"535353",x"515151",x"545353",x"545252",x"4a4847",x"4a4847",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"1e160d",x"21170b",x"1d1208",x"1a1107",x"160f07",x"1b1108",x"1d130b",x"1c130a",x"1c140b",x"1a130c",x"1a130c",x"19120c",x"1c140b",x"1b130c",x"1b130c",x"19120b",x"1c1309",x"1c130a",x"1f140b",x"261a0b",x"181007",x"170f07",x"160f07",x"180f07",x"160f07",x"1b1108",x"180f07",x"170f07",x"191007",x"1d1208",x"1d1308",x"1e1308",x"201408",x"1e1308",x"180f07",x"1b1108",x"1e1308",x"211508",x"1f1408",x"211508",x"1a1107",x"150e07",x"150e07",x"1d1208",x"1c1208",x"1a1107",x"181007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211508",x"211508",x"201408",x"201508",x"221608",x"241708",x"221508",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160f07",x"170f07",x"160f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19130c",x"19130c",x"19120c",x"19120b",x"19120b",x"17110a",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"4e3017",x"4f3115",x"4b2d13",x"563416",x"4f2f13",x"4c2d15",x"3f2410",x"3f2410",x"402410",x"3e220f",x"3c210f",x"3a220f",x"3e2310",x"3a210f",x"3f2410",x"3e2410",x"3c2210",x"3e2411",x"3f2512",x"402511",x"3e2310",x"402410",x"3b220f",x"3b210f",x"39210f",x"3a210f",x"381f0e",x"381f0d",x"371f0d",x"3a210f",x"3d220f",x"38200e",x"3a210f",x"3b210f",x"3a210f",x"341d0d",x"311b0b",x"2f190b",x"301b0b",x"361d0d",x"361e0d",x"351d0d",x"341d0c",x"321c0c",x"311a0b",x"2b170a",x"2e180a",x"321c0c",x"361e0d",x"351d0c",x"2f1a0b",x"351e0d",x"351d0d",x"331c0c",x"331c0c",x"331c0c",x"311b0c",x"371f0d",x"331c0d",x"3a210f",x"3e2310",x"3b210f",x"351e0d",x"38200e",x"3e2411",x"3d2310",x"3d2310",x"3b2210",x"38200f",x"3b2310",x"392110",x"3b2210",x"3d2411",x"432712",x"432812",x"462912",x"41240f",x"4b2b14",x"4d2c15",x"000000",x"563417",x"533215",x"583516",x"37200e",x"2a190a",x"3c210e",x"512c14",x"442610",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"201309",x"2f1b0c",x"24150a",x"3a200f",x"211509",x"34200c",x"563316",x"583416",x"533216",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d322a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494949",x"464646",x"535353",x"505050",x"3e3e3e",x"454545",x"414141",x"4e4e4e",x"4e4e4e",x"515151",x"545454",x"545353",x"433932",x"3f3329",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f4e4d",x"4a4948",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"514e4e",x"514e4e",x"3f3d3c",x"343231",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"1f1408",x"1c1208",x"1a1107",x"160f07",x"191007",x"191007",x"181007",x"191007",x"150e07",x"150e07",x"150e07",x"181007",x"170f07",x"170f07",x"150e07",x"181007",x"1a1107",x"1c1208",x"241708",x"181007",x"170f07",x"160f07",x"170f07",x"170f07",x"1a1107",x"170f07",x"170f07",x"191007",x"1c1208",x"1c1208",x"1d1308",x"1f1408",x"1d1308",x"170f07",x"1a1108",x"1d1208",x"201408",x"1d1308",x"201408",x"191007",x"150e07",x"150e07",x"1c1208",x"1b1108",x"191007",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"1c1208",x"1b1208",x"1d1208",x"211508",x"231608",x"201508",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"190f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160f07",x"170f07",x"160f07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120c",x"19120c",x"1a130c",x"19120b",x"19120b",x"17110a",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"452910",x"42270f",x"513015",x"4d2d14",x"492b13",x"432510",x"472913",x"402411",x"3c210f",x"402511",x"432612",x"452813",x"402410",x"432712",x"412511",x"3c2210",x"3c2310",x"412511",x"412612",x"452813",x"3e2411",x"3d2310",x"3c2210",x"3f2511",x"3e2411",x"3a2210",x"3e2411",x"3e2411",x"371f0e",x"3a200e",x"371f0d",x"341d0d",x"38200e",x"3a220f",x"3b2210",x"3b220f",x"3b220f",x"3f2411",x"3d2310",x"3a210f",x"3b210f",x"361e0d",x"3c220f",x"3c220f",x"3a210f",x"3c2310",x"381f0e",x"3f2511",x"3a210f",x"3a210f",x"3a2210",x"3c220f",x"3a210f",x"402511",x"3b220f",x"3a210f",x"3b210f",x"381f0d",x"3c220f",x"3f2411",x"3f2410",x"3d2210",x"412511",x"472a15",x"462914",x"442813",x"3f2511",x"412612",x"402612",x"3a210f",x"39200f",x"3f2310",x"412612",x"472a14",x"3d210e",x"41240f",x"41240f",x"000000",x"000000",x"000000",x"4b2b10",x"4b2a11",x"3d240f",x"201309",x"2f1a0b",x"29170a",x"251509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1208",x"1e1208",x"29170a",x"241409",x"301a0b",x"201309",x"442810",x"4e2e14",x"563316",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"40352c",x"3d322a",x"3d322a",x"3a2f27",x"3f362f",x"423830",x"3e3631",x"413831",x"403832",x"3f3832",x"3f3631",x"413933",x"433931",x"403832",x"3f3630",x"403833",x"3d3632",x"3e3632",x"3e3630",x"3d2f26",x"3f3731",x"413832",x"423831",x"3f3630",x"433932",x"443932",x"433931",x"3f352e",x"3f3630",x"423831",x"433831",x"453a31",x"433932",x"3f3329",x"3f3329",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f4e4d",x"4f4e4d",x"4a4948",x"353332",x"2f2116",x"323131",x"000000",x"000000",x"000000",x"515050",x"514e4e",x"353332",x"353433",x"353434",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"1d1308",x"1b1108",x"191007",x"160f07",x"191007",x"191107",x"181007",x"191007",x"150e07",x"150e07",x"150e07",x"181007",x"170f07",x"170f07",x"150e07",x"191007",x"191007",x"1b1108",x"231608",x"181007",x"170f07",x"160f07",x"170f07",x"160f07",x"1a1107",x"170f07",x"170f07",x"181007",x"1b1108",x"1c1208",x"1c1208",x"1d1308",x"1c1208",x"170f07",x"1a1107",x"1c1208",x"1d1308",x"1c1208",x"1e1308",x"181007",x"150e07",x"150e07",x"1a1107",x"1a1107",x"191007",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"1b1108",x"1b1108",x"1c1208",x"1f1408",x"211508",x"1f1408",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"160e07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19120b",x"19120b",x"19120b",x"19120b",x"19120b",x"17110a",x"171009",x"17100a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"39230e",x"331e0b",x"4a2a13",x"422610",x"3c210f",x"402411",x"412511",x"3b210f",x"3d220f",x"3c210f",x"3a200e",x"3d220f",x"3b210f",x"39200e",x"3a200e",x"3a210f",x"381f0d",x"361e0d",x"3b210e",x"391f0e",x"351d0c",x"361e0d",x"331c0c",x"3a210f",x"39210f",x"38200e",x"39200e",x"381f0e",x"38210f",x"3a200f",x"39210f",x"38200e",x"361e0e",x"361e0d",x"3a200e",x"381f0e",x"3a200e",x"351d0d",x"341d0c",x"341d0c",x"361e0d",x"39200e",x"38200e",x"3b210f",x"391f0e",x"39200e",x"39200e",x"39200e",x"3a200f",x"3a210f",x"3e2410",x"3c2310",x"3f2511",x"37200e",x"3c210f",x"361e0d",x"371e0d",x"351d0d",x"391f0d",x"361e0d",x"371e0d",x"3d220f",x"412411",x"38200e",x"37200f",x"37200f",x"371f0e",x"39210f",x"361f0e",x"37200e",x"3d2310",x"3f2310",x"422511",x"3c200d",x"3d210e",x"000000",x"000000",x"000000",x"000000",x"40220e",x"472810",x"492911",x"24160b",x"3e2310",x"381f0e",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1007",x"1b1008",x"2c170a",x"29160a",x"191008",x"1f1309",x"4b2b14",x"472910",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"44382e",x"40352c",x"3a3029",x"40362e",x"3f362f",x"423830",x"3e3631",x"453a32",x"403832",x"3f3832",x"3f3631",x"413933",x"433931",x"403832",x"3f3630",x"403833",x"3d3632",x"3e3632",x"3e3630",x"3d2f26",x"3f3731",x"413832",x"423831",x"3f3731",x"433932",x"443932",x"413831",x"3f362f",x"3f362f",x"423831",x"433830",x"473b32",x"433a33",x"3f3229",x"473729",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494747",x"494747",x"343332",x"383634",x"323131",x"323131",x"000000",x"000000",x"535252",x"535252",x"414141",x"333232",x"333332",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191007",x"1c1208",x"1a1107",x"181007",x"160e07",x"181007",x"191007",x"180f07",x"181007",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"160f07",x"150e07",x"181007",x"181007",x"1a1107",x"201508",x"170f07",x"160f07",x"160e07",x"170f07",x"160f07",x"1a1107",x"170f07",x"160f07",x"170f07",x"1a1107",x"1b1108",x"1b1108",x"1c1208",x"1a1107",x"170f07",x"191007",x"1a1107",x"1c1208",x"1a1107",x"1c1208",x"170f07",x"150e07",x"150e07",x"191007",x"191007",x"180f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1107",x"1a1107",x"191107",x"1a1107",x"1d1308",x"1f1408",x"1d1308",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"26160a",x"27170a",x"28170a",x"28170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19130c",x"19130c",x"19120c",x"19130c",x"19130c",x"17100a",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331e0b",x"38210c",x"351f0d",x"3c220f",x"3f2511",x"3c220f",x"3c220f",x"3d2310",x"3c220f",x"351e0d",x"3b210f",x"361f0e",x"38200f",x"371f0e",x"3a200e",x"361e0e",x"361e0d",x"351d0d",x"371f0e",x"331d0d",x"351d0d",x"341d0d",x"341c0d",x"361e0e",x"341d0d",x"331c0c",x"231107",x"2d190a",x"2b180b",x"331c0d",x"351d0d",x"331d0d",x"321c0c",x"361e0d",x"361f0e",x"361f0e",x"351e0d",x"351d0d",x"371f0e",x"351f0e",x"38200f",x"37200e",x"3a220f",x"39210f",x"39210f",x"3b2210",x"38200f",x"361f0e",x"371f0e",x"331d0d",x"331d0d",x"351f0e",x"38200f",x"3a220f",x"38200f",x"3c2310",x"3b2210",x"341e0e",x"3b2311",x"36200f",x"3a2210",x"3b2311",x"361f0d",x"331d0d",x"301c0d",x"311c0d",x"331d0e",x"371f0e",x"351d0d",x"311a0b",x"321b0b",x"2f190b",x"2f1a0b",x"3a200e",x"1c150f",x"1c150f",x"1c150e",x"1c150e",x"1c150e",x"1c150e",x"472811",x"361e0e",x"27160a",x"3c220f",x"381f0e",x"150e07",x"150e07",x"150e07",x"1c150d",x"150e07",x"150e07",x"150e07",x"150e07",x"614c3d",x"665344",x"635043",x"58473b",x"39200e",x"482812",x"482812",x"1a130c",x"19120b",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"171009",x"150e08",x"150e07",x"160f07",x"160f07",x"170f07",x"170f07",x"160f07",x"181007",x"150e07",x"160f07",x"191107",x"170f07",x"1b1108",x"181007",x"1a1008",x"180f07",x"191007",x"181007",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"554c47",x"493f37",x"433932",x"443931",x"3f3631",x"3f3631",x"3e3631",x"3d3631",x"463a32",x"403730",x"3c3632",x"403832",x"413933",x"443a33",x"3f3832",x"423831",x"3b342f",x"3a3430",x"3d3632",x"3b3532",x"403832",x"413831",x"433831",x"423831",x"433932",x"40342b",x"453a32",x"413730",x"42372f",x"423933",x"453b33",x"443930",x"443930",x"453a31",x"433a33",x"453a32",x"4f453f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"373737",x"373737",x"353332",x"383533",x"343332",x"343332",x"000000",x"000000",x"585858",x"585858",x"4f4f4f",x"323131",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1107",x"181007",x"170f07",x"160e07",x"170f07",x"170f07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"170f07",x"160f07",x"160f07",x"150e07",x"170f07",x"170f07",x"181007",x"1d1308",x"170f07",x"160f07",x"160e07",x"160f07",x"160e07",x"181007",x"160f07",x"160f07",x"170f07",x"181007",x"191007",x"191007",x"1a1107",x"191007",x"160f07",x"170f07",x"181007",x"191007",x"191007",x"1a1107",x"170f07",x"150e07",x"150e07",x"180f07",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181007",x"181007",x"181007",x"191007",x"1b1108",x"1c1208",x"1b1108",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"231509",x"28170b",x"2a190b",x"2a190b",x"2a190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19130c",x"19130c",x"19120b",x"19130c",x"19130c",x"1a130c",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"482711",x"40230f",x"462611",x"482913",x"4b2b14",x"4e2e16",x"4e2e16",x"4a2a13",x"452712",x"4c2c15",x"4a2b15",x"4e2e16",x"4a2a15",x"4a2b15",x"4e2d16",x"4a2b15",x"492a14",x"472913",x"452712",x"4d2d16",x"4b2c16",x"4c2c15",x"4c2c15",x"4b2b15",x"472914",x"452813",x"4a2b14",x"472813",x"482914",x"472812",x"4a2b15",x"452813",x"432612",x"452712",x"412510",x"442511",x"452612",x"472812",x"442712",x"452712",x"472913",x"4a2b15",x"452712",x"492a14",x"462813",x"452712",x"462712",x"442611",x"432611",x"462712",x"462812",x"422612",x"442712",x"4a2b15",x"4d2d16",x"452813",x"472914",x"482a14",x"4b2c15",x"452611",x"4a2a14",x"4a2913",x"4c2c14",x"462812",x"462813",x"442611",x"442511",x"432511",x"4b2a13",x"4e2c14",x"1c150f",x"1c150f",x"1c150f",x"1c150e",x"1c150e",x"1c150e",x"1c150e",x"1c150e",x"1c160e",x"422d1f",x"5d4a3c",x"544235",x"524338",x"54453a",x"1c150e",x"1c150d",x"1c150e",x"1c150e",x"150e07",x"150e07",x"1b140d",x"1b140d",x"1b140c",x"1a130d",x"1b140c",x"1b140d",x"1c140d",x"1a130c",x"19120b",x"19120b",x"150e07",x"150e07",x"170f07",x"171009",x"171009",x"171009",x"150e08",x"150e07",x"160f07",x"160f07",x"170f07",x"170f07",x"160f07",x"181007",x"150e07",x"160f07",x"191107",x"170f07",x"1b1108",x"181007",x"1a1008",x"180f07",x"191007",x"181007",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"4f4740",x"534b45",x"58504b",x"5e5956",x"544e4a",x"41362f",x"403831",x"3f3833",x"3e3631",x"413832",x"403833",x"3e3631",x"403831",x"3e3732",x"3f3631",x"433932",x"3e3732",x"413730",x"3d3733",x"3b3531",x"3d3733",x"403730",x"443830",x"433831",x"423830",x"433932",x"443a33",x"463b33",x"443a33",x"403730",x"453930",x"433830",x"433931",x"423932",x"564d47",x"58504b",x"58504b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b4a4a",x"4b4a4a",x"302e2d",x"363331",x"333232",x"333232",x"000000",x"000000",x"4e4e4e",x"545454",x"3a3a3a",x"313131",x"2f2f2f",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"160f07",x"160f07",x"150e07",x"160f07",x"160f07",x"160e07",x"160f07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160f07",x"160f07",x"160f07",x"191007",x"160e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160f07",x"160e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"150e07",x"160f07",x"160f07",x"170f07",x"160f07",x"170f07",x"160e07",x"150e07",x"150e07",x"160f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160f07",x"160f07",x"170f07",x"180f07",x"181007",x"180f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"29180b",x"2c190b",x"2c190b",x"2e1b0c",x"2e1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130c",x"1a130c",x"1a130c",x"1a130c",x"19120c",x"19120b",x"17100a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160e07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160e07",x"160f07",x"160e07",x"160e07",x"150e07",x"160f07",x"160f07",x"160e07",x"150e07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"181007",x"170f07",x"181007",x"170f07",x"170f07",x"160f07",x"180f07",x"170f07",x"160f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"564d48",x"564d48",x"524943",x"554f4a",x"5e5955",x"5a5553",x"463f3b",x"3f3832",x"3f362f",x"3f3833",x"3b342f",x"3f3832",x"3e3732",x"413832",x"3e3632",x"413831",x"615e5b",x"544e4a",x"3e3834",x"322b26",x"362d27",x"3a2f26",x"40342c",x"3f3630",x"67615d",x"625c58",x"5e5854",x"5f5854",x"5f5955",x"5d5651",x"544e49",x"57504b",x"534b45",x"473b33",x"59514c",x"584f4a",x"584f4a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d4c4c",x"474545",x"323131",x"353433",x"363433",x"bbbbbb",x"000000",x"000000",x"464646",x"464646",x"333333",x"333333",x"323232",x"343434",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"1d1208",x"22150a",x"24160a",x"24150a",x"24150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a130d",x"1a130d",x"19130c",x"19120b",x"19120b",x"19120b",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160e07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"564d48",x"534b47",x"544f4b",x"57524f",x"595452",x"57514e",x"423b35",x"443e3a",x"453f3a",x"45403c",x"514d4a",x"4a433f",x"47403c",x"4a4440",x"4f4945",x"5e5956",x"544e4b",x"443d39",x"332b26",x"362d27",x"3a2f26",x"40342c",x"3f3630",x"67615d",x"625c58",x"5e5854",x"5f5854",x"5f5955",x"5d5651",x"544e49",x"57504b",x"534b45",x"473b33",x"59514c",x"584f4a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"464545",x"464545",x"353332",x"323131",x"333332",x"343332",x"343332",x"3f3f3f",x"3f3f3f",x"343434",x"323232",x"333333",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"1b1108",x"1f1209",x"221509",x"211409",x"211409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1c150e",x"19130c",x"19130c",x"19130c",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160e07",x"150e07",x"160e07",x"150e07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"4a4949",x"4a4949",x"4e4e4e",x"3d3d3d",x"000000",x"000000",x"59534f",x"595451",x"595451",x"57514e",x"423b35",x"443e3a",x"453f3a",x"45403c",x"514d4a",x"4a433f",x"47403c",x"4a4440",x"4f4945",x"5e5956",x"544e4b",x"443d39",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f4e4e",x"5b5a5a",x"30302f",x"30302f",x"000000",x"000000",x"000000",x"4d4c4c",x"4d4c4c",x"363331",x"343231",x"323131",x"343333",x"343333",x"393939",x"393939",x"303030",x"343434",x"343434",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"4b2c15",x"3e2310",x"3c2310",x"371f0e",x"381f0e",x"2f1a0b",x"2c190b",x"361f0d",x"412919",x"412919",x"3c230f",x"321c0c",x"3a200f",x"341d0d",x"2b180a",x"311b0b",x"332116",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"1b1108",x"201309",x"22150a",x"23150a",x"23150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"19130c",x"19130c",x"19130c",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"150e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"150e07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"343332",x"343332",x"4a4949",x"4a4a4a",x"323233",x"373737",x"3a3a3a",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b4a4a",x"5d5c5c",x"575655",x"4b4a4a",x"585858",x"30302f",x"2c2c2b",x"000000",x"000000",x"000000",x"525151",x"525151",x"363332",x"333231",x"373534",x"373534",x"373534",x"000000",x"424242",x"424242",x"333333",x"2d2d2d",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"4b2c15",x"4b2c15",x"3e2310",x"3c2310",x"371f0e",x"381f0e",x"2f1a0b",x"2c190b",x"361f0d",x"150e07",x"412919",x"3c230f",x"321c0c",x"3a200f",x"341d0d",x"2b180a",x"311b0b",x"332116",x"332116",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b140e",x"1b140e",x"1b140e",x"19130c",x"19130c",x"19120c",x"17100a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"343333",x"343433",x"312f2d",x"333231",x"323232",x"363636",x"3d3d3d",x"343434",x"323232",x"3b3b3b",x"3e3c3c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"444444",x"474746",x"4a4949",x"504f4f",x"5d5d5d",x"424140",x"353433",x"343332",x"313030",x"31302f",x"000000",x"000000",x"545353",x"545353",x"343332",x"353433",x"363433",x"343232",x"343232",x"000000",x"4b4b4b",x"4b4b4b",x"2f2f2f",x"303030",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"311c0d",x"311c0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29160a",x"523b2d",x"594638",x"574437",x"5c4333",x"553f31",x"563f31",x"473a30",x"422c1f",x"422c1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"1b150e",x"1a130c",x"1a130c",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"180f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"191008",x"181008",x"180f08",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f08",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"180f08",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"333332",x"323232",x"323231",x"343434",x"343434",x"303030",x"343434",x"323232",x"343434",x"3d3c3c",x"3d3a39",x"3c3835",x"4a4643",x"4e4b49",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434141",x"474646",x"434343",x"444343",x"3e3c3b",x"343332",x"373534",x"363331",x"343332",x"353332",x"31302f",x"2d2c2c",x"000000",x"000000",x"515050",x"515050",x"343333",x"383533",x"333232",x"323130",x"323130",x"000000",x"4e4e4e",x"4e4e4e",x"2f2e2e",x"313131",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"221409",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331e0e",x"483223",x"544336",x"594232",x"583f2d",x"543c2b",x"533a2a",x"44372d",x"3f2819",x"3f2819",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"bcbcbc",x"bcbcbc",x"bcbcbc",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b140d",x"1b140d",x"1b150e",x"1b150e",x"19120c",x"19120c",x"17100a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"180f07",x"1a1008",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1d1108",x"1d1108",x"1e1208",x"1e1209",x"1e1208",x"1c1108",x"1c1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"201309",x"221409",x"241509",x"26160a",x"251509",x"251509",x"251509",x"26150a",x"28170a",x"2a180b",x"2a190b",x"2b190b",x"2a180b",x"28170b",x"27160a",x"251509",x"251509",x"25150a",x"26160a",x"25150a",x"211308",x"1d1007",x"221309",x"241509",x"231509",x"241509",x"241509",x"25150a",x"26170a",x"27170b",x"28170b",x"28170b",x"28180b",x"28180b",x"28170b",x"28170b",x"28170b",x"27170a",x"25160a",x"201308",x"201309",x"211409",x"221409",x"211409",x"211409",x"201309",x"201309",x"1f1309",x"1f1208",x"1f1208",x"1e1208",x"1c1108",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"1e1208",x"1d1108",x"1e1208",x"1f1208",x"1f1209",x"1f1209",x"1f1209",x"1f1309",x"1f1309",x"1f1309",x"201309",x"1f1309",x"211409",x"221509",x"221409",x"1f1309",x"1f1309",x"1f1309",x"1f1209",x"1e1209",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"180f08",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"2e2d2d",x"2d2c2c",x"333231",x"2e2b29",x"323232",x"303030",x"2f2f2f",x"313131",x"333333",x"353433",x"343332",x"3f3c39",x"4a4643",x"4e4b49",x"4b4845",x"504d4b",x"514f4d",x"454240",x"3c3a38",x"44413f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"55514f",x"433e3b",x"423e3b",x"434240",x"454544",x"323130",x"353434",x"343332",x"363433",x"393533",x"4d4c4b",x"353433",x"343333",x"333332",x"333332",x"000000",x"000000",x"484746",x"484746",x"353433",x"363433",x"343333",x"343332",x"343332",x"000000",x"4b4b4b",x"4b4b4b",x"2e2e2e",x"2e2e2e",x"323232",x"323232",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"666463",x"393939",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"343434",x"333333",x"000000",x"000000"),
(x"000000",x"331d0d",x"331d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1a0c",x"4d382a",x"544235",x"513c2f",x"583f2e",x"503727",x"4d3729",x"4d3b2e",x"4d311f",x"4d311f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"180f08",x"180f08",x"180f08",x"180f08",x"1a1008",x"28170b",x"351e0d",x"3c2310",x"38200f",x"402511",x"3e2410",x"3c2210",x"3f2310",x"402511",x"412411",x"422612",x"452813",x"422612",x"452814",x"462913",x"4b2b15",x"492a14",x"492a13",x"422611",x"482913",x"462913",x"412612",x"472913",x"422511",x"3a1f0d",x"341c0c",x"3d210e",x"402410",x"482a14",x"4b2b15",x"4b2c15",x"4b2d15",x"482a14",x"472812",x"482a13",x"462813",x"492a14",x"432711",x"3c210f",x"3e220f",x"452711",x"422511",x"402310",x"3e220f",x"40240f",x"40230f",x"3e220f",x"412410",x"422410",x"422511",x"432611",x"452813",x"482913",x"462711",x"432611",x"341d0c",x"3f230f",x"422510",x"422511",x"452812",x"422510",x"3f2410",x"432611",x"402410",x"432611",x"371e0d",x"3a1f0d",x"371d0c",x"3a1f0d",x"381e0c",x"371d0c",x"3b200d",x"3c210e",x"3f230f",x"371d0c",x"3a200e",x"3c210f",x"381f0e",x"3c210f",x"3e230f",x"3b210f",x"3c220f",x"381f0e",x"39200e",x"39200f",x"351e0d",x"3a210f",x"321d0d",x"29180b",x"1a1008",x"201309",x"241509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b150e",x"1b150e",x"19120c",x"19130c",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"1a1008",x"1e1208",x"231409",x"26160a",x"27170a",x"27170a",x"27170a",x"27170a",x"27170a",x"27160a",x"28170a",x"29180b",x"28180b",x"28180b",x"27170b",x"26160a",x"27170a",x"27170b",x"25160a",x"25150a",x"26160a",x"28170b",x"2b190b",x"2d1a0c",x"2c190b",x"29170a",x"2b180a",x"2c180b",x"2e1a0c",x"321d0d",x"331d0e",x"331d0e",x"331e0e",x"331d0d",x"311c0c",x"311c0d",x"301c0d",x"301c0d",x"2e1a0c",x"2b180b",x"2b180b",x"2d190b",x"2d190b",x"2a180a",x"29170a",x"29170a",x"29170a",x"2a170a",x"2b180b",x"2d190b",x"2e1a0c",x"301c0d",x"321d0d",x"301c0c",x"2f1b0c",x"2e1a0b",x"2d190b",x"2d190b",x"2e1a0c",x"2e1a0c",x"2d190b",x"2a180b",x"2b180b",x"2a180b",x"29170a",x"27160a",x"221409",x"221309",x"211308",x"211309",x"201208",x"1f1208",x"1d1108",x"1c1108",x"191008",x"170f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1c1108",x"1d1208",x"1e1208",x"1f1208",x"201309",x"221309",x"231409",x"251509",x"26160a",x"28170a",x"29180b",x"29180b",x"28170b",x"29180b",x"29180b",x"2a180b",x"29180b",x"29180b",x"28170a",x"27170a",x"26160a",x"2a190b",x"2c1a0b",x"29180b",x"27170b",x"27170a",x"26160a",x"26160a",x"26160a",x"25160a",x"25160a",x"25160a",x"24160a",x"24150a",x"231409",x"201308",x"201208",x"201309",x"201309",x"221409",x"23150a",x"221409",x"211409",x"1f1309",x"1c1108",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"180f07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"2e2d2d",x"2c2b2b",x"313131",x"303030",x"313131",x"303030",x"333333",x"343434",x"323131",x"333231",x"3b3734",x"3a3532",x"393431",x"3a3633",x"474340",x"504d4b",x"514f4d",x"454240",x"3c3a38",x"454341",x"403d3b",x"3e3c3b",x"444343",x"454343",x"454343",x"454343",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5d5b5a",x"54514f",x"56514e",x"55514f",x"3e3937",x"403c39",x"373433",x"343231",x"343231",x"363332",x"383534",x"363230",x"373533",x"585655",x"363332",x"323232",x"353332",x"333332",x"000000",x"000000",x"504b4a",x"504b4a",x"343231",x"343332",x"313131",x"353433",x"000000",x"000000",x"4f4e4e",x"4f4e4e",x"343433",x"333232",x"333333",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545453",x"666463",x"393939",x"323232",x"646464",x"575757",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f3f3f",x"383838",x"343434",x"323232",x"323232",x"333333",x"333333",x"000000"),
(x"000000",x"361f0e",x"361f0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1a0b",x"3c2414",x"584232",x"4f3a2c",x"51392b",x"543a29",x"523a2c",x"4c382b",x"533623",x"533623",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"180f07",x"180f07",x"180f08",x"191008",x"1c1108",x"1f1208",x"221409",x"24150a",x"24150a",x"25160a",x"211409",x"1f1309",x"201309",x"191008",x"191008",x"201309",x"24160a",x"27170b",x"25160a",x"27170a",x"26160a",x"28170a",x"29170a",x"27160a",x"28160a",x"251509",x"241409",x"221409",x"251509",x"261509",x"1e1208",x"251509",x"28170a",x"27170a",x"26160a",x"27160a",x"29170a",x"29180b",x"2f1c0d",x"24160a",x"2e1d0d",x"36200f",x"311d0e",x"311d0e",x"2d1a0c",x"2c1a0c",x"25160a",x"2f1b0c",x"321d0e",x"2d1a0c",x"301c0d",x"331e0e",x"311d0e",x"2e1b0c",x"2a180b",x"2c1a0c",x"311c0d",x"2d1a0c",x"2f1c0c",x"2d1a0b",x"2e1a0c",x"2b190b",x"2c180b",x"2c190b",x"29170a",x"2c190b",x"2a180b",x"241509",x"28170a",x"241509",x"2a180b",x"231509",x"241509",x"221409",x"27160a",x"2b180b",x"251509",x"231409",x"27160a",x"2b180b",x"231409",x"241509",x"25150a",x"25150a",x"24150a",x"1c1108",x"201309",x"231409",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"211409",x"25160a",x"41230f",x"432712",x"3f2411",x"3f2410",x"3d220f",x"3c220f",x"422611",x"412511",x"442712",x"3d2210",x"3e2310",x"432712",x"3c210f",x"3c220f",x"3a200e",x"3d220f",x"3f2411",x"432712",x"3e2411",x"442712",x"3b210f",x"3e2310",x"3c220f",x"3f2410",x"3c210e",x"371e0d",x"3d230f",x"402411",x"412511",x"432612",x"3f2410",x"432612",x"3e230f",x"3c220f",x"3d210f",x"371e0d",x"402411",x"3d230f",x"3d2310",x"3e2411",x"3e2310",x"3d2310",x"3b210f",x"351e0d",x"361d0d",x"381f0e",x"371e0d",x"321b0b",x"361e0d",x"361e0d",x"2c190b",x"402511",x"402511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1c150e",x"1c150e",x"19130c",x"19130c",x"19130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"191008",x"1e1208",x"221409",x"28170a",x"2c190b",x"2d190b",x"2f1b0c",x"301b0d",x"2f1b0c",x"311c0d",x"311d0d",x"321d0e",x"321d0e",x"311d0e",x"321d0d",x"2f1b0c",x"2e1a0c",x"2c190b",x"29180a",x"29170a",x"28170a",x"29170a",x"2a170a",x"2b180b",x"2c180a",x"2b180a",x"2c180b",x"301a0c",x"311c0c",x"321c0d",x"311c0c",x"2f1a0b",x"2f1a0b",x"331c0d",x"341f0e",x"331f0e",x"331e0e",x"33200f",x"36210f",x"351f0e",x"35200f",x"361f0f",x"361f0e",x"351f0e",x"351f0e",x"36200f",x"351f0f",x"37200f",x"37200f",x"37210f",x"371f0f",x"371f0e",x"3a210f",x"3b2210",x"3b2210",x"3a210f",x"38200e",x"38200f",x"361f0e",x"321c0c",x"341d0d",x"321c0c",x"321c0d",x"311c0c",x"2f1a0b",x"2f1b0c",x"2e1a0c",x"2b180b",x"28170a",x"27160a",x"251509",x"27170a",x"26160a",x"201308",x"1d1108",x"1d1108",x"1b1008",x"1a1008",x"1c1108",x"1d1108",x"1d1108",x"1d1208",x"1c1108",x"1a1008",x"1a1008",x"191008",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1c1108",x"1f1209",x"211309",x"221409",x"241509",x"251509",x"28170a",x"2c1a0c",x"2e1b0c",x"2e1a0c",x"301c0d",x"301b0d",x"2f1b0c",x"2e1a0c",x"2e1a0c",x"2e1a0b",x"301c0c",x"2e1a0c",x"2f1b0d",x"2d1a0b",x"2e1a0c",x"2d1a0c",x"2e1b0d",x"301d0c",x"301d0c",x"2f1b0c",x"2c190b",x"29180b",x"28170a",x"28170a",x"26160a",x"27160a",x"27160a",x"26160a",x"251509",x"251509",x"251509",x"241409",x"251509",x"26160a",x"27170a",x"27160a",x"25150a",x"241409",x"241509",x"231509",x"201409",x"1b1108",x"191008",x"160f07",x"150e07",x"150e07",x"150e07",x"160e07",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"4c4c4c",x"313131",x"313131",x"333333",x"333333",x"343333",x"363331",x"38322f",x"383432",x"3b3532",x"3a3531",x"3d3733",x"36322f",x"3a332f",x"332d29",x"373331",x"373331",x"393736",x"3a3736",x"444343",x"454343",x"464545",x"353434",x"444242",x"545454",x"555555",x"5a5959",x"5f5f5f",x"5f5f5f",x"616161",x"656565",x"595858",x"696969",x"656464",x"605f5f",x"635f5d",x"52514f",x"504b49",x"605d5b",x"3f3832",x"3b3633",x"3b3532",x"393533",x"373534",x"363433",x"373534",x"343231",x"373432",x"363534",x"3d3a39",x"4f4f4f",x"353535",x"353535",x"000000",x"000000",x"3a3838",x"313131",x"2f2e2e",x"303030",x"323131",x"323131",x"000000",x"000000",x"4d4c4c",x"4d4c4c",x"2f2f2e",x"2f2f2f",x"282828",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"323232",x"464646",x"323232",x"333333",x"646464",x"4d4d4d",x"4e4e4e",x"555555",x"595959",x"353434",x"3e3e3e",x"333231",x"353433",x"444343",x"686868",x"656565",x"5e5e5e",x"515151",x"3f3f3f",x"383838",x"3e3e3e",x"5f5f5f",x"333333",x"313131",x"323232",x"000000"),
(x"000000",x"351e0d",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d190b",x"4d382a",x"594536",x"533c2e",x"513727",x"543a29",x"4e372a",x"4b382b",x"523521",x"523521",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"170f07",x"180f07",x"1b1008",x"1f1208",x"241509",x"27160a",x"25150a",x"231409",x"231409",x"211309",x"1b1008",x"1c1108",x"241509",x"27170a",x"25150a",x"261509",x"241409",x"2a180b",x"29180b",x"2b190b",x"2d1b0c",x"2d1a0c",x"311c0d",x"221409",x"2b180b",x"211409",x"2d190b",x"28170a",x"261509",x"221309",x"231409",x"2e1a0c",x"2c1a0c",x"29180b",x"2c1a0c",x"2b190b",x"29170a",x"2c190b",x"29180b",x"2d190b",x"2e1a0c",x"2a180b",x"2d1a0b",x"2d1a0b",x"321d0d",x"2d1a0c",x"2d1a0c",x"2e1b0c",x"321d0d",x"351f0f",x"351f0f",x"311c0d",x"311d0d",x"2d1a0c",x"311c0d",x"331d0d",x"2c1a0c",x"2b190b",x"2f1b0c",x"26160a",x"26150a",x"27160a",x"29170a",x"2d1a0b",x"29180a",x"27170a",x"28170a",x"28170a",x"221409",x"221409",x"27160a",x"241509",x"27160a",x"241509",x"231409",x"231409",x"26160a",x"251509",x"1f1208",x"211309",x"231409",x"1d1108",x"1c1008",x"1e1108",x"1b1008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1e1208",x"221309",x"41230f",x"432712",x"3f2411",x"3f2410",x"3d220f",x"3c220f",x"422611",x"412511",x"442712",x"3d2210",x"3e2310",x"432712",x"3c210f",x"3c220f",x"3a200e",x"3d220f",x"3f2411",x"432712",x"3e2411",x"442712",x"3b210f",x"3e2310",x"3c220f",x"3f2410",x"3c210e",x"371e0d",x"3d230f",x"402411",x"412511",x"432612",x"3f2410",x"432612",x"3e230f",x"3c220f",x"3d210f",x"371e0d",x"402411",x"3d230f",x"3d2310",x"3e2411",x"3e2310",x"3d2310",x"3b210f",x"351e0d",x"361d0d",x"381f0e",x"371e0d",x"321b0b",x"361e0d",x"361e0d",x"2c190b",x"402511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1c150f",x"1c150e",x"1b140d",x"19130c",x"1a130c",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f07",x"191008",x"191008",x"191008",x"190f07",x"180f07",x"191008",x"191008",x"191008",x"191008",x"191008",x"180f08",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"3b3b3b",x"5b5b5b",x"555555",x"565656",x"323232",x"343433",x"333232",x"353230",x"383432",x"3e3835",x"393431",x"3b3633",x"38312d",x"342f2c",x"353230",x"383432",x"3b3633",x"373330",x"2e2a28",x"343332",x"383432",x"332117",x"333232",x"434342",x"545454",x"555555",x"5a5959",x"5f5f5f",x"5f5f5f",x"616161",x"656565",x"595858",x"696969",x"656464",x"5b5959",x"4e4946",x"3a3735",x"3a3633",x"393532",x"3a3532",x"363432",x"363331",x"373534",x"373534",x"343231",x"343231",x"333231",x"373737",x"343434",x"373737",x"3e3e3e",x"303030",x"313131",x"000000",x"000000",x"32302f",x"32302f",x"323131",x"313131",x"353332",x"353332",x"000000",x"000000",x"504f4f",x"504f4f",x"2f2e2e",x"313131",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"686867",x"333333",x"343434",x"343434",x"616161",x"5e5e5e",x"555555",x"505050",x"353434",x"333333",x"333231",x"353433",x"444343",x"4d4d4d",x"6b6b6b",x"5d5d5d",x"535353",x"424242",x"313131",x"303030",x"343434",x"312f2e",x"323131",x"323131",x"000000"),
(x"000000",x"38200f",x"38200f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"4a3527",x"4f3f33",x"503a2c",x"51392a",x"513929",x"513928",x"583f2e",x"492d1b",x"492d1b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"160e07",x"190f07",x"1e1208",x"24150a",x"29180b",x"2a180b",x"28170a",x"251509",x"241409",x"251509",x"201309",x"25160a",x"24150a",x"25150a",x"1d1208",x"29180b",x"2c190b",x"2b190b",x"2e1b0c",x"2b180b",x"2d1a0b",x"29180b",x"26160a",x"2b190b",x"27170a",x"29180b",x"25150a",x"26160a",x"26160a",x"26160a",x"241509",x"241509",x"1f1208",x"27160a",x"26160a",x"2b180b",x"251509",x"2b180b",x"2b180b",x"2d190b",x"29170a",x"2a180a",x"2b180b",x"2d190b",x"2e1b0c",x"2e1b0c",x"2c190c",x"2f1b0c",x"29170a",x"29170b",x"2d1a0b",x"2a180b",x"241509",x"29170a",x"2f1a0c",x"2f1c0d",x"2f1b0c",x"2e1b0c",x"2f1b0d",x"2d1a0c",x"2a190b",x"201309",x"2b190b",x"2a180b",x"29180b",x"2d1a0b",x"211409",x"251509",x"241509",x"25160a",x"2e1b0c",x"201309",x"231509",x"221309",x"221308",x"26160a",x"27160a",x"27170a",x"2c1a0b",x"29170b",x"231409",x"251509",x"211309",x"1e1209",x"191008",x"24160a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"211409",x"27170a",x"27170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"474545",x"4d4c4c",x"474747",x"3d3d3d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"393939",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1b140d",x"1b150e",x"1b150e",x"19130c",x"19120b",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f07",x"180f08",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"180f07",x"1a1008",x"1c1108",x"1d1208",x"1e1208",x"1e1208",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"191008",x"190f08",x"190f08",x"190f08",x"191008",x"191008",x"190f08",x"180f08",x"180f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f08",x"180f08",x"180f08",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"180f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"160e07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"323232",x"313131",x"343434",x"393939",x"565656",x"535353",x"4e4e4e",x"4a4949",x"35312f",x"373533",x"393532",x"353230",x"363330",x"343130",x"33302e",x"3a3532",x"353230",x"3c3633",x"32302f",x"3a3633",x"343332",x"343231",x"353433",x"373331",x"353433",x"343231",x"323232",x"333333",x"3a3a3a",x"3f3f3f",x"484848",x"484848",x"373432",x"342b25",x"373534",x"333333",x"413730",x"373432",x"3d3632",x"403832",x"38322f",x"393431",x"3a3532",x"363432",x"383432",x"363636",x"333333",x"363636",x"323232",x"313131",x"323232",x"2e2f2f",x"323232",x"2e2e2e",x"2f2f2f",x"000000",x"323131",x"323131",x"343332",x"313030",x"31241c",x"323232",x"000000",x"000000",x"575757",x"535353",x"3a3a3a",x"323232",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"5b5b5b",x"333333",x"323232",x"343434",x"333333",x"5f5f5f",x"313131",x"313131",x"333333",x"343333",x"333232",x"373534",x"343333",x"323232",x"343333",x"343434",x"333333",x"323232",x"333333",x"333333",x"373737",x"333333",x"312f2e",x"323131",x"323131",x"000000"),
(x"000000",x"2e1a0b",x"2e1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301b0b",x"4c392c",x"604839",x"5b4333",x"5b402d",x"513a2a",x"4e3829",x"523d2d",x"4e3220",x"4e3220",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"160f07",x"191008",x"1f1208",x"221409",x"29170b",x"2b180b",x"2a180b",x"29170b",x"28170a",x"25160a",x"26160a",x"1f1208",x"1e1108",x"1c1108",x"1e1108",x"231409",x"231409",x"27160a",x"29170a",x"2b180b",x"231409",x"251509",x"261509",x"28160a",x"27160a",x"2b190b",x"2c1a0b",x"29180b",x"2b180b",x"221409",x"27160a",x"27160a",x"29170a",x"1f1209",x"221409",x"2c190b",x"221409",x"2d190b",x"2b180b",x"28160a",x"26150a",x"28160a",x"28160a",x"2b180b",x"29170b",x"2d1a0c",x"2a180b",x"2f1b0c",x"29180b",x"331d0e",x"2d1a0c",x"2a180b",x"251509",x"251509",x"29170a",x"2f1b0c",x"2e1b0c",x"2e1b0c",x"2b180b",x"26150a",x"2a180b",x"2e1a0b",x"2d1a0c",x"29180b",x"2d190b",x"26160a",x"29170b",x"29170a",x"26160a",x"29170b",x"26160a",x"24150a",x"1f1309",x"241509",x"201309",x"2b190b",x"28170b",x"2a190b",x"26160a",x"2a180b",x"26160a",x"26170a",x"22150a",x"1e1209",x"150e07",x"180f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f08",x"211409",x"26160a",x"26160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"605e5e",x"605f5f",x"4e4d4d",x"4d4c4c",x"474747",x"3d3d3d",x"323232",x"333332",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"505050",x"4a4746",x"515151",x"4c4c4b",x"393939",x"353535",x"353535",x"343434",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"454545",x"535353",x"545454",x"424242",x"323232",x"333333",x"333333",x"434343",x"3a3a3a",x"323232",x"333333",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"1c150e",x"1c150e",x"1b140e",x"19120b",x"19120b",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"180f07",x"190f08",x"191008",x"190f08",x"180f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"170f07",x"191008",x"1d1108",x"201309",x"221409",x"221409",x"221409",x"211309",x"201309",x"201309",x"201309",x"201309",x"201309",x"1f1209",x"1f1209",x"1f1209",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1d1108",x"1d1208",x"1d1108",x"1d1208",x"1d1208",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"180f08",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f08",x"190f08",x"180f07",x"180f07",x"180f07",x"180f08",x"180f08",x"180f08",x"180f08",x"190f08",x"191008",x"180f07",x"180f08",x"180f07",x"190f08",x"191008",x"1b1107",x"180f07",x"181007",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"343434",x"2c2c2c",x"313131",x"303030",x"323232",x"292929",x"2d2d2d",x"323131",x"4a4848",x"454444",x"464543",x"34302e",x"353230",x"363230",x"393533",x"353230",x"363330",x"383432",x"393532",x"373332",x"383432",x"363433",x"323131",x"353433",x"343332",x"343333",x"323232",x"303030",x"333232",x"313131",x"333333",x"333333",x"313131",x"313131",x"353332",x"3c3a39",x"52514f",x"4f4e4d",x"3e3b39",x"413c38",x"3b3632",x"383432",x"363332",x"3b3532",x"3a3a3a",x"3b3b3b",x"323232",x"272828",x"343434",x"313131",x"323232",x"2b2c2c",x"2f2f2f",x"303030",x"2c2c2c",x"2c2c2c",x"000000",x"363331",x"363331",x"33312f",x"333231",x"31302f",x"31302f",x"000000",x"000000",x"4e4e4e",x"4e4e4e",x"333333",x"323232",x"2f2f2f",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"343434",x"4b4b4b",x"555555",x"4d4d4d",x"323232",x"303030",x"313131",x"333333",x"323130",x"353432",x"333232",x"313131",x"323232",x"333333",x"323232",x"323232",x"343434",x"373737",x"323232",x"323232",x"000000",x"000000",x"000000"),
(x"000000",x"2d1a0b",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"523d2e",x"665040",x"5e4636",x"5c4331",x"573d2c",x"533b2b",x"553d2f",x"472f1f",x"472f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"160f07",x"1b1108",x"201309",x"24150a",x"27160a",x"2b180b",x"2d1a0b",x"2e1b0c",x"2b190b",x"28180b",x"231509",x"22150a",x"191008",x"28170b",x"2c1a0c",x"2a190b",x"311c0d",x"2a190b",x"2c1a0b",x"2b190b",x"2b180b",x"29180b",x"2e1b0c",x"311c0d",x"2c1a0c",x"2a180b",x"2a180b",x"211409",x"2b190b",x"2d1a0c",x"241509",x"28160a",x"1f1209",x"2e1a0b",x"25160a",x"24150a",x"2c1a0c",x"2a180b",x"2b190c",x"301c0d",x"2d1a0c",x"2b190b",x"321d0d",x"2d1a0c",x"311c0d",x"2c1a0b",x"2e1b0c",x"301c0d",x"2d1a0c",x"27170b",x"2a180b",x"25150a",x"2b180b",x"26170b",x"2a1a0c",x"2e1b0d",x"301c0d",x"2e1b0d",x"2c1a0c",x"2d1b0c",x"2d1b0c",x"2b190c",x"2c1a0c",x"2c1a0c",x"2d1a0c",x"2e1b0c",x"27170a",x"2d1a0b",x"2b190b",x"29170a",x"26160a",x"201309",x"29180b",x"27170a",x"29180b",x"26160a",x"29170b",x"28170a",x"211409",x"241509",x"25160a",x"29180b",x"221409",x"201209",x"160f07",x"191008",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"24150a",x"2a190b",x"2a190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e5e5d",x"5f5d5d",x"616060",x"545252",x"5d5c5c",x"5a5959",x"4c4b4b",x"323131",x"343333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"333333",x"000000",x"616160",x"595959",x"323232",x"333333",x"000000",x"5c5c5c",x"5d5d5d",x"5a5a5a",x"4a4746",x"515151",x"4c4c4b",x"4c4c4c",x"4a4a4a",x"3d3d3d",x"323232",x"323232",x"333333",x"313232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"444444",x"434343",x"363636",x"484848",x"414141",x"454545",x"565656",x"515151",x"4a4a4a",x"333333",x"323232",x"323232",x"494949",x"3a3a3a",x"323232",x"333333",x"323232",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"1b140d",x"1b140d",x"1b150e",x"19120c",x"19120b",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"171009",x"171009",x"171009",x"17110a",x"171009",x"171009",x"17100a",x"171009",x"171009",x"17110a",x"17100a",x"17100a",x"171009",x"17110a",x"17110a",x"17110a",x"17100a",x"17110a",x"171009",x"171009",x"171009",x"171009",x"17110a",x"17110a",x"171009",x"171009",x"17110a",x"17110a",x"17110a",x"17110a",x"171009",x"17110a",x"171009",x"17110a",x"171009",x"171009",x"171009",x"171009",x"171009",x"171009",x"171009",x"17110a",x"171009",x"171009",x"171009",x"171009",x"17110a",x"17110a",x"17110a",x"171009",x"171009",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"303030",x"313131",x"333333",x"2e2e2e",x"5e5e5e",x"313131",x"313131",x"333231",x"363433",x"383635",x"474544",x"494847",x"484745",x"42403f",x"4b4a49",x"393431",x"363330",x"383432",x"373331",x"373332",x"363230",x"333232",x"353333",x"343332",x"333232",x"333232",x"303030",x"343434",x"404040",x"4a4a4a",x"515151",x"515151",x"514e4c",x"524f4d",x"515050",x"555454",x"595553",x"545251",x"403f3e",x"3c3835",x"3b3532",x"4d4d4d",x"4e4e4e",x"414141",x"313131",x"39261d",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"2f2f2f",x"323232",x"333333",x"303030",x"000000",x"363331",x"383432",x"2f2c2a",x"35312e",x"2a2a28",x"2a2a28",x"000000",x"000000",x"343434",x"343434",x"2f2f2f",x"292929",x"323232",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"565656",x"3e3e3e",x"323232",x"323232",x"323232",x"333333",x"333232",x"343331",x"313030",x"313131",x"333333",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"311b0c",x"311b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"241309",x"462f21",x"604a3c",x"584032",x"5a3f2d",x"5b3c29",x"573d2b",x"483223",x"4c311e",x"4c311e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"160f07",x"1a1008",x"201309",x"26160a",x"29170a",x"2d1a0b",x"2d1a0b",x"2c190b",x"28170a",x"231509",x"201309",x"27160a",x"26160a",x"25160a",x"29180b",x"27160a",x"29180b",x"24150a",x"25150a",x"2a190b",x"2c1a0c",x"2e1b0d",x"2e1b0c",x"2f1b0c",x"29180b",x"2c190b",x"2e1b0c",x"29180b",x"29180b",x"2b190b",x"28170b",x"29180b",x"27170a",x"2a190b",x"28180b",x"29170b",x"2a180b",x"29180b",x"25160a",x"2c190c",x"361f0f",x"2b190c",x"2b190b",x"331d0e",x"2f1b0c",x"2b190b",x"311c0d",x"301c0d",x"311d0e",x"2b190c",x"2a190c",x"301c0d",x"2d1b0c",x"2a180b",x"2c1a0c",x"28180b",x"2c1a0c",x"2c1a0c",x"27170b",x"2a180b",x"2e1a0c",x"26160a",x"28180b",x"29180b",x"2d1a0c",x"2f1b0d",x"27170a",x"2a180b",x"29180b",x"29180b",x"28170a",x"26160a",x"28180b",x"211309",x"2a190b",x"29180b",x"27160a",x"29170a",x"201309",x"24150a",x"23150a",x"28170b",x"211409",x"201309",x"1c1108",x"1c1108",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"180f08",x"221409",x"28170b",x"28170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"605f5f",x"5d5d5c",x"5e5e5d",x"5a5856",x"575656",x"4c4b4b",x"535252",x"494949",x"535151",x"323232",x"303030",x"333232",x"000000",x"000000",x"5b5a59",x"383737",x"333333",x"333333",x"5c5b5a",x"595959",x"323232",x"333333",x"585858",x"5d5d5d",x"606060",x"636363",x"5c5c5c",x"474747",x"303030",x"464646",x"565656",x"5c5c5c",x"656565",x"484848",x"323232",x"333333",x"323232",x"333333",x"000000",x"000000",x"616161",x"545454",x"474747",x"434343",x"3a3a3a",x"484848",x"494949",x"545454",x"424242",x"434343",x"494949",x"4f4f4f",x"333333",x"3c3c3c",x"454545",x"5a5a5a",x"3d3d3d",x"333333",x"333333",x"323232",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c150e",x"1c150e",x"1b150e",x"1b140d",x"1b150e",x"1a130c",x"19120c",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"17110a",x"17100a",x"17110a",x"17110a",x"171009",x"171009",x"17110a",x"171009",x"17110a",x"17110a",x"171009",x"17110a",x"171009",x"17110a",x"17110a",x"17110a",x"17110a",x"17110a",x"171009",x"17100a",x"171009",x"171009",x"171009",x"17100a",x"171009",x"171009",x"171009",x"171009",x"17110a",x"171009",x"17110a",x"17110a",x"171009",x"171009",x"171009",x"171009",x"171009",x"171009",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"363432",x"363432",x"3d3d3d",x"323232",x"31302f",x"333333",x"302d2c",x"343231",x"353332",x"322f2d",x"363332",x"454443",x"42403f",x"4f4d4d",x"515050",x"565656",x"5b5b5b",x"000000",x"000000",x"353332",x"333232",x"343332",x"343332",x"333232",x"333232",x"303030",x"343434",x"3c3c3c",x"4d4d4d",x"525252",x"515151",x"4e4e4e",x"545351",x"4f4e4e",x"444342",x"484645",x"474545",x"464646",x"5c5b5b",x"444444",x"333333",x"323232",x"333333",x"333333",x"2b2b2b",x"313131",x"343434",x"2f2219",x"323131",x"333333",x"313131",x"363432",x"373533",x"363331",x"000000",x"000000",x"3a3736",x"3a3736",x"3a3633",x"363230",x"342f2d",x"211f1d",x"000000",x"000000",x"3e3e3e",x"323232",x"2f2f2f",x"323232",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a3a3a",x"616161",x"5c5c5c",x"616161",x"525252",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"333232",x"343331",x"313030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"331c0c",x"331c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"261409",x"533e31",x"5d493a",x"573f2f",x"5d402b",x"563826",x"573a27",x"463123",x"52321c",x"52321c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"181007",x"181007",x"170f07",x"1a1108",x"201409",x"27170b",x"2a180b",x"2c190b",x"2f1b0c",x"2e1b0d",x"2c1a0c",x"26160a",x"211409",x"27170b",x"25160a",x"29180b",x"26160a",x"27170b",x"180f08",x"28170b",x"2a190b",x"2e1b0c",x"2c190b",x"2c190b",x"2d1a0b",x"2c190b",x"2e1b0c",x"2f1b0d",x"311c0d",x"2e1b0c",x"2b190b",x"2e1a0c",x"331e0e",x"27170b",x"22150a",x"2b190b",x"2c190b",x"2f1b0d",x"301c0d",x"311c0d",x"2f1c0d",x"311c0d",x"341e0e",x"29170b",x"2a180b",x"2d1a0c",x"311c0d",x"311c0d",x"301c0d",x"2d1a0c",x"301c0d",x"2f1b0c",x"2f1b0c",x"321d0e",x"321d0e",x"331e0e",x"351f0f",x"321d0e",x"341f0f",x"301c0d",x"2d1a0c",x"2c190c",x"2f1c0d",x"321d0d",x"311c0d",x"2c190b",x"2e1b0c",x"2e1b0c",x"2f1b0c",x"2d1a0b",x"26160a",x"2b190b",x"28170a",x"26160a",x"251509",x"26160a",x"24150a",x"29180b",x"2a180b",x"26160a",x"29180b",x"241509",x"201309",x"241509",x"27170a",x"1e1209",x"24150a",x"1c1108",x"1c1108",x"1a1108",x"180f08",x"160e07",x"150e07",x"150e07",x"1a1008",x"23150a",x"29180b",x"29180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"666564",x"646363",x"6a6969",x"343433",x"383533",x"383735",x"565555",x"535353",x"4e4d4d",x"363534",x"323232",x"343333",x"474747",x"3a3a3a",x"616060",x"5b5a59",x"313131",x"5d5d5d",x"515151",x"575757",x"303030",x"333333",x"5d5d5d",x"5a5a5a",x"5e5e5e",x"2c2c2d",x"382820",x"2f3030",x"323232",x"3f3f40",x"4a4a4a",x"535353",x"655f5d",x"585757",x"606060",x"323232",x"323232",x"333333",x"000000",x"646464",x"656565",x"5a5a5a",x"505050",x"5b5b5b",x"5a5a5a",x"4f4f4f",x"484848",x"414141",x"464646",x"4c4c4c",x"454545",x"3c3c3c",x"494949",x"4c4c4c",x"494949",x"4b4b4b",x"454545",x"494949",x"4f4f4f",x"353535",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b150e",x"1b150e",x"1c160f",x"1b150e",x"1b140d",x"1a140d",x"19120c",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"17100a",x"171009",x"171009",x"17110a",x"171009",x"171009",x"17110a",x"17110a",x"171009",x"171009",x"171009",x"171009",x"17100a",x"17110a",x"171009",x"171009",x"17110a",x"171009",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"363332",x"353331",x"343230",x"5d5956",x"605e5c",x"5e5d5c",x"393939",x"333232",x"343231",x"363433",x"353231",x"32302f",x"332e2c",x"353332",x"4f4e4e",x"525151",x"565656",x"5b5b5b",x"575757",x"5b5a5a",x"646464",x"595959",x"606060",x"5e5e5e",x"5b5b5b",x"5a5a5a",x"5b5b5b",x"4b4b4b",x"4a4a4a",x"464545",x"434242",x"515050",x"4d4c4c",x"4b4a49",x"3f3e3e",x"353433",x"343231",x"343332",x"313131",x"323232",x"303030",x"313131",x"333333",x"313131",x"333333",x"313131",x"333333",x"252525",x"313131",x"3a332f",x"39332f",x"363230",x"373534",x"363331",x"373533",x"000000",x"4f4d4a",x"4f4d4a",x"3c3938",x"433a33",x"353332",x"383331",x"383331",x"000000",x"000000",x"323232",x"323232",x"313131",x"313131",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"333333",x"3a3a3a",x"616161",x"5c5c5c",x"616161",x"525252",x"4c4c4c",x"525252",x"585858",x"5c5c5c",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2d190b",x"2d190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251409",x"4a3223",x"5a4537",x"593f2e",x"523727",x"573926",x"5b3b25",x"483021",x"4c301a",x"4c301a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c1108",x"1c1108",x"1c1108",x"180f08",x"1d1208",x"231509",x"28170a",x"2a180a",x"2a180a",x"28170a",x"251509",x"201208",x"221309",x"201309",x"241509",x"201309",x"28170b",x"29180b",x"211409",x"2d1b0d",x"2f1c0d",x"2f1c0d",x"311d0e",x"2e1b0d",x"2f1b0d",x"311c0d",x"311c0d",x"321d0d",x"2d1a0c",x"321c0d",x"2e1b0c",x"2f1b0c",x"341f0f",x"321e0e",x"331f0f",x"2d1a0d",x"311d0e",x"2c1a0c",x"311c0d",x"2d1a0c",x"2d190b",x"2e1a0c",x"2b190b",x"351f0e",x"2b190c",x"2f1b0d",x"331d0e",x"341e0e",x"2c1a0c",x"29180b",x"29180b",x"2c190c",x"2c190b",x"2e1b0c",x"321e0e",x"331f0f",x"321d0e",x"331e0e",x"321d0e",x"321d0e",x"301c0d",x"311d0d",x"36200f",x"2e1b0c",x"321d0d",x"28160a",x"301b0c",x"2f1b0c",x"331d0d",x"2e1b0c",x"2d1a0c",x"2a180a",x"261509",x"29170a",x"27160a",x"27170a",x"28170a",x"25150a",x"241509",x"251509",x"211308",x"231409",x"261509",x"28170a",x"2a190b",x"25160a",x"211409",x"211409",x"211309",x"1f1208",x"1b1008",x"170f07",x"150e07",x"150e07",x"180f07",x"211309",x"26160a",x"26160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"686564",x"666564",x"686767",x"353433",x"343333",x"373533",x"5a5959",x"5f5d5c",x"575554",x"504f4f",x"595858",x"333333",x"323232",x"474747",x"424242",x"4f4f4f",x"5e5e5e",x"323232",x"4d4d4d",x"505050",x"4c4d4d",x"323232",x"353535",x"575757",x"5a5a5a",x"2d2d2d",x"303030",x"323232",x"303030",x"313131",x"3f3f40",x"4a4a4a",x"545454",x"585757",x"414141",x"464646",x"616161",x"333333",x"333333",x"5f5f5f",x"656564",x"5f5f5f",x"535353",x"4b4b4b",x"515151",x"424242",x"494949",x"424242",x"373737",x"464646",x"4e4e4e",x"4b4b4b",x"484848",x"424242",x"454545",x"484848",x"4a4a4a",x"3f3f3f",x"4a4a4a",x"515151",x"5a5a5a",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1610",x"1d1610",x"1d1610",x"1c150f",x"1c150e",x"1b150e",x"1a130c",x"19120b",x"171009",x"17100a",x"150e07",x"150e07",x"150e07",x"1b130b",x"1e130b",x"2a1c12",x"2c1e15",x"332316",x"372517",x"3b2617",x"3d2819",x"3f2816",x"3b2515",x"3e2817",x"422a18",x"412817",x"3b2516",x"3c2617",x"3d2515",x"3e2515",x"412717",x"422716",x"442916",x"482c17",x"4a2e18",x"4c2f19",x"4e301a",x"4b2e19",x"4d2f1a",x"4b2e1b",x"4b2d19",x"4b2e1a",x"4b2e1a",x"492d1a",x"472c19",x"492e1c",x"462b19",x"4e321d",x"4e321e",x"4e331d",x"4c311d",x"4d321d",x"4b301c",x"492d1a",x"472d1b",x"482d1a",x"452c1a",x"4b301c",x"4d311c",x"4d301b",x"4a2e1b",x"4c2e19",x"4c2f1a",x"482c19",x"472c19",x"472c19",x"492d18",x"492d19",x"50311c",x"51341e",x"52361f",x"533620",x"543620",x"513621",x"513620",x"4f3321",x"4e321f",x"4e331e",x"49301f",x"472f1f",x"462e1f",x"4b3120",x"4a3220",x"4c3322",x"49301f",x"4d3320",x"472f1f",x"432d1e",x"482f1f",x"4c3321",x"4a321f",x"4a3222",x"4b3321",x"452f1f",x"452f20",x"432d1f",x"3f2a1d",x"422e20",x"432e1f",x"463020",x"453020",x"443021",x"453022",x"432f20",x"423023",x"3e2c1f",x"2c1e15",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"363534",x"363432",x"353331",x"383432",x"332f2c",x"373331",x"666564",x"504c49",x"53504d",x"353332",x"353332",x"353332",x"302f2e",x"363534",x"353433",x"333332",x"353434",x"323232",x"383838",x"515151",x"5b5b5b",x"585858",x"595959",x"5f5f5f",x"5e5e5e",x"5b5b5b",x"5b5b5b",x"5b5b5b",x"4b4b4b",x"4a4a4a",x"343434",x"343333",x"343332",x"353433",x"38271e",x"333232",x"353433",x"353433",x"323232",x"2f2f2f",x"313131",x"343434",x"323232",x"333333",x"303030",x"2a2a2a",x"323232",x"39312c",x"3e3732",x"3b3532",x"3e3733",x"3b3532",x"353230",x"353331",x"353332",x"343231",x"2f2d2b",x"000000",x"565351",x"56514f",x"352f2b",x"343231",x"333231",x"333231",x"000000",x"000000",x"2f2f2f",x"2f2f2f",x"282929",x"333434",x"2c1d0f",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"323232",x"333333",x"313131",x"323231",x"2f3030",x"4f4440",x"646363",x"4e4e4e",x"525252",x"585858",x"5c5c5c",x"333333",x"333333",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2f1a0b",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251409",x"513b2d",x"5a4536",x"5c412f",x"533928",x"563827",x"553827",x"483325",x"4d301d",x"4d301d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221508",x"221508",x"231608",x"201509",x"1d1208",x"25160a",x"2b190b",x"311d0d",x"311c0d",x"2d1a0c",x"2b190c",x"27170b",x"1e1208",x"1c1108",x"211409",x"221409",x"25160a",x"27170b",x"27170b",x"25160a",x"2b180b",x"28170a",x"2c190b",x"2b180b",x"2b180b",x"2e1a0b",x"2d190b",x"2e1a0b",x"2b180a",x"29170a",x"2e1a0b",x"2b190b",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"27170a",x"2a180b",x"2c1a0c",x"27170b",x"2c1a0c",x"2c190c",x"29180b",x"221409",x"2a190b",x"2c1a0c",x"2a180b",x"28170b",x"2d1a0c",x"2e1b0c",x"2f1c0d",x"29180b",x"2a180b",x"2b180b",x"2a180b",x"2d190b",x"2a180b",x"2d1a0b",x"2d1a0b",x"2d1a0b",x"2e1a0c",x"2c190b",x"2c190b",x"2d190b",x"2d190b",x"2c190b",x"2d190b",x"2b180b",x"2c190b",x"28170a",x"2b180b",x"271609",x"251509",x"241409",x"241409",x"221308",x"1d1108",x"1f1108",x"1c1108",x"1d1108",x"211308",x"241409",x"211309",x"231409",x"221409",x"221409",x"221409",x"221409",x"241409",x"231409",x"221309",x"1e1208",x"191008",x"160f07",x"150e07",x"191008",x"24150a",x"29180b",x"29180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"6b6764",x"6b6764",x"565554",x"333231",x"333231",x"000000",x"5e5c5b",x"5e5c5b",x"565454",x"545252",x"4b4b4b",x"575656",x"696969",x"6b6b6b",x"5e5e5e",x"585858",x"4f4f4f",x"494949",x"484848",x"4c4c4c",x"515151",x"545454",x"4f4f4f",x"505151",x"333333",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"464646",x"5c5b5b",x"5a5a5a",x"434343",x"333333",x"535353",x"5b5b5b",x"404040",x"313131",x"323232",x"333333",x"313131",x"484848",x"323232",x"323232",x"343434",x"444444",x"484848",x"515151",x"505050",x"4c4c4c",x"4e4e4e",x"505050",x"535353",x"4d4d4d",x"3f3f3f",x"373737",x"444444",x"373737",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d160f",x"1d160f",x"1d1710",x"1d1610",x"1b140e",x"1b150e",x"19120b",x"19120b",x"17110a",x"17100a",x"150e07",x"150e07",x"150e07",x"51463c",x"51473d",x"493e34",x"44362a",x"403328",x"413226",x"413226",x"453528",x"463528",x"48372a",x"4a382b",x"4a382a",x"4e3b2c",x"48362a",x"49382d",x"4d3c2f",x"4e3c30",x"4c3b2f",x"514034",x"4c3a2c",x"564539",x"5a4a3d",x"554537",x"57473b",x"534133",x"523f32",x"4f3c2e",x"4f3b2d",x"513c2e",x"4d3a2c",x"4b3b2f",x"4a3a2e",x"4a392d",x"48362a",x"4b392b",x"4a3729",x"493628",x"4b382b",x"4d392c",x"4b382a",x"4b382a",x"4c382a",x"4f3b2c",x"4e3b2c",x"503b2c",x"4e392b",x"4c3829",x"513f30",x"533f31",x"544133",x"574333",x"574334",x"544132",x"544235",x"523e30",x"523f31",x"503b2d",x"4e392a",x"4d3828",x"4c3727",x"4d3829",x"4f3a2b",x"4c382a",x"4e3a2c",x"4f3d30",x"4e3c2f",x"48382b",x"4a392b",x"49362a",x"493729",x"48362a",x"49372a",x"48362a",x"453428",x"453427",x"483628",x"423225",x"413026",x"3f2f24",x"3d2e24",x"3d2d22",x"3f3126",x"3f3025",x"3e3025",x"3c2f25",x"3c2f26",x"3d3126",x"392f26",x"342a21",x"342a21",x"3a2e24",x"3b2e24",x"40352b",x"4c4239",x"564d43",x"554b40",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"160e07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"322f2e",x"322f2e",x"35312e",x"383432",x"363332",x"363331",x"363433",x"373432",x"383431",x"44403d",x"514e4c",x"353433",x"333332",x"343433",x"333232",x"323232",x"303030",x"323232",x"343434",x"323232",x"313131",x"343434",x"313131",x"303030",x"323232",x"333333",x"313131",x"2f2f2f",x"333333",x"323232",x"343332",x"353434",x"333231",x"343333",x"323131",x"333232",x"333333",x"343434",x"313131",x"313131",x"333333",x"535353",x"323232",x"333333",x"3c342f",x"3b342f",x"3f362f",x"423831",x"3c3633",x"3a3531",x"3b3632",x"393533",x"383431",x"373331",x"302f2e",x"322f2e",x"322f2e",x"000000",x"51504e",x"51504e",x"342d29",x"353230",x"383532",x"383532",x"000000",x"000000",x"343434",x"343434",x"333333",x"313131",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"3e3e3e",x"343434",x"323232",x"333333",x"323232",x"333333",x"343535",x"353535",x"323232",x"333333",x"303030",x"313131",x"494745",x"333333",x"323232",x"333333",x"323232",x"323232",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"301a0b",x"301a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"221308",x"4f392a",x"594437",x"5f432f",x"533b2b",x"5a3f2d",x"583d2d",x"513829",x"4e301c",x"4e301c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231608",x"231608",x"231608",x"231609",x"1d1208",x"211409",x"251509",x"28170a",x"2b190b",x"2a180b",x"28170a",x"24150a",x"1f1309",x"1c1108",x"1e1209",x"201309",x"201309",x"22150a",x"24150a",x"28170b",x"2b190c",x"2d1a0c",x"2e1b0c",x"301c0d",x"311c0d",x"321d0d",x"311c0d",x"311c0d",x"2e1a0c",x"2f1b0c",x"2f1b0d",x"2c190b",x"2c190b",x"2d1b0c",x"2e1b0d",x"2d1b0c",x"2b190c",x"29180b",x"29190b",x"2a190b",x"2b190c",x"2a190b",x"2a190b",x"29180b",x"311c0d",x"2c1a0c",x"2a190c",x"29180b",x"26160a",x"201309",x"211309",x"231409",x"28170b",x"2d1a0c",x"2d1a0c",x"301c0d",x"311c0d",x"311c0d",x"301c0d",x"321d0e",x"2f1b0c",x"2d1a0b",x"2b180b",x"29170a",x"2f1b0c",x"2f1b0c",x"2f1c0c",x"2e1a0c",x"2e1a0c",x"2b190b",x"29180a",x"261509",x"261509",x"241409",x"241509",x"221409",x"201309",x"201208",x"1f1208",x"201308",x"221409",x"251509",x"28170a",x"29180b",x"2a180b",x"29170b",x"28170a",x"251509",x"221309",x"221409",x"201308",x"1d1208",x"181008",x"160e07",x"1a1008",x"24150a",x"2a180b",x"2a180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"615d59",x"615d59",x"4a4744",x"373331",x"373331",x"000000",x"616060",x"616060",x"565656",x"504e4e",x"323131",x"333332",x"343333",x"434343",x"494949",x"515151",x"535353",x"474747",x"464646",x"484848",x"414141",x"444444",x"444444",x"464646",x"414141",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"383838",x"383838",x"313131",x"333333",x"555453",x"5a5958",x"565656",x"333333",x"4f4f4f",x"454545",x"313131",x"333333",x"323232",x"323232",x"323232",x"383838",x"323232",x"333333",x"393939",x"4a4a4a",x"4a4a4a",x"4d4d4d",x"434343",x"474747",x"454545",x"4c4c4c",x"3a3a3a",x"333333",x"323232",x"323232",x"414141",x"3c3c3c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1d1710",x"1c160f",x"1b150e",x"1b150e",x"1b150e",x"19130c",x"171009",x"18110a",x"150e07",x"150e07",x"150e07",x"51473d",x"52483e",x"4c3f33",x"45382c",x"3e3126",x"413326",x"3f3024",x"433325",x"443326",x"463629",x"453528",x"4a3829",x"47372a",x"433227",x"443429",x"4a3a2e",x"4c3b2e",x"49392d",x"4a392d",x"4d3d31",x"504034",x"534337",x"58473a",x"574639",x"544033",x"533f31",x"543f30",x"543e2e",x"543e2d",x"533f30",x"4f3c2d",x"4a382a",x"4a3729",x"473427",x"473426",x"473426",x"493527",x"4a3728",x"4e3829",x"4c3728",x"4d382a",x"4c3829",x"4a3526",x"4c3829",x"4d3829",x"513d2c",x"523d2d",x"523c2d",x"4e3a2a",x"4f3b2e",x"4f3b2d",x"4e3b2c",x"4f3c2e",x"523e30",x"523d2d",x"533f2f",x"503a2b",x"4e392a",x"503a2b",x"503928",x"503a29",x"513a2b",x"4e3828",x"4d392b",x"4f3c2f",x"4e3b2d",x"4c3b2e",x"4d3b2e",x"4d3a2c",x"4b3829",x"4b3729",x"4c382a",x"4a3628",x"4b3728",x"4a3729",x"473528",x"483527",x"413125",x"3f2f22",x"3f3025",x"413125",x"3e2e24",x"3f3125",x"3b2d22",x"3e3126",x"3d3026",x"3c2e24",x"3a2e25",x"382d24",x"342a22",x"362b22",x"372c22",x"3c2f25",x"493f36",x"564b41",x"594f45",x"594f45",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"322f2e",x"322f2d",x"353230",x"393633",x"373330",x"4f4c4a",x"3a3633",x"393431",x"3b3532",x"3c3531",x"3b342f",x"403731",x"4e4946",x"313131",x"313131",x"323232",x"3a3a3a",x"444444",x"505050",x"515151",x"575757",x"555555",x"4c4c4c",x"343434",x"323232",x"3b3b3b",x"323232",x"4c4c4c",x"454545",x"342e2a",x"313131",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"333333",x"333333",x"5c5451",x"554e4a",x"544f4c",x"47403c",x"3b3531",x"403731",x"3e3632",x"3d3531",x"3b342f",x"362c25",x"39312c",x"3a3633",x"39322e",x"393431",x"363331",x"302d2c",x"353332",x"322f2e",x"474442",x"474442",x"46423f",x"393533",x"35312f",x"383432",x"383432",x"000000",x"000000",x"323232",x"323232",x"333333",x"323232",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"3c3c3c",x"5c5b5b",x"4d4d4d",x"323232",x"323232",x"323232",x"333333",x"323131",x"333333",x"323232",x"313130",x"454342",x"605f5d",x"393939",x"323232",x"3c3c3c",x"353535",x"323232",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2e1a0b",x"2e1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"271509",x"473021",x"604533",x"59402f",x"543e30",x"583f2f",x"543c2c",x"513b2c",x"4e301c",x"4e301c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1a0a",x"2a1a0a",x"2c1b0a",x"201409",x"1e1308",x"211509",x"28170b",x"2b190c",x"2d1a0c",x"2c1a0c",x"28180b",x"25160b",x"201309",x"1f1309",x"201409",x"211409",x"22150a",x"231509",x"25150a",x"26160a",x"2c1a0c",x"2f1b0d",x"2d190b",x"2e1a0c",x"311c0d",x"321d0d",x"321d0d",x"321d0d",x"321d0e",x"321d0e",x"311d0d",x"2e1b0c",x"2e1b0c",x"2f1b0d",x"2d1a0c",x"2c190c",x"2a190b",x"2a190b",x"29180b",x"28180b",x"28180b",x"28170b",x"27170a",x"25150a",x"25150a",x"25160a",x"24150a",x"241509",x"231509",x"23150a",x"25160a",x"26160a",x"2a190b",x"2e1b0d",x"311d0d",x"331e0e",x"311c0d",x"301c0d",x"321d0d",x"321c0d",x"311c0d",x"311c0d",x"321d0d",x"331e0e",x"2d190b",x"2c190b",x"2b180a",x"2a170a",x"271509",x"251409",x"231308",x"271609",x"231408",x"211208",x"201208",x"211208",x"221309",x"211309",x"231409",x"231409",x"25150a",x"27170a",x"27160a",x"27160a",x"27160a",x"29170a",x"28170a",x"29170a",x"28160a",x"26160a",x"221409",x"1e1208",x"191008",x"160e07",x"191008",x"221409",x"26150a",x"26150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"6c6763",x"5c5a59",x"373432",x"373432",x"383432",x"373331",x"616060",x"616161",x"565555",x"393737",x"353433",x"333332",x"5b5b5b",x"585858",x"5d5d5d",x"4c4c4c",x"4a4a4a",x"424242",x"414141",x"454545",x"323232",x"323232",x"363636",x"494949",x"505050",x"575757",x"333333",x"333333",x"333333",x"000000",x"575757",x"565656",x"383838",x"313131",x"323232",x"434343",x"4b4b4b",x"4e4e4e",x"545454",x"4b4b4b",x"4a4a4a",x"343434",x"333333",x"35312f",x"352e2c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4a4a",x"494949",x"494949",x"474747",x"454545",x"4c4c4c",x"3a3a3a",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d160f",x"1d160f",x"1d160f",x"1c150e",x"1d160f",x"1b140d",x"1c150f",x"19120b",x"19130c",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"52483e",x"4c3f33",x"45382c",x"3e3126",x"413326",x"3f3024",x"433325",x"443326",x"463629",x"453528",x"4a3829",x"47372a",x"433227",x"443429",x"4a3a2e",x"4c3b2e",x"49392d",x"4a392d",x"4d3d31",x"504034",x"534337",x"58473a",x"574639",x"544033",x"533f31",x"543f30",x"543e2e",x"543e2d",x"533f30",x"4f3c2d",x"4a382a",x"4a3729",x"473427",x"473426",x"473426",x"493527",x"4a3728",x"4e3829",x"4c3728",x"4d382a",x"4c3829",x"4a3526",x"4c3829",x"4d3829",x"513d2c",x"523d2d",x"523c2d",x"4e3a2a",x"4f3b2e",x"4f3b2d",x"4e3b2c",x"4f3c2e",x"523e30",x"523d2d",x"533f2f",x"503a2b",x"4e392a",x"503a2b",x"503928",x"503a29",x"513a2b",x"4e3828",x"4d392b",x"4f3c2f",x"4e3b2d",x"4c3b2e",x"4d3b2e",x"4d3a2c",x"4b3829",x"4b3729",x"4c382a",x"4a3628",x"4b3728",x"4a3729",x"473528",x"483527",x"413125",x"3f2f22",x"3f3025",x"413125",x"3e2e24",x"3f3125",x"3b2d22",x"3e3126",x"3d3026",x"3c2e24",x"3a2e25",x"382d24",x"342a22",x"362b22",x"372c22",x"3c2f25",x"493f36",x"564b41",x"594f45",x"594f45",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"333333",x"333434",x"3a3736",x"36322f",x"3b3633",x"3b3532",x"3f3631",x"403933",x"3f3832",x"3f3630",x"443a33",x"423932",x"463c35",x"564e48",x"59534e",x"4b4b4b",x"525252",x"5b5a5a",x"5a5a5a",x"494949",x"4d4d4d",x"4d4d4d",x"4d4d4d",x"575757",x"5b5b5b",x"545454",x"4b433f",x"363636",x"323232",x"323232",x"313131",x"59504a",x"594f47",x"564b43",x"53473f",x"584d46",x"4c4440",x"635c58",x"4c4541",x"403731",x"413730",x"3e3733",x"3e3834",x"413831",x"413832",x"403831",x"423831",x"3c3530",x"3c3531",x"3d3631",x"333333",x"333333",x"323232",x"000000",x"000000",x"444342",x"444342",x"373433",x"333232",x"333333",x"353432",x"343332",x"000000",x"000000",x"353535",x"353535",x"343434",x"312f2c",x"333333",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"3d3d3d",x"383838",x"333333",x"313131",x"333333",x"303030",x"343434",x"333333",x"313131",x"323232",x"313131",x"5f5f5f",x"636363",x"424242",x"313131",x"323232",x"323232",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"28170a",x"28170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"28160a",x"4c3425",x"5f422f",x"593d2c",x"513828",x"573a27",x"4f3727",x"50392b",x"4e311e",x"4e311e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"291a09",x"291a09",x"291a09",x"211508",x"1f1308",x"27170b",x"2b190c",x"2a180b",x"26160a",x"1e1209",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"191008",x"1a1008",x"191008",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1f1408",x"150e07",x"150e07",x"150e07",x"160e07",x"1a1108",x"1f1209",x"231509",x"231409",x"231409",x"221409",x"211309",x"1e1208",x"1a1008",x"170f07",x"160e07",x"1c1108",x"251509",x"201208",x"211208",x"221309",x"211309",x"231409",x"231409",x"25150a",x"27160a",x"27160a",x"27160a",x"27160a",x"29170a",x"28170a",x"29170a",x"28160a",x"26160a",x"221409",x"1e1208",x"191008",x"160e07",x"191008",x"231409",x"27160a",x"27160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5f5d5c",x"555453",x"575655",x"535252",x"373433",x"373432",x"373534",x"474545",x"3f3d3c",x"3e3d3d",x"515151",x"565656",x"5d5d5d",x"585858",x"4d4d4d",x"4a4a4a",x"4c4c4c",x"3f3f3f",x"333333",x"383838",x"353535",x"333333",x"616160",x"595959",x"535353",x"595959",x"3c3c3c",x"323232",x"323232",x"000000",x"525251",x"575757",x"505050",x"3f3f3f",x"333333",x"414141",x"535353",x"4a4a4a",x"343434",x"545454",x"525252",x"4d4d4d",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1c150f",x"1d1610",x"1c160f",x"1c150e",x"1b140e",x"19120b",x"19120b",x"171009",x"171009",x"150e07",x"150e07",x"170f07",x"180f07",x"1b1108",x"1b1108",x"1a1108",x"191008",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1c1208",x"1d1208",x"1e1209",x"1f1309",x"201309",x"1f1208",x"1d1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"180f07",x"170f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181009",x"1b140c",x"1d150b",x"1d150c",x"1c130a",x"1d1308",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f08",x"191008",x"1b1008",x"1c1108",x"1d1108",x"1e1209",x"1f1309",x"211409",x"211409",x"221409",x"23150a",x"22140a",x"23150a",x"201309",x"201409",x"1f1209",x"1f1209",x"201309",x"1f1309",x"1f1309",x"1d1108",x"1f1309",x"1e1309",x"1d1208",x"1d1209",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1209",x"1d1209",x"1d1208",x"1e1208",x"1e1209",x"1e1309",x"1e1209",x"1e1209",x"1d1209",x"1b1108",x"1a1008",x"180f08",x"170f07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d190a",x"2f1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c2c2c",x"323232",x"333333",x"343434",x"343434",x"333333",x"333333",x"3a3430",x"3d3632",x"3d3631",x"3e3732",x"3d3631",x"3e3733",x"3d352e",x"413831",x"423831",x"554e4a",x"5b5654",x"5d5a58",x"625c58",x"585553",x"585453",x"5b5856",x"4d4d4d",x"4f4f4f",x"585858",x"605b59",x"5c5856",x"5d5955",x"4f4741",x"4c433d",x"483d36",x"564e4a",x"4b4038",x"473a31",x"4b3c32",x"493b31",x"473a30",x"463b32",x"433830",x"433932",x"413832",x"413831",x"403832",x"3f3833",x"413933",x"403732",x"403732",x"403832",x"5c5c5c",x"565656",x"4a4a4a",x"343434",x"323232",x"333333",x"303030",x"000000",x"4d4b4a",x"4d4b4a",x"343433",x"33302e",x"343332",x"343333",x"343333",x"000000",x"000000",x"505050",x"505050",x"424242",x"323232",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"383838",x"333333",x"333333",x"343434",x"333333",x"343434",x"342e2b",x"34302e",x"323232",x"343434",x"333333",x"313131",x"333333",x"363636",x"333333",x"343434",x"333333",x"323232",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f4f4f",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2a180b",x"2a180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"3d2513",x"5c3f2c",x"563927",x"583c29",x"543824",x"4d3424",x"4b3426",x"4b2f1d",x"4b2f1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a1b09",x"2a1b09",x"221508",x"1f1308",x"231509",x"27170a",x"27160a",x"24150a",x"1e1209",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"180f08",x"1a1008",x"1b1108",x"1a1008",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181007",x"1e1308",x"150e07",x"150e07",x"150e07",x"160e07",x"190f07",x"201309",x"25160a",x"26160a",x"26160a",x"241509",x"211309",x"1f1208",x"1b1108",x"180f07",x"160e07",x"1e1208",x"27160a",x"27160a",x"211208",x"221309",x"211309",x"231409",x"231409",x"25150a",x"27160a",x"27160a",x"27160a",x"27160a",x"29170a",x"28170a",x"29170a",x"28160a",x"26160a",x"221409",x"1e1208",x"191008",x"160e07",x"191008",x"231409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"575655",x"5c5b59",x"636261",x"666564",x"494848",x"454443",x"474545",x"4a4948",x"565656",x"616161",x"515151",x"595959",x"575757",x"4e4e4e",x"3f3f3f",x"343434",x"333333",x"333333",x"373737",x"363635",x"000000",x"646464",x"606060",x"484848",x"4b4b4b",x"363636",x"323232",x"323232",x"000000",x"51504e",x"575654",x"5c5c5c",x"515151",x"595959",x"4b4b4b",x"474747",x"323232",x"313131",x"5f5e5e",x"595959",x"363636",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1711",x"1d1711",x"1e1711",x"1c150e",x"1c150f",x"1c160f",x"1b150e",x"1b150e",x"1a130c",x"17110a",x"17110a",x"150e07",x"170f07",x"170f07",x"180f07",x"1b1108",x"1b1108",x"1a1108",x"191008",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"170f07",x"180f07",x"191008",x"1a1008",x"1c1208",x"1d1208",x"1e1209",x"1f1309",x"201309",x"1f1208",x"1d1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"180f07",x"170f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181009",x"1b140c",x"1d150b",x"1d150c",x"1c130a",x"1d1308",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f08",x"191008",x"1b1008",x"1c1108",x"1d1108",x"1e1209",x"1f1309",x"211409",x"211409",x"221409",x"23150a",x"22140a",x"23150a",x"201309",x"201409",x"1f1209",x"1f1209",x"201309",x"1f1309",x"1f1309",x"1d1108",x"1f1309",x"1e1309",x"1d1208",x"1d1209",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1209",x"1d1209",x"1d1208",x"1e1208",x"1e1209",x"1e1309",x"1e1209",x"1e1209",x"1d1209",x"1b1108",x"1a1008",x"180f08",x"170f07",x"160e07",x"160e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d190a",x"2f1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"303131",x"313131",x"333333",x"343434",x"323232",x"313131",x"333333",x"313131",x"323232",x"3b3430",x"38302b",x"3e3632",x"3c3531",x"3f362f",x"413831",x"413831",x"403832",x"3b3531",x"433e3a",x"5b5755",x"686564",x"5f5d5c",x"666361",x"605d5b",x"5b5856",x"635f5d",x"625e5c",x"4d4946",x"413b36",x"403832",x"453931",x"413832",x"443a32",x"463a31",x"473a31",x"493b31",x"493b32",x"473b32",x"473c34",x"443a33",x"514943",x"3e3732",x"413831",x"3e3732",x"403731",x"3e3732",x"414141",x"555555",x"484848",x"606060",x"333333",x"303030",x"313131",x"292929",x"2d2d2d",x"323232",x"000000",x"4f4f4f",x"4f4f4f",x"343434",x"373533",x"302f2f",x"323131",x"323131",x"000000",x"000000",x"000000",x"585858",x"4f4f4f",x"323232",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"343434",x"333333",x"33312f",x"323130",x"343333",x"333130",x"333231",x"323232",x"333130",x"343434",x"353535",x"323232",x"333333",x"333333",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"636363",x"323232",x"4b4b4b",x"4f4f4f",x"6c6a68",x"000000",x"000000",x"000000"),
(x"000000",x"2f1a0b",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"4a3222",x"5b3f2c",x"5d3f2a",x"563925",x"4d3323",x"4c3323",x"483123",x"52331d",x"52331d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c1b09",x"2c1b09",x"231608",x"211409",x"231509",x"27170a",x"26150a",x"26160a",x"1d1208",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"191008",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181007",x"1e1308",x"150e07",x"150e07",x"150e07",x"170f07",x"1c1108",x"221409",x"251509",x"28170a",x"28170a",x"26160a",x"221409",x"201309",x"1c1108",x"180f07",x"160e07",x"1e1208",x"27160a",x"27160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e5d5b",x"656362",x"595756",x"666564",x"565452",x"5d5b5a",x"595858",x"515050",x"464545",x"3e3d3d",x"353535",x"3c3c3c",x"424242",x"3b3b3b",x"343434",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"60605f",x"5b5b5b",x"3e3e3e",x"323232",x"333333",x"333333",x"000000",x"606060",x"575757",x"504f4f",x"525252",x"484848",x"343434",x"323232",x"323232",x"323232",x"5d5d5d",x"4c4c4c",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1710",x"1d1710",x"1d1610",x"1c160f",x"1d160f",x"1d1610",x"1c150e",x"1c150e",x"19120c",x"19120b",x"18110a",x"160f07",x"170f07",x"170f07",x"170f07",x"180f08",x"191008",x"180f08",x"180f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"191008",x"1a1008",x"1b1108",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1108",x"1a1008",x"191008",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"18110a",x"1a120b",x"1c140c",x"1a120b",x"20150a",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"180f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1c1108",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"1a1008",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"191008",x"1a1008",x"1a1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f08",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"1c1108",x"1c1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"303030",x"2c2c2c",x"303030",x"333333",x"313131",x"313131",x"323232",x"333333",x"363433",x"373331",x"393431",x"3f3731",x"403731",x"413730",x"413831",x"403833",x"3c3531",x"3e3733",x"393532",x"3a3633",x"33312f",x"3a3532",x"3b3735",x"3e3631",x"3a3634",x"3a3431",x"3a3633",x"423a34",x"3a3531",x"423932",x"423830",x"453a32",x"463a32",x"473a31",x"473a31",x"483c33",x"453a32",x"453a33",x"423831",x"514a45",x"3d3633",x"423831",x"3d3632",x"494949",x"4c4a4a",x"414141",x"343434",x"323232",x"333333",x"313131",x"323232",x"323232",x"313131",x"333333",x"333333",x"000000",x"4b4b4b",x"464646",x"333333",x"2f2f2f",x"303030",x"323232",x"323232",x"000000",x"000000",x"4f4f4f",x"4f4f4f",x"4e4e4e",x"333333",x"303030",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333131",x"333131",x"323232",x"3c3c3c",x"3b3b3b",x"414141",x"474747",x"515151",x"5b5b5b",x"666666",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"525252",x"4f4f4f",x"4e4e4e",x"636363",x"434343",x"353535",x"6c6a68",x"353535",x"323232",x"000000",x"000000"),
(x"000000",x"29170a",x"29170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"49301f",x"60412b",x"593c28",x"513523",x"543926",x"543826",x"483224",x"52321d",x"52321d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d1c0a",x"2d1c0a",x"221508",x"211509",x"201309",x"25150a",x"26160a",x"231409",x"1c1108",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f08",x"1c1108",x"1d1108",x"201309",x"1f1309",x"1d1108",x"191008",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f08",x"190f08",x"180f08",x"190f07",x"1c1107",x"1e1308",x"170f07",x"170f07",x"180f07",x"1a1008",x"1d1108",x"231409",x"261509",x"261509",x"251509",x"231409",x"211309",x"1e1108",x"1a1008",x"170f07",x"160e07",x"1b1008",x"231308",x"231308",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595756",x"5a5858",x"565452",x"5d5b5a",x"595858",x"515050",x"464545",x"3e3d3d",x"323131",x"3c3c3c",x"414141",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"60605f",x"555555",x"3e3e3e",x"353535",x"333333",x"000000",x"000000",x"000000",x"5b5b5b",x"545454",x"393939",x"342d2a",x"333333",x"333333",x"323232",x"323232",x"000000",x"4c4c4c",x"323232",x"333232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d160f",x"1d160f",x"1d160f",x"1d1610",x"1d1711",x"1d1710",x"1d160f",x"1b150e",x"1c150e",x"19120c",x"19110a",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"180f07",x"190f08",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"181009",x"1a130c",x"18110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"180f07",x"190f07",x"1a1008",x"1b1108",x"1b1108",x"1b1008",x"1c1108",x"1c1108",x"1b1108",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"191008",x"1a1008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"190f08",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"190f08",x"190f07",x"191008",x"191008",x"180f07",x"180f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"241409",x"241409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"303030",x"2e2e2e",x"323232",x"323232",x"343434",x"343434",x"313131",x"323131",x"333231",x"373432",x"3d3632",x"3d352f",x"433f3c",x"55514e",x"3f3732",x"3f3935",x"47413d",x"4b4744",x"524f4d",x"51504e",x"4d4a48",x"423f3e",x"484340",x"464340",x"413e3d",x"484340",x"413d3b",x"3e3732",x"3b3531",x"3e3834",x"443a33",x"453930",x"443931",x"483b31",x"473a31",x"473b31",x"453a31",x"453a32",x"423831",x"515151",x"3d3d3d",x"424242",x"474747",x"383838",x"323232",x"333333",x"303030",x"323232",x"313131",x"313131",x"333333",x"323232",x"323232",x"333333",x"333333",x"000000",x"434343",x"434343",x"323232",x"313131",x"323232",x"313131",x"313131",x"000000",x"000000",x"4f4f4f",x"4f4f4f",x"4e4e4e",x"343434",x"323232",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"353535",x"2f2f2f",x"535353",x"494949",x"545454",x"5a5a5a",x"666666",x"696969",x"5f5f5f",x"333333",x"313131",x"323232",x"4f4f4f",x"474747",x"565656",x"5d5d5d",x"4f4f4f",x"464646",x"313131",x"332f2c",x"313131",x"323232",x"323232",x"000000",x"000000"),
(x"000000",x"261609",x"261609",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"4e3321",x"5a3e2a",x"5b3e28",x"563a26",x"543825",x"503423",x"473124",x"51321d",x"51321d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b1b0a",x"2b1b0a",x"221508",x"1f1308",x"221409",x"2b180b",x"2b190b",x"2d1a0c",x"2f1c0d",x"2a180b",x"2e1b0c",x"311d0d",x"2f1b0d",x"321d0d",x"351f0e",x"341e0e",x"37200f",x"3a2210",x"39210f",x"351e0e",x"311c0d",x"331c0d",x"361e0d",x"371f0e",x"351e0d",x"351e0d",x"331d0d",x"2d1a0c",x"341d0d",x"321c0c",x"331c0c",x"38200f",x"3b2210",x"36200f",x"38200f",x"38200e",x"361f0e",x"351e0d",x"321c0c",x"331c0c",x"351d0d",x"361e0d",x"38200e",x"38200f",x"39200f",x"3a210f",x"361f0e",x"351e0d",x"39200f",x"38200e",x"361f0e",x"341d0d",x"38200e",x"38200e",x"37200d",x"341d0c",x"2e1a0b",x"2c180a",x"2d190a",x"2b180a",x"2a170a",x"2e190b",x"331c0c",x"2e1a0b",x"321c0c",x"311c0c",x"2f1b0c",x"2d190b",x"231509",x"1c1108",x"160e07",x"1d1108",x"251509",x"251509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"333333",x"434242",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"313131",x"323232",x"363636",x"3d3d3d",x"393939",x"342d2a",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"393939",x"3f3f3f",x"404040",x"5b5b5b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c160f",x"1c160f",x"1d1710",x"1d1610",x"1c160f",x"1d1710",x"1d160f",x"1a140d",x"1b150e",x"19130c",x"1a120b",x"191109",x"180f08",x"191008",x"191008",x"191008",x"191008",x"180f08",x"180f07",x"180f08",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1008",x"1d1208",x"1e1209",x"1e1209",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"1a1008",x"180f08",x"170f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"191008",x"191008",x"190f07",x"190f07",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"1a1008",x"191008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1208",x"1c1108",x"1b1108",x"1a1008",x"191008",x"191008",x"170f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"25150a",x"25150a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e2e2e",x"313131",x"333333",x"333333",x"333333",x"333333",x"323131",x"343333",x"373432",x"3c3734",x"393431",x"3b3531",x"3c3734",x"3b3531",x"373331",x"585553",x"3b3531",x"3d3531",x"484543",x"4f4b49",x"433f3c",x"474443",x"41403f",x"4c4a48",x"474443",x"44403e",x"403d3c",x"3d3733",x"3b3530",x"3e3733",x"433932",x"453930",x"433932",x"483b31",x"525252",x"585858",x"5c5c5c",x"585858",x"515151",x"535353",x"393939",x"333333",x"333333",x"313131",x"333333",x"303030",x"313131",x"323232",x"333333",x"323232",x"4f4f4f",x"323232",x"333333",x"000000",x"000000",x"000000",x"3f3f3f",x"3f3f3f",x"303030",x"323232",x"323232",x"313131",x"313131",x"000000",x"000000",x"515050",x"515050",x"515050",x"323232",x"313131",x"282828",x"282828",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"333333",x"323232",x"313131",x"323232",x"323232",x"323232",x"343434",x"333333",x"5f5f5f",x"333333",x"313131",x"313131",x"323232",x"474747",x"313131",x"313131",x"313131",x"323232",x"323232",x"333232",x"323232",x"494949",x"323232",x"000000",x"000000"),
(x"000000",x"2a170a",x"2a170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"4a3121",x"573f2c",x"523926",x"513423",x"553725",x"513625",x"473124",x"50321d",x"50321d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c1b0a",x"2c1b0a",x"221508",x"211509",x"26160a",x"29180b",x"27170b",x"29170a",x"2b190b",x"2a180b",x"2e1a0c",x"341f0e",x"2e1a0b",x"321c0c",x"38210f",x"38210f",x"39210f",x"38200f",x"38200f",x"3c220f",x"381f0e",x"371f0e",x"38200e",x"39200f",x"38200f",x"371f0e",x"371f0f",x"38200f",x"3a200f",x"361f0e",x"38200f",x"351e0d",x"351e0d",x"38200f",x"331d0d",x"351e0e",x"351e0e",x"38200f",x"37200e",x"351e0d",x"341d0d",x"351d0d",x"361e0d",x"39200f",x"3e2511",x"3f2511",x"3c2210",x"39200f",x"3a200e",x"3c220f",x"3b2210",x"3b210f",x"3b220f",x"3b230f",x"3a210f",x"38200e",x"321c0c",x"321c0c",x"331c0c",x"2f1a0b",x"2e190b",x"311b0b",x"321c0c",x"341d0d",x"331d0d",x"361f0e",x"311c0d",x"2d1a0b",x"26160a",x"1b1108",x"160e07",x"1d1108",x"27170a",x"27170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"323232",x"323232",x"3a3a3a",x"434343",x"313131",x"333333",x"333333",x"353535",x"4b4b4b",x"575757",x"424242",x"3c3c3c",x"404040",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"313131",x"323232",x"363636",x"3d3d3d",x"3c3c3c",x"434343",x"4f4d4d",x"5c5c5c",x"000000",x"000000",x"000000",x"343434",x"494949",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"313131",x"393939",x"3f3f3f",x"4a4a4a",x"595959",x"515151",x"494949",x"000000",x"000000",x"000000",x"000000",x"301b0b",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1610",x"1d1610",x"1d1610",x"1d1710",x"1d1710",x"1d160f",x"1d1610",x"1c150e",x"1b150e",x"19130c",x"1a130b",x"191109",x"180f07",x"180f07",x"191008",x"191008",x"191008",x"180f07",x"180f07",x"180f08",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"170f07",x"170f07",x"191008",x"191008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1a1008",x"190f08",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f08",x"191008",x"190f08",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"191008",x"191008",x"190f08",x"191008",x"180f07",x"191008",x"190f08",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"1c1108",x"1a1008",x"190f08",x"191008",x"191008",x"180f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"2a190a",x"29180a",x"29180a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"333333",x"333232",x"333332",x"353332",x"3c342e",x"3b3531",x"373533",x"3a3633",x"443a32",x"3b3632",x"393533",x"3f3732",x"3b3531",x"3b3531",x"393431",x"373432",x"393532",x"383331",x"474341",x"413d3b",x"46433f",x"545150",x"524f4d",x"5d5a59",x"5d5b5a",x"605e5d",x"595959",x"5b5b5b",x"5a5a5a",x"525252",x"585858",x"5c5c5c",x"575757",x"474747",x"292929",x"272727",x"323232",x"313131",x"313131",x"333333",x"343434",x"323232",x"313131",x"313131",x"313131",x"383838",x"000000",x"000000",x"000000",x"000000",x"000000",x"444444",x"444444",x"323232",x"313131",x"323232",x"333231",x"333231",x"000000",x"000000",x"4c4b4b",x"4c4b4b",x"484747",x"302f2f",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"333333",x"313131",x"323232",x"323232",x"323232",x"323232",x"323232",x"343434",x"323232",x"323232",x"333333",x"333333",x"323232",x"343434",x"313131",x"323232",x"484848",x"373736",x"323131",x"323232",x"323232",x"505050",x"000000",x"000000",x"000000"),
(x"000000",x"2c180a",x"2c180a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"26150a",x"41291a",x"583d2a",x"523a27",x"4e3624",x"543623",x"533624",x"452e20",x"51321c",x"51321c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1d0b",x"2f1d0b",x"251709",x"2c1b0c",x"2c190b",x"321d0d",x"331d0d",x"341d0d",x"331d0d",x"371f0e",x"37200e",x"371f0e",x"3a210f",x"3b2310",x"3f2511",x"3b2210",x"3e2310",x"3d230f",x"402511",x"402511",x"3e2410",x"412612",x"3f2511",x"3c220f",x"402411",x"3b210f",x"3c210f",x"3d2310",x"3b2210",x"402511",x"3e2311",x"3c220f",x"3c220f",x"3f2612",x"3a2210",x"402512",x"3f2411",x"402511",x"432713",x"422713",x"452914",x"412612",x"3e2410",x"3e2310",x"3e2410",x"402511",x"3d2310",x"3f2410",x"3f2410",x"3e2310",x"402511",x"3e2310",x"432712",x"402512",x"3e2410",x"381f0d",x"331c0c",x"351d0d",x"38200e",x"3a210f",x"3a200e",x"351e0d",x"381f0e",x"381f0e",x"38200f",x"371f0e",x"371f0e",x"341d0d",x"321c0d",x"27170a",x"201309",x"1f1309",x"29180b",x"29180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"323232",x"323232",x"323232",x"3a3a3a",x"434343",x"313232",x"333333",x"404040",x"4b4b4b",x"3b3b3b",x"555555",x"424242",x"3c3c3c",x"404040",x"3c3b3b",x"393939",x"414141",x"4b4b4b",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"333333",x"3d3d3d",x"414141",x"515151",x"585858",x"656565",x"626262",x"4f5050",x"504f4f",x"5e5e5e",x"595858",x"5b5b5b",x"323232",x"343434",x"494949",x"5a5a5a",x"5c5c5c",x"343434",x"3b3b3b",x"000000",x"000000",x"000000",x"313232",x"323232",x"323232",x"343434",x"535353",x"555555",x"595959",x"5a5a5a",x"565656",x"494949",x"515151",x"565656",x"000000",x"000000",x"301b0b",x"301b0b",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1710",x"1d160f",x"1d160f",x"1d160f",x"1d160f",x"1d1710",x"1c150e",x"1b150e",x"1b140d",x"1a130b",x"191109",x"180f07",x"180f08",x"191008",x"191008",x"191008",x"190f08",x"180f08",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160f07",x"170f07",x"170f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"160f07",x"170f07",x"180f08",x"191008",x"1a1008",x"1c1108",x"1d1209",x"1e1209",x"1f1309",x"1f1309",x"1e1209",x"1e1209",x"1d1209",x"1c1108",x"1b1108",x"1a1008",x"180f08",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"180f07",x"180f08",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"1b1108",x"1b1108",x"1a1008",x"190f07",x"180f07",x"180f07",x"190f07",x"191008",x"191008",x"191008",x"191008",x"190f08",x"191008",x"180f08",x"180f08",x"180f08",x"190f08",x"180f08",x"191008",x"191008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"231608",x"331e0d",x"321d0c",x"321d0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"343333",x"363432",x"383431",x"3d3630",x"393532",x"3d3733",x"3d3733",x"3e3631",x"3c3632",x"39332f",x"3c3531",x"3c3633",x"383431",x"383533",x"383432",x"3a3633",x"393431",x"3c3531",x"3b3531",x"37322f",x"363432",x"56524f",x"646160",x"605e5d",x"616161",x"656362",x"5d5d5d",x"605e5d",x"535353",x"3a3a3a",x"343434",x"323232",x"333333",x"313131",x"323232",x"333333",x"323232",x"313131",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"444444",x"444444",x"313131",x"323232",x"323232",x"343230",x"343230",x"000000",x"000000",x"4d4b4a",x"4d4b4a",x"42403f",x"353332",x"333232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"323232",x"323232",x"333333",x"313131",x"333333",x"333333",x"323232",x"333333",x"333333",x"313132",x"343434",x"343434",x"323232",x"414140",x"3d3d3d",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"261509",x"261509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"4f3524",x"593e2c",x"5a3e29",x"4b3423",x"573924",x"503523",x"412b1e",x"50311b",x"50311b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"35210b",x"35210b",x"281909",x"211509",x"1e1209",x"23150a",x"27170b",x"24150a",x"24150a",x"231509",x"25160a",x"2c1a0c",x"2c1a0c",x"2e1a0c",x"2d1a0b",x"321c0c",x"321c0c",x"331d0d",x"361e0d",x"361f0e",x"38200e",x"38200e",x"361e0e",x"371f0e",x"38200f",x"3a2210",x"351e0e",x"311c0c",x"321c0d",x"321d0d",x"341e0e",x"331d0e",x"36200f",x"36200f",x"321d0d",x"2d1a0b",x"2d190b",x"2f1a0c",x"301b0c",x"331d0d",x"37200e",x"39210f",x"3a220f",x"371f0e",x"371f0e",x"361e0d",x"351e0d",x"381f0e",x"38200e",x"371f0e",x"381f0e",x"371f0e",x"39210e",x"361e0d",x"37200e",x"321d0d",x"2f1b0b",x"2c190b",x"2d1a0b",x"2c190b",x"2f1b0b",x"2c190b",x"2f1a0b",x"331e0e",x"301c0d",x"311c0d",x"2d190b",x"2a180b",x"24150a",x"1c1108",x"170f07",x"1d1108",x"28170a",x"28170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"313131",x"333333",x"323232",x"323232",x"353535",x"4b4b4b",x"494949",x"3c3c3c",x"333333",x"4a4a4a",x"464646",x"424242",x"3e3e3e",x"494949",x"595959",x"5e5e5e",x"494949",x"404040",x"454545",x"535353",x"5b5b5b",x"5d5d5d",x"000000",x"343434",x"323231",x"313131",x"323232",x"454545",x"515151",x"4c4c4c",x"474747",x"515151",x"313131",x"363636",x"323232",x"4b4b4b",x"464646",x"595959",x"4b4b4b",x"323232",x"353535",x"3a3a3a",x"575656",x"5b5b5b",x"343434",x"3b3b3b",x"575757",x"000000",x"000000",x"323333",x"323232",x"323232",x"3f3f3f",x"474747",x"3e3e3e",x"353535",x"313131",x"363636",x"474747",x"565656",x"5d5c5b",x"000000",x"000000",x"261609",x"261609",x"1e1208",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"191008",x"180f08",x"170f07",x"160f07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"1b1108",x"1d1208",x"1e1209",x"1e1209",x"1e1209",x"1e1208",x"1e1208",x"1d1208",x"1d1208",x"1d1108",x"1d1108",x"1d1208",x"1e1208",x"1d1108",x"1e1208",x"1e1209",x"1f1309",x"1e1208",x"1e1208",x"1e1209",x"201409",x"201309",x"211409",x"22150a",x"211409",x"201309",x"1f1208",x"1f1208",x"1f1209",x"201309",x"221409",x"231509",x"24150a",x"24150a",x"221409",x"211409",x"201309",x"201309",x"1f1208",x"1e1208",x"1c1108",x"1b1108",x"191008",x"180f08",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211508",x"1d130a",x"1d1409",x"1b1209",x"1f140b",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f07",x"180f07",x"190f07",x"190f07",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1c1108",x"1e1208",x"201308",x"1d1108",x"211309",x"201309",x"1f1208",x"1e1208",x"1e1209",x"1d1208",x"1b1108",x"1a1008",x"191008",x"180f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"180f08",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"160f07",x"150e07",x"150e07",x"1c1208",x"221508",x"2d1a0b",x"2e1b0b",x"2e1b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a3532",x"403732",x"373432",x"3d3733",x"3e352f",x"433b35",x"3b322b",x"3a3532",x"3a3633",x"3b3632",x"373331",x"3a3431",x"3a3532",x"393431",x"353230",x"3b3531",x"3a3430",x"3c3633",x"353231",x"383533",x"343231",x"373432",x"333232",x"333333",x"333333",x"323232",x"323232",x"323232",x"353535",x"303030",x"333333",x"323232",x"333333",x"343434",x"333333",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"474747",x"474747",x"35312d",x"262626",x"313131",x"2e2e2e",x"333333",x"000000",x"000000",x"575553",x"575553",x"484645",x"333130",x"333232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"333333",x"333333",x"323232",x"333333",x"333333",x"313132",x"343434",x"343434",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"26160a",x"26160a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251409",x"462d1d",x"553a28",x"583b28",x"513622",x"513523",x"503421",x"432e22",x"50311d",x"50311d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38291c",x"38291c",x"302317",x"281d14",x"2c1f15",x"2d1d13",x"2c1c12",x"2a1b10",x"2e1d11",x"2a1b10",x"311e11",x"342012",x"361f10",x"311d0f",x"341f10",x"351f0f",x"301c0e",x"321d0f",x"2d190d",x"311c0e",x"331c0f",x"351f10",x"361e0f",x"371f0f",x"361e0f",x"381f0f",x"362010",x"362010",x"372011",x"3a2211",x"371f10",x"3b2211",x"372010",x"3b2413",x"392313",x"392314",x"3a2414",x"382313",x"382113",x"382214",x"382212",x"372012",x"372011",x"392212",x"3d2514",x"3b2312",x"3b2110",x"392010",x"382010",x"381f0f",x"3a2110",x"3a2111",x"3a2110",x"371e0f",x"331c0e",x"311c0d",x"361f10",x"371f10",x"361e0f",x"321c0e",x"351f10",x"352011",x"351f10",x"341f12",x"301d11",x"362011",x"382213",x"362314",x"312013",x"231810",x"1d150e",x"25190f",x"312014",x"312014",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"313131",x"333333",x"3f3f3f",x"414141",x"424242",x"414141",x"414141",x"414141",x"464646",x"474747",x"3d3d3d",x"454545",x"4d4d4d",x"4c4c4c",x"4c4c4c",x"444444",x"464646",x"545454",x"595959",x"595959",x"5d5d5d",x"575656",x"545353",x"333333",x"343434",x"343434",x"646464",x"4b4b4a",x"585858",x"4c4c4c",x"424242",x"515151",x"313131",x"323333",x"323232",x"333333",x"303030",x"454545",x"494949",x"3f3e3d",x"313131",x"4d4d4d",x"454545",x"5a5a5a",x"333333",x"575757",x"5f5f5e",x"353535",x"434343",x"343434",x"333334",x"343434",x"3d3d3d",x"474747",x"595857",x"353535",x"333333",x"333333",x"323232",x"545454",x"565656",x"565656",x"000000",x"1a1107",x"1a1107",x"191107",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"180f08",x"1a1008",x"1a1008",x"191008",x"190f08",x"180f08",x"180f07",x"170f07",x"170f07",x"180f07",x"190f08",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"190f07",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201208",x"211309",x"211309",x"221409",x"221409",x"221409",x"23150a",x"23150a",x"221409",x"221409",x"211409",x"211309",x"221409",x"221409",x"221409",x"221409",x"231509",x"24150a",x"231509",x"221409",x"201309",x"1f1209",x"1e1208",x"1d1108",x"1b1108",x"191008",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"271809",x"231608",x"1c1108",x"191007",x"190f07",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f08",x"1a1008",x"1b1008",x"1d1108",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1d1208",x"1e1208",x"1d1108",x"1e1208",x"211309",x"1f1208",x"221409",x"211409",x"201309",x"1e1208",x"1d1208",x"1b1108",x"1a1008",x"1a1008",x"191008",x"191008",x"180f07",x"180f08",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f08",x"150e07",x"160e07",x"160e07",x"170f07",x"191007",x"160f07",x"170f07",x"160f07",x"160e07",x"231608",x"33200a",x"37210d",x"321e0c",x"321e0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e352f",x"433b35",x"39332f",x"3a3532",x"3a3633",x"3c3632",x"393431",x"38332f",x"3b3531",x"383432",x"393431",x"3b3633",x"383533",x"3a3634",x"373432",x"343231",x"3f3c3a",x"434241",x"3c3b3b",x"3d3a38",x"393939",x"454545",x"3f3f3f",x"3f3936",x"393939",x"323232",x"312f2e",x"323232",x"333333",x"343434",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d4d4d",x"4d4d4d",x"454442",x"323232",x"2e2f2f",x"313131",x"323232",x"000000",x"000000",x"000000",x"43413f",x"43413f",x"383534",x"343332",x"343434",x"343434",x"3b3b3b",x"434343",x"494949",x"3d3d3d",x"333333",x"000000",x"474747",x"383838",x"323232",x"323232",x"313131",x"323232",x"4b4b4b",x"4a4a4a",x"545454",x"4a4a4a",x"464646",x"373737",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2b180b",x"2b180b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"241409",x"4d3526",x"4d382a",x"5d402b",x"543724",x"573824",x"4c3222",x"3f2d22",x"4e301c",x"4e301c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"52453a",x"52453a",x"43362b",x"3a3026",x"3b322a",x"392f26",x"352b22",x"332921",x"32271f",x"332820",x"33281f",x"35281e",x"322419",x"352419",x"362519",x"3e2c20",x"412f21",x"412d20",x"412d21",x"412d1f",x"412d20",x"402c1f",x"3c2819",x"382315",x"352113",x"362418",x"38261a",x"342317",x"36251a",x"342215",x"342114",x"331f13",x"301f13",x"2e1d12",x"2f1f15",x"302117",x"2f2117",x"2f1f15",x"312217",x"372519",x"39271a",x"3c281b",x"3e2a1b",x"3a2719",x"372216",x"392415",x"382112",x"382211",x"3b2616",x"3a2517",x"3c2618",x"3b2618",x"3c2719",x"392618",x"362316",x"362316",x"362419",x"322318",x"312217",x"332318",x"34251a",x"352519",x"36261b",x"3a2a1f",x"3a2a1f",x"38271b",x"3b291d",x"38281c",x"34261c",x"2f261d",x"302820",x"342b23",x"40352b",x"40352b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"3f3f3f",x"434343",x"3e3e3e",x"454545",x"383838",x"373737",x"3e3e3e",x"434343",x"454545",x"4d4d4d",x"474747",x"404040",x"343434",x"333333",x"3d3d3d",x"363636",x"333333",x"313131",x"444444",x"464646",x"545353",x"585858",x"323232",x"313131",x"5d5d5d",x"51504e",x"4f4f4f",x"4b4b4a",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"333333",x"353636",x"434343",x"3f3f3f",x"323232",x"3d3d3d",x"464646",x"454545",x"424242",x"4d4d4d",x"484848",x"353535",x"434343",x"363636",x"313131",x"545454",x"414141",x"474747",x"4c4c4b",x"595756",x"333333",x"323232",x"323333",x"4a4a4a",x"5d5c5a",x"5d5c5a",x"000000",x"181007",x"181007",x"1c1208",x"1d1308",x"181007",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"170f07",x"160e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"241708",x"201408",x"1b1108",x"1f1309",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"191008",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1d1208",x"1e1209",x"1e1208",x"1e1208",x"1f1209",x"1f1309",x"201309",x"211409",x"201309",x"221409",x"221409",x"231409",x"24150a",x"231509",x"231409",x"231409",x"231409",x"221409",x"231409",x"241509",x"24150a",x"231409",x"211309",x"201208",x"201208",x"1f1208",x"201309",x"211309",x"231409",x"24150a",x"241509",x"26160a",x"27170a",x"241509",x"231409",x"241509",x"24150a",x"231409",x"211409",x"201309",x"1f1209",x"1d1208",x"1b1108",x"190f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1e0a",x"311f0a",x"2c1c09",x"261809",x"1d1308",x"1b1107",x"180f07",x"180f07",x"180f08",x"180f08",x"191008",x"1c1108",x"1d1108",x"1f1208",x"1d1108",x"1f1208",x"1e1208",x"1d1108",x"1c1108",x"1c1108",x"1e1208",x"201208",x"1d1108",x"211309",x"1e1108",x"23150a",x"221409",x"201309",x"1f1309",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1108",x"1a1008",x"150e07",x"150e07",x"170f07",x"170f07",x"181007",x"180f07",x"180f07",x"180f07",x"170f07",x"291a09",x"311f0b",x"3b240c",x"3a230d",x"3a230d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"393431",x"3a3431",x"3b3531",x"393532",x"393432",x"393533",x"3a3533",x"373432",x"363331",x"353332",x"3c3a39",x"3d3a39",x"3a322c",x"404040",x"3a3a3a",x"454545",x"434343",x"3f3936",x"3a3a3a",x"353535",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"575757",x"575757",x"464443",x"333232",x"333332",x"323232",x"333232",x"333232",x"000000",x"000000",x"3f3c3a",x"3f3c3a",x"363433",x"333232",x"333232",x"333232",x"3b3b3b",x"434343",x"494949",x"333333",x"333333",x"525252",x"474747",x"383838",x"323232",x"323232",x"313131",x"323232",x"4b4b4b",x"4a4a4a",x"545454",x"4b4b4b",x"464646",x"373737",x"5c5c5c",x"5c5c5c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"331c0c",x"331c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"4d3829",x"503b2e",x"664630",x"573c28",x"5c3d29",x"4f3422",x"412f24",x"4b2e1a",x"4b2e1a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"51463a",x"51463a",x"42382e",x"3d332a",x"352c24",x"362c24",x"33291f",x"30261e",x"32271f",x"342921",x"362b22",x"3a2d24",x"38291f",x"39291f",x"3b2a1e",x"412f24",x"443225",x"433123",x"412e21",x"412c1e",x"402c1f",x"412c1d",x"432f22",x"453121",x"3b281b",x"3e2c1f",x"38271b",x"38261a",x"352316",x"372418",x"342114",x"332014",x"321f13",x"331f12",x"322014",x"332216",x"301f14",x"312116",x"322015",x"362316",x"382416",x"3a2516",x"3c2717",x"3c2719",x"3b2516",x"3b2415",x"3c2618",x"3d271a",x"3e2b1d",x"402c1f",x"412e21",x"3d2b1e",x"3e2a1d",x"3f2b1d",x"3a281c",x"3e2b1d",x"39291e",x"39291d",x"38291e",x"36281e",x"37291f",x"3c2e24",x"392a20",x"3a2b21",x"39291f",x"38271c",x"3a2a1e",x"37261a",x"36281e",x"332820",x"3e352d",x"4e433a",x"52473c",x"52473c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"3b3b3b",x"333333",x"333333",x"313131",x"3f3f3f",x"474747",x"4b4b4b",x"494949",x"484848",x"474747",x"414141",x"393939",x"323232",x"333333",x"333333",x"3d3d3d",x"323232",x"333333",x"333333",x"323232",x"474747",x"444444",x"545454",x"333333",x"323232",x"464646",x"585756",x"585756",x"323232",x"393837",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"323232",x"323232",x"4a4a4a",x"373737",x"434343",x"3e3e3e",x"3c3c3c",x"3d3d3d",x"3e3e3e",x"3a3b3b",x"4b4b4b",x"555555",x"484848",x"393939",x"343434",x"363636",x"434343",x"494949",x"505050",x"555453",x"555453",x"323232",x"323232",x"303030",x"4f4e4d",x"55524f",x"000000",x"1c1208",x"1c1208",x"201508",x"211508",x"241708",x"160e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"190f07",x"180f07",x"150e07",x"150e07",x"150e07",x"170f07",x"191007",x"1d1308",x"211508",x"331f0b",x"271809",x"271809",x"251709",x"1e1208",x"1d1208",x"1c1108",x"1c1108",x"1b1108",x"1a1108",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"201309",x"211409",x"221409",x"231509",x"25160a",x"241509",x"27170b",x"26160a",x"26160a",x"25150a",x"25160a",x"231409",x"241509",x"241509",x"25160a",x"241509",x"221409",x"221409",x"231509",x"221409",x"221409",x"211409",x"221409",x"24150a",x"25160a",x"26160a",x"27160a",x"27170a",x"26160a",x"26160a",x"25150a",x"231409",x"221409",x"211309",x"201309",x"1f1208",x"1d1108",x"1c1108",x"1a1008",x"180f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"171007",x"251708",x"21150b",x"1d1308",x"1f1309",x"1a1008",x"1c1108",x"1b1108",x"1c1108",x"1d1108",x"1d1208",x"1f1208",x"1e1208",x"201308",x"1f1208",x"201309",x"1e1208",x"1b1008",x"1b1008",x"1b1008",x"1d1108",x"1f1208",x"1d1108",x"211309",x"1e1108",x"201309",x"1f1309",x"1f1208",x"1c1108",x"1b1008",x"1b1008",x"1b1008",x"1a1008",x"190f07",x"191008",x"1a1008",x"191008",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"191008",x"1a1008",x"1b1108",x"1c1108",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1b1108",x"1b1108",x"1b1008",x"1c1108",x"1c1108",x"1b1108",x"150e07",x"150e07",x"160f07",x"170f07",x"181007",x"181007",x"181007",x"180f07",x"1b1108",x"2c1c0a",x"34200b",x"3d250e",x"3b230e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"555555",x"363331",x"363433",x"3c3a39",x"3d3a39",x"3c3b3b",x"404040",x"3a3a3a",x"454545",x"323232",x"333333",x"313131",x"4b4b4b",x"505050",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b3b3b",x"444444",x"444444",x"363636",x"313131",x"323232",x"000000",x"000000",x"000000",x"4f4f4f",x"4d4d4d",x"363433",x"343332",x"322e2b",x"333232",x"333232",x"000000",x"000000",x"504e4d",x"504e4d",x"353433",x"353433",x"313131",x"333332",x"323232",x"323232",x"333333",x"313131",x"383838",x"595858",x"5d5956",x"323232",x"343434",x"333333",x"313131",x"333333",x"313131",x"333333",x"333333",x"313131",x"313131",x"3d3b38",x"3c3c3b",x"3c3c3b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2c190b",x"2c190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"4f3727",x"533f33",x"5f422e",x"5a3e29",x"583a26",x"4f3524",x"453024",x"4b2d19",x"4b2d19",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"53483e",x"53483e",x"4b4138",x"473e36",x"382e26",x"392f27",x"392f26",x"362c23",x"342a21",x"32271f",x"372c23",x"3d3026",x"3a2b21",x"3d2c20",x"3c2a1e",x"3c2c21",x"3f2d21",x"3a291e",x"3c2a1e",x"392619",x"3a271b",x"3b281c",x"433227",x"403024",x"3e2e23",x"3b2c21",x"3e2f25",x"3c2c22",x"35251b",x"38271c",x"392619",x"39271b",x"382517",x"392619",x"39291d",x"3d2e23",x"3d2f25",x"3d2f26",x"3b2d23",x"3b2c21",x"3c2b20",x"3c2b20",x"423024",x"402d21",x"372416",x"362012",x"392619",x"3f2c20",x"412f22",x"433023",x"422f22",x"402c1f",x"402d1e",x"443121",x"433023",x"412e20",x"3b2b20",x"3b2b20",x"3a2b21",x"3c2e24",x"3b2c22",x"3c2e24",x"3b2b21",x"392b21",x"392a20",x"37281e",x"3d2f26",x"382a20",x"3e3228",x"352b22",x"3c332b",x"4f453c",x"584d43",x"584d43",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a3a3a",x"333333",x"323232",x"333333",x"323232",x"383838",x"3c3c3c",x"3c3c3c",x"393939",x"3f3f3f",x"414141",x"464646",x"353535",x"333333",x"000000",x"000000",x"000000",x"323232",x"333333",x"323232",x"343130",x"353535",x"494949",x"4c4c4c",x"525252",x"4d4d4d",x"4c4c4c",x"332e2d",x"323232",x"393837",x"464646",x"575857",x"000000",x"000000",x"323232",x"323232",x"333333",x"434343",x"353636",x"323232",x"333333",x"343434",x"333333",x"2e2e2e",x"323232",x"3b3b3b",x"525251",x"3a3a3a",x"353535",x"333333",x"323232",x"343434",x"313131",x"434343",x"595959",x"5e5d5c",x"000000",x"323232",x"323232",x"323232",x"504d4b",x"504d4b",x"000000",x"201308",x"201308",x"271809",x"3b230d",x"37200c",x"2d1a0b",x"301c0d",x"2e1a0c",x"2d190b",x"28170a",x"28160a",x"2b170a",x"29170a",x"1d1108",x"1a1008",x"180f08",x"170f07",x"160e07",x"191007",x"201408",x"2d1c09",x"2f1d0a",x"2d1c0a",x"2b1a0a",x"2d1b0a",x"291709",x"251509",x"261509",x"261509",x"27160a",x"28170a",x"28170a",x"27170a",x"2a180b",x"29170b",x"2b190b",x"29170a",x"27170a",x"28170a",x"28170a",x"28170a",x"2b190c",x"2c190b",x"2b190b",x"28170b",x"2b190b",x"29180b",x"27160a",x"28160a",x"251509",x"26160a",x"251509",x"241509",x"27160a",x"27160a",x"29170a",x"251509",x"28160a",x"27160a",x"2a180a",x"27160a",x"2a180a",x"27160a",x"2a180b",x"2a180b",x"28160a",x"261609",x"261509",x"29170a",x"251509",x"261509",x"231409",x"27160a",x"26160a",x"261509",x"241509",x"241409",x"251509",x"1f1208",x"1e1109",x"1a1008",x"170f07",x"150e07",x"150e07",x"27160a",x"2e1a0b",x"301b0c",x"311b0c",x"321d0e",x"341f10",x"2e1c0d",x"2e1b0c",x"2c180a",x"2b180b",x"301b0c",x"2e190b",x"2d190b",x"2f1a0c",x"2f1a0b",x"2f1a0a",x"2e190a",x"2f1a0b",x"2e1a0b",x"2f1a0b",x"311b0c",x"2e1a0b",x"331c0d",x"301a0c",x"341d0d",x"321d0d",x"321d0d",x"341d0d",x"351e0e",x"341d0d",x"351e0d",x"38200e",x"371f0e",x"38200f",x"3a210f",x"361f0e",x"341e0e",x"341d0d",x"2e1a0b",x"311b0b",x"2e1a0b",x"2d190b",x"301b0b",x"321b0b",x"321b0c",x"361d0c",x"361d0c",x"341c0b",x"381e0d",x"361e0d",x"381f0e",x"381f0d",x"3f230f",x"38200e",x"3c220f",x"3b210f",x"371e0d",x"331c0c",x"371e0c",x"361d0c",x"331c0b",x"331c0c",x"2f1a0a",x"3a210e",x"351d0d",x"341c0c",x"351d0c",x"29170a",x"29180b",x"2d1a0c",x"2f1b0c",x"2f1a0b",x"27170a",x"29180b",x"311c0c",x"2c190b",x"321c0d",x"2d1a0b",x"3d250e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"313131",x"555555",x"333333",x"000000",x"313131",x"3b3b3b",x"474747",x"545454",x"323232",x"313131",x"323232",x"333333",x"313131",x"4b4b4b",x"3b3b3b",x"4f4f4f",x"4b4b4b",x"505050",x"494949",x"393939",x"333333",x"343434",x"484848",x"474747",x"444444",x"343434",x"363636",x"323232",x"323232",x"323232",x"000000",x"000000",x"474646",x"4c4a4a",x"4a4949",x"353332",x"343230",x"333232",x"000000",x"000000",x"000000",x"525050",x"525050",x"393736",x"353433",x"313131",x"333333",x"333333",x"323232",x"333333",x"323232",x"303030",x"534f4c",x"393736",x"333232",x"333333",x"333333",x"333333",x"323232",x"343434",x"332e2c",x"333333",x"323232",x"333333",x"4b4540",x"433f3b",x"363332",x"373432",x"343231",x"363432",x"4c4b4b",x"504e4e",x"5b5a5a",x"4c4b4b",x"424141",x"4f4f4f",x"535353",x"4d4d4d",x"4d4d4d",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2c190b",x"2c190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"533a29",x"573f30",x"61432f",x"573a28",x"593a27",x"523523",x"433024",x"482b19",x"482b19",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574d43",x"574d43",x"564c42",x"574d42",x"50463c",x"4f4439",x"52473e",x"4c4137",x"4b4036",x"473b32",x"483d33",x"4b3e34",x"45362b",x"3f2f23",x"3e2e22",x"3f2f24",x"443226",x"463428",x"49372a",x"453326",x"453326",x"483628",x"503e31",x"503e31",x"503f33",x"524033",x"524135",x"524235",x"504034",x"503e31",x"4b3a2d",x"4d3d32",x"433126",x"413024",x"413125",x"413226",x"423429",x"3f3024",x"403328",x"423328",x"433428",x"46362a",x"463528",x"433328",x"382619",x"362418",x"352317",x"3a291f",x"3d2d22",x"402f25",x"433328",x"413126",x"443224",x"4a392b",x"433429",x"44362a",x"423328",x"42352b",x"41352b",x"40342b",x"3f3329",x"42362c",x"43362d",x"423429",x"3f3026",x"413228",x"493b31",x"42352a",x"55493f",x"4f443a",x"4c4136",x"554b40",x"594e43",x"594e43",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"343434",x"323232",x"383838",x"3c3c3c",x"3c3c3c",x"3b3b3b",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"484848",x"494949",x"383838",x"434343",x"4a4a4a",x"454646",x"362f2a",x"313131",x"333333",x"575857",x"555454",x"000000",x"323232",x"323232",x"333333",x"565656",x"474747",x"414141",x"3d3c3b",x"323232",x"323131",x"333333",x"313131",x"323232",x"333333",x"373737",x"444444",x"535353",x"4a4a4a",x"4a4a4a",x"323232",x"333333",x"444444",x"585858",x"323232",x"323232",x"313131",x"313131",x"383838",x"444343",x"494746",x"000000",x"000000",x"201308",x"271809",x"3b230d",x"37200c",x"2d1a0b",x"301c0d",x"2e1a0c",x"2d190b",x"28170a",x"28160a",x"361d0d",x"29170a",x"1c1108",x"1d1108",x"221409",x"211309",x"211309",x"221409",x"231409",x"211309",x"1f1308",x"1c1108",x"1d1108",x"1d1108",x"1d1208",x"1e1208",x"1f1309",x"1f1309",x"1f1309",x"1e1208",x"150e07",x"1e1208",x"1e1208",x"1c1108",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"190f07",x"190f07",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"201308",x"201308",x"201208",x"211309",x"211309",x"211309",x"211308",x"211308",x"201308",x"201208",x"1f1208",x"201208",x"201308",x"201208",x"201308",x"1f1208",x"1e1208",x"1f1208",x"1e1108",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"190f08",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"1e1208",x"1e1208",x"1f1208",x"231409",x"231409",x"231409",x"1c1108",x"28160a",x"221308",x"25150a",x"1f1208",x"201308",x"231409",x"231409",x"241409",x"251509",x"26150a",x"251509",x"27160a",x"241509",x"231409",x"241409",x"25150a",x"27160a",x"26150a",x"25150a",x"26160a",x"25160a",x"29180b",x"27160a",x"28170a",x"251509",x"241509",x"26160a",x"251509",x"231409",x"221409",x"241409",x"241409",x"241409",x"251509",x"29170a",x"2a180b",x"2a180b",x"29170a",x"27160a",x"2b180b",x"26160a",x"25160a",x"2a180a",x"231509",x"2d190b",x"26160a",x"2b180b",x"26160a",x"2c190b",x"221409",x"25150a",x"28170a",x"28160a",x"28160a",x"2c180a",x"2d1a0b",x"2b190a",x"2f1c0b",x"311d0b",x"351f0c",x"38200d",x"3a220d",x"3c230d",x"3b230e",x"41270e",x"40260e",x"3d240d",x"331e0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"323232",x"333333",x"404040",x"4b4b4b",x"313131",x"3b3b3b",x"474747",x"343535",x"323232",x"333333",x"313131",x"333333",x"333333",x"313131",x"313131",x"4f4f4f",x"4b4b4b",x"505050",x"494949",x"343434",x"333333",x"343434",x"343434",x"313131",x"333333",x"303030",x"393939",x"323232",x"323232",x"323232",x"000000",x"000000",x"4c4a4a",x"4c4a4a",x"4a4949",x"343332",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"525050",x"000000",x"000000",x"000000",x"333333",x"333333",x"312823",x"323232",x"313131",x"323232",x"524f4b",x"504b45",x"2f2b29",x"333333",x"333333",x"333333",x"33302f",x"4d4e4e",x"4a4a4a",x"525252",x"5a5a5a",x"5e5e5e",x"5b5a5a",x"535151",x"363332",x"373432",x"343231",x"363432",x"4c4b4b",x"504e4e",x"5e5d5d",x"4c4b4b",x"343232",x"4f4f4f",x"525252",x"4d4d4d",x"5a5a5a",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2e1a0b",x"2e1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29170a",x"432917",x"5d4331",x"5f422d",x"5d3e2a",x"553826",x"563a26",x"473326",x"4e311e",x"4e311e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584e44",x"584e44",x"544a3e",x"554a3f",x"544a3e",x"554a40",x"54493e",x"574b41",x"584c42",x"51453b",x"4e4138",x"4e4034",x"4e3f33",x"48382c",x"4a3b2f",x"4d3c30",x"48392d",x"48362a",x"47382c",x"48392d",x"4d3e32",x"4e3e32",x"544438",x"544438",x"58493d",x"564538",x"5a493b",x"5a493c",x"5e4e41",x"5d4e42",x"5c4b3e",x"605043",x"5b4a3e",x"564438",x"55463a",x"534236",x"554539",x"564537",x"544436",x"574537",x"5a493c",x"584739",x"544334",x"564538",x"554439",x"514135",x"503f33",x"524337",x"534338",x"55463a",x"5b4d41",x"534336",x"57473a",x"57483a",x"524337",x"55473a",x"54473a",x"514337",x"52463c",x"53473c",x"55493f",x"584c41",x"53473b",x"594d42",x"584b40",x"56483d",x"52453a",x"514338",x"54473b",x"594d42",x"5a4f45",x"584c42",x"594f44",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"525252",x"4c4c4c",x"434343",x"323232",x"323232",x"414141",x"444444",x"3b3b3b",x"404040",x"4e4e4e",x"494949",x"525151",x"525151",x"323333",x"323333",x"333333",x"4d4d4d",x"454545",x"4c4c4c",x"4e4e4e",x"323232",x"323232",x"333333",x"323232",x"323232",x"323232",x"313131",x"323232",x"343434",x"494949",x"515151",x"4f4f4f",x"3f3f3f",x"393939",x"333333",x"323232",x"323232",x"323232",x"505050",x"484848",x"4d4d4d",x"4a4949",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"160e07",x"170f07",x"180f07",x"190f08",x"191008",x"1a1008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"1f1309",x"1f1209",x"1e1208",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1a1008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1008",x"1b1108",x"1b1008",x"1c1108",x"1d1108",x"1e1208",x"1f1208",x"1f1309",x"201309",x"201309",x"211309",x"211309",x"201309",x"201208",x"221409",x"231509",x"241509",x"25160a",x"25160a",x"25150a",x"25160a",x"25160a",x"25150a",x"25160a",x"25150a",x"241509",x"221409",x"211309",x"211309",x"211309",x"211309",x"221409",x"221409",x"211309",x"201208",x"1f1208",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"180f07",x"170f07",x"160e07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f07",x"1a1008",x"190f07",x"1b1108",x"1a1008",x"1c1108",x"1c1108",x"1b1008",x"1c1108",x"1d1108",x"1e1108",x"1f1208",x"201308",x"201309",x"201309",x"211309",x"211409",x"211409",x"221409",x"221409",x"221409",x"211309",x"231409",x"24150a",x"231409",x"221409",x"231509",x"24150a",x"24150a",x"231509",x"221409",x"221409",x"231409",x"241509",x"241509",x"231409",x"231409",x"241509",x"231409",x"201208",x"201208",x"201308",x"201308",x"1f1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1b1008",x"1a1008",x"191008",x"190f08",x"180f08",x"180f07",x"180f07",x"2c180a",x"2c180a",x"2d1a0b",x"2b190a",x"2f1c0b",x"311d0b",x"351f0c",x"38200d",x"3a220d",x"3c230d",x"3b230e",x"41270e",x"40260e",x"3d240d",x"331e0c",x"331e0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e3a39",x"3e3a39",x"393532",x"363432",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"333333",x"373737",x"3c3c3c",x"363636",x"313131",x"484848",x"323232",x"323232",x"323232",x"313131",x"323232",x"323232",x"343434",x"333333",x"333333",x"333333",x"343434",x"323232",x"333333",x"454545",x"333333",x"343434",x"333333",x"333333",x"313131",x"323232",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"323232",x"524f4b",x"504b45",x"000000",x"000000",x"000000",x"000000",x"373635",x"373635",x"413e3b",x"333333",x"323232",x"363534",x"353331",x"353433",x"393533",x"3a3532",x"33312f",x"373534",x"333130",x"5f5955",x"6a6661",x"5a5858",x"333232",x"343332",x"313131",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"351e0d",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"553b29",x"563f2f",x"583d2b",x"62432d",x"5b3b27",x"563c2b",x"4c3629",x"4b2f1c",x"4b2f1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"343434",x"424140",x"5c5c5c",x"333333",x"333333",x"2f2f2f",x"353535",x"474747",x"4d4d4d",x"4e4e4e",x"595959",x"5a5958",x"535251",x"323232",x"323232",x"313131",x"3c3d3d",x"3a3a3a",x"4e4e4e",x"4e4d4d",x"000000",x"000000",x"333333",x"333333",x"323232",x"323232",x"333333",x"323232",x"333333",x"343434",x"353535",x"505050",x"595959",x"4f4f4f",x"505050",x"5d5d5d",x"636363",x"5d5d5d",x"5c5c5c",x"525252",x"4b4b4b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"180f08",x"180f08",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f08",x"191008",x"191008",x"190f08",x"191008",x"191008",x"1a1008",x"191008",x"1a1008",x"1b1108",x"1b1108",x"1c1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1008",x"1a1008",x"1b1008",x"1c1108",x"1c1108",x"1c1108",x"1e1208",x"1f1209",x"201309",x"201309",x"201309",x"211409",x"221409",x"221409",x"211309",x"211309",x"211309",x"211409",x"231409",x"231409",x"231409",x"231409",x"231509",x"241509",x"231509",x"231409",x"221409",x"211309",x"231409",x"201309",x"211309",x"221409",x"211309",x"201208",x"1f1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"190f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"180f07",x"170f07",x"180f07",x"170f07",x"170f07",x"170f07",x"180f07",x"190f07",x"180f07",x"1a1008",x"191008",x"1b1108",x"1a1008",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1d1108",x"1f1208",x"201308",x"211309",x"211409",x"211409",x"221409",x"231509",x"231509",x"211409",x"211309",x"211309",x"221409",x"221409",x"211409",x"221409",x"231509",x"231409",x"231509",x"231409",x"211309",x"231509",x"241509",x"241509",x"221309",x"221409",x"25150a",x"241509",x"241509",x"211309",x"211309",x"201309",x"201309",x"1e1108",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1a1008",x"191008",x"180f08",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"1e1208",x"1e1208",x"1e1208",x"1f1309",x"231609",x"2b190a",x"301d0b",x"331f0c",x"37200c",x"3b220d",x"38210c",x"3e260d",x"39220c",x"37220c",x"331d0c",x"331d0c",x"000000",x"000000",x"000000",x"504b47",x"4d4844",x"453a33",x"3e3630",x"423831",x"393431",x"3f3935",x"3e3a39",x"393532",x"363432",x"363432",x"000000",x"000000",x"383431",x"3e3a37",x"383431",x"000000",x"000000",x"3a3431",x"36302c",x"393533",x"413a35",x"3a3431",x"3b3531",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"333333",x"3f3f3f",x"5d5d5d",x"323232",x"414141",x"363636",x"333333",x"333333",x"333333",x"323232",x"323232",x"313131",x"363636",x"3c3c3c",x"424242",x"323232",x"313131",x"333333",x"323232",x"333333",x"333333",x"323232",x"444444",x"323232",x"323232",x"323232",x"323232",x"313131",x"000000",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"626262",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"45413e",x"45413e",x"47423f",x"343333",x"343332",x"343332",x"363332",x"343231",x"393532",x"38332f",x"363433",x"353332",x"38312d",x"3f3b38",x"5d564f",x"353231",x"353332",x"343433",x"323232",x"343333",x"343333",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2b190b",x"2b190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"4e3525",x"584032",x"583c2b",x"6a4932",x"563d2b",x"553d2c",x"4c382c",x"50321f",x"50321f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323130",x"383432",x"5c5c5c",x"333333",x"333333",x"333333",x"323232",x"323232",x"303030",x"3e3e3e",x"4e4e4e",x"504f4f",x"000000",x"000000",x"323232",x"333333",x"373737",x"525252",x"545454",x"4e4e4e",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"333333",x"343434",x"323232",x"323232",x"323232",x"343434",x"3e3e3e",x"4a4a4a",x"4b4b4b",x"4e4e4e",x"5f5f5f",x"555555",x"565656",x"585858",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"180f07",x"190f08",x"1a1008",x"1b1008",x"1b1108",x"1b1108",x"1a1008",x"190f07",x"180f07",x"180f07",x"191008",x"1a1008",x"1b1008",x"1b1108",x"1c1108",x"1c1108",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1d1108",x"1d1108",x"1e1208",x"1f1309",x"1e1208",x"1f1209",x"1f1208",x"201208",x"221409",x"221409",x"221409",x"221409",x"211309",x"231409",x"24150a",x"241509",x"241509",x"241509",x"24150a",x"241509",x"241509",x"24150a",x"241509",x"241509",x"231409",x"231409",x"211309",x"221409",x"221409",x"201309",x"211409",x"211309",x"201309",x"1f1209",x"1c1108",x"1d1108",x"1b1108",x"1a1008",x"191008",x"180f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"191007",x"1a1109",x"191109",x"18100a",x"160f07",x"170f07",x"180f07",x"190f07",x"190f07",x"1a1008",x"191008",x"1b1108",x"1c1108",x"1d1108",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1e1208",x"201308",x"201309",x"211309",x"211309",x"211409",x"221409",x"211409",x"201208",x"1f1208",x"211309",x"221409",x"221409",x"221409",x"201308",x"201308",x"201208",x"211309",x"211309",x"231409",x"231409",x"221409",x"201308",x"201308",x"201208",x"221409",x"231409",x"231409",x"221409",x"221409",x"221409",x"221409",x"201309",x"1f1208",x"1d1108",x"1c1108",x"1a1008",x"191008",x"180f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"211309",x"231509",x"251609",x"2c190b",x"321d0c",x"39220e",x"3b220e",x"3d240f",x"40250e",x"3d230e",x"422810",x"3c240e",x"38210d",x"311d0c",x"311d0c",x"000000",x"000000",x"54504d",x"524d4a",x"4d4844",x"453a33",x"3e3630",x"423831",x"393431",x"3d3734",x"5d5b5a",x"676361",x"353231",x"353231",x"575654",x"3d3a39",x"383431",x"3e3a37",x"3a3633",x"3b3632",x"393532",x"3a3431",x"36302c",x"393533",x"413a35",x"3a3431",x"3b3531",x"000000",x"000000",x"333333",x"333333",x"313131",x"333333",x"303030",x"323232",x"595959",x"504f4f",x"414141",x"323232",x"313131",x"313131",x"333333",x"343434",x"333333",x"323232",x"313131",x"3c3a38",x"333130",x"323232",x"333333",x"323232",x"323232",x"33312f",x"3f3f3f",x"4d4d4d",x"535353",x"323232",x"323232",x"333333",x"343434",x"313131",x"585858",x"454545",x"5c5c5c",x"696969",x"606060",x"494949",x"5e5e5e",x"4b4b4b",x"353535",x"333333",x"3e3e3e",x"4e4e4e",x"353535",x"626262",x"626262",x"505050",x"3a3a3a",x"3f3f3f",x"5d5d5d",x"333333",x"323232",x"474747",x"595959",x"3f3f3f",x"3f3f3f",x"60605f",x"5a5a5a",x"3f3f3f",x"545454",x"45413e",x"47423f",x"343333",x"343332",x"343332",x"363332",x"343231",x"393532",x"383533",x"363433",x"353332",x"38312d",x"3f3b38",x"55504b",x"363332",x"353332",x"333332",x"323232",x"343333",x"343333",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"28170a",x"28170a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2a170b",x"4d3525",x"563f2f",x"583e2d",x"6a4831",x"5d4130",x"5a3f2d",x"4f3e31",x"4d3322",x"4d3322",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"170f07",x"170f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323130",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"323232",x"323232",x"393939",x"464646",x"000000",x"000000",x"000000",x"000000",x"373737",x"373737",x"484848",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"343434",x"3e3e3e",x"4a4a4a",x"4b4b4b",x"4e4e4e",x"585858",x"555555",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"645242",x"504134",x"635241",x"605342",x"5e5241",x"5f5241",x"625444",x"635443",x"615443",x"5e5241",x"38200e",x"311c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"1f140a",x"1f130a",x"1d1208",x"1d1108",x"1c1108",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1b1008",x"1b1008",x"1b1008",x"1b1008",x"1c1108",x"1c1108",x"1d1108",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1f1208",x"201309",x"211309",x"211409",x"221409",x"221409",x"201208",x"201308",x"221409",x"221409",x"231409",x"24150a",x"241509",x"241509",x"231409",x"231409",x"231409",x"221409",x"231509",x"231509",x"231509",x"221409",x"221409",x"221409",x"211409",x"201209",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"180f07",x"170f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"1e1308",x"1c1309",x"1a130c",x"1a120b",x"1a130c",x"191109",x"170f07",x"170f07",x"180f08",x"191008",x"1a1008",x"1b1108",x"1d1208",x"1d1208",x"1e1208",x"1e1208",x"1f1208",x"1f1308",x"1d1108",x"201309",x"211409",x"231509",x"221409",x"221409",x"231409",x"24150a",x"24160a",x"24150a",x"221409",x"241509",x"231409",x"221409",x"241509",x"25150a",x"24150a",x"25150a",x"241509",x"241509",x"241509",x"241509",x"24150a",x"241509",x"231409",x"221409",x"211309",x"201308",x"201208",x"1f1208",x"201208",x"1f1208",x"1e1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1a1008",x"191008",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"695444",x"28160a",x"281609",x"2d190b",x"311c0b",x"351e0c",x"3b220e",x"3f2510",x"3e240f",x"3e240f",x"3d220e",x"3f250e",x"3b220d",x"39220d",x"301c0c",x"301c0c",x"000000",x"686563",x"696564",x"63605d",x"56504c",x"59534f",x"5d5956",x"5c5856",x"5d5a58",x"605c59",x"5b5653",x"5d5a58",x"3a3431",x"3a3431",x"5c5b5b",x"575654",x"5f5c5b",x"636160",x"575250",x"3b3634",x"3d3a37",x"4f4c4a",x"54504e",x"575351",x"585654",x"3b3531",x"3b3633",x"3b3633",x"000000",x"333333",x"333333",x"313131",x"313131",x"323232",x"323232",x"323232",x"494949",x"4a4949",x"494949",x"505050",x"343434",x"343434",x"323232",x"4c4c4c",x"323232",x"616161",x"6c6966",x"616161",x"626262",x"313131",x"323232",x"606060",x"5a5a5a",x"323232",x"323232",x"434343",x"393939",x"3d3d3d",x"323232",x"333333",x"323232",x"515151",x"626161",x"616060",x"636363",x"4b4b4b",x"494949",x"5e5e5e",x"323232",x"353535",x"333333",x"444444",x"565656",x"353535",x"626262",x"616161",x"505050",x"3a3a3a",x"3f3f3f",x"5d5d5d",x"333333",x"3b3b3b",x"333333",x"595959",x"3f3f3f",x"3f3f3f",x"60605f",x"5a5a5a",x"434343",x"545454",x"545454",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f3b38",x"55504b",x"363332",x"353332",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"311c0d",x"311c0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"4e3424",x"563f31",x"5e412f",x"5a402d",x"5f4332",x"5e4534",x"584334",x"533727",x"533727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"180f07",x"180f07",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"343434",x"3c3c3c",x"333333",x"333333",x"383635",x"343130",x"323232",x"323131",x"353433",x"353535",x"393939",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"353535",x"353535",x"343434",x"343434",x"333232",x"323232",x"3a3a3a",x"393939",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"4e4e4e",x"4b4b4b",x"373737",x"373737",x"323232",x"353535",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"645242",x"504134",x"635241",x"605342",x"5e5241",x"5f5241",x"625444",x"635443",x"615443",x"5e5241",x"5d503f",x"5d4f3f",x"5f5241",x"655543",x"675544",x"645745",x"655746",x"645746",x"645746",x"645745",x"615543",x"645544",x"655545",x"655443",x"665544",x"625444",x"655645",x"665444",x"645644",x"665443",x"5f5241",x"5e5040",x"615040",x"675141",x"635242",x"685342",x"695243",x"655141",x"5e4e3e",x"5d4b3c",x"605040",x"625040",x"604e3e",x"614c3d",x"594839",x"5a4b3c",x"564839",x"4b3e31",x"473b2f",x"4b3e32",x"4d4133",x"4b3e32",x"4c4033",x"5a4c3e",x"5f4b3d",x"645141",x"614f3f",x"685444",x"655041",x"645040",x"685645",x"615443",x"6b5746",x"6a5b49",x"665646",x"675646",x"625443",x"625242",x"635443",x"675847",x"685847",x"685847",x"665747",x"655645",x"655645",x"655747",x"665847",x"645646",x"655747",x"675949",x"645848",x"645848",x"665848",x"6a5544",x"695545",x"685544",x"665546",x"655545",x"655546",x"615243",x"645444",x"635747",x"645847",x"665747",x"645747",x"605445",x"625647",x"645848",x"5f5344",x"635848",x"5e5142",x"5b4d3d",x"5d4b3c",x"625040",x"605041",x"625142",x"625242",x"675747",x"6c5c4c",x"645645",x"645645",x"645745",x"645745",x"625545",x"625141",x"5b4f3f",x"5c4f3f",x"594c3d",x"5b4f3f",x"5d503f",x"564a3b",x"5a4e3e",x"564939",x"594d3d",x"594d3c",x"584b3b",x"554537",x"614f3f",x"635142",x"605140",x"5e5140",x"615442",x"5f5141",x"615342",x"635444",x"655645",x"645544",x"605341",x"5f5241",x"5e5140",x"645343",x"675543",x"675645",x"675645",x"655746",x"625545",x"655846",x"645747",x"625645",x"635645",x"665848",x"665645",x"665645",x"685646",x"695747",x"685647",x"625444",x"685645",x"635242",x"635242",x"665443",x"695444",x"695444",x"311b0b",x"311b0c",x"331c0c",x"38200e",x"3b210e",x"3b210e",x"3c230e",x"3d230f",x"3f240f",x"3e230f",x"3b230f",x"39220e",x"311d0b",x"311d0b",x"000000",x"605d5c",x"605d5c",x"585451",x"3a3430",x"5d5651",x"3e3631",x"3e3733",x"3e3631",x"3e3632",x"5a5653",x"5c5856",x"393431",x"393431",x"5a5957",x"63615f",x"3b3634",x"4d4b4a",x"605d5c",x"5b5856",x"5a5957",x"5a5856",x"5a5856",x"585756",x"4d4c4b",x"353332",x"333131",x"333131",x"000000",x"000000",x"323232",x"323232",x"333333",x"333333",x"33312f",x"333333",x"313131",x"313131",x"333333",x"464646",x"3a3a3a",x"464646",x"545454",x"636363",x"5f5f5f",x"5c5c5c",x"535353",x"3b3b3b",x"4f4e4e",x"333333",x"535251",x"676564",x"313131",x"323232",x"323232",x"333333",x"4b4b4b",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"4c4c4c",x"313131",x"323232",x"323231",x"303131",x"333333",x"333333",x"313131",x"323232",x"383838",x"323232",x"313131",x"323232",x"323232",x"333333",x"313131",x"5e5b59",x"313131",x"313131",x"333333",x"343434",x"313131",x"323232",x"303030",x"322e2c",x"313131",x"343434",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"341e0d",x"341e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"41291a",x"4e3a2d",x"5e412f",x"664732",x"624531",x"654937",x"5b4637",x"513320",x"513320",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"160e07",x"160e07",x"170f07",x"180f08",x"191008",x"190f07",x"190f08",x"180f08",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"180f07",x"1b1108",x"1b1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"414141",x"3e3e3e",x"333333",x"343434",x"3c3c3c",x"333333",x"333333",x"4d4c4b",x"383635",x"323232",x"333333",x"333333",x"3c3c3c",x"464646",x"3b3a38",x"363434",x"322a26",x"312d2a",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434343",x"3a3a3a",x"353535",x"393939",x"353535",x"333232",x"323232",x"3a3a3a",x"393939",x"323232",x"333333",x"333333",x"313131",x"000000",x"545454",x"474747",x"393837",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"555555",x"5d5d5c",x"595959",x"4b4b4b",x"4a4a4a",x"353535",x"343434",x"373737",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"615342",x"615342",x"5f5342",x"655443",x"655443",x"665342",x"665443",x"665544",x"695444",x"645544",x"635645",x"645444",x"605140",x"605442",x"625543",x"645443",x"655241",x"615241",x"615140",x"625241",x"625443",x"615242",x"605343",x"655442",x"665343",x"695443",x"685444",x"645645",x"645644",x"625444",x"625342",x"675242",x"5f5141",x"5a4d3e",x"5a4e3d",x"635141",x"695141",x"615040",x"625141",x"5a493a",x"5a4a3a",x"5b4a3b",x"564839",x"574739",x"594b3b",x"574a3b",x"594a3c",x"524637",x"493e31",x"463b2f",x"453a2e",x"514437",x"514033",x"4b3c30",x"5a4b3c",x"614e3e",x"695444",x"615141",x"635443",x"5b4c3d",x"615242",x"5d4e3e",x"605040",x"645443",x"635645",x"5d4d3e",x"695646",x"695444",x"685343",x"6b5545",x"6d5645",x"6c5645",x"695646",x"645746",x"675343",x"625545",x"625444",x"635445",x"635746",x"675a4a",x"67594a",x"645847",x"615344",x"605040",x"605040",x"605141",x"5f5040",x"5d5140",x"5d5140",x"605140",x"5f5243",x"615445",x"625445",x"605343",x"615243",x"5d5142",x"615141",x"605344",x"635443",x"655243",x"635445",x"695b4c",x"635645",x"5c4e3f",x"5d5141",x"645443",x"615544",x"625645",x"685847",x"665645",x"655745",x"645645",x"635343",x"645343",x"655544",x"544235",x"655040",x"594c3c",x"5a4c3c",x"625140",x"5e4d3d",x"604f3e",x"5b4c3b",x"5f4d3d",x"5f4d3d",x"5f4e3e",x"5a4d3d",x"5e4e3f",x"605040",x"645242",x"5f5241",x"665342",x"615241",x"5f5140",x"615342",x"625544",x"625645",x"675544",x"675544",x"665443",x"605140",x"665342",x"625242",x"635443",x"605241",x"5c503f",x"605241",x"625544",x"625545",x"625545",x"635545",x"625645",x"645846",x"655848",x"655847",x"665947",x"635444",x"655443",x"645443",x"615443",x"615342",x"665443",x"625443",x"615443",x"371f0d",x"381f0d",x"341c0c",x"371f0d",x"3e2310",x"3f240f",x"3f2410",x"412510",x"402510",x"402611",x"3a210e",x"351f0d",x"2e1a0b",x"2e1a0b",x"000000",x"676462",x"676462",x"55504d",x"423931",x"5c5551",x"605954",x"5d5753",x"514842",x"493e36",x"544d49",x"534d4a",x"3a332f",x"3a332f",x"616161",x"545454",x"343332",x"333333",x"494542",x"4c4847",x"444241",x"3d3a3a",x"383432",x"494341",x"4c4b4b",x"333333",x"343434",x"343434",x"000000",x"000000",x"313131",x"2f2f2f",x"333333",x"343434",x"333333",x"545454",x"353535",x"382319",x"323232",x"404040",x"5f5f5f",x"4b4b4b",x"494949",x"454545",x"343434",x"323232",x"333333",x"333333",x"323232",x"333333",x"333333",x"514f4d",x"5c5b5b",x"323232",x"323232",x"4d4d4d",x"323232",x"303030",x"323232",x"343434",x"343434",x"343434",x"333333",x"454545",x"4e4e4e",x"434343",x"323232",x"333333",x"313131",x"323232",x"323232",x"494745",x"525252",x"323232",x"323232",x"313131",x"333333",x"323232",x"333333",x"5f5c5b",x"323232",x"333333",x"323232",x"313131",x"333333",x"323232",x"333333",x"434343",x"3c3a39",x"333333",x"323232",x"5b5b5b",x"454545",x"343434",x"323232",x"323232",x"333333",x"505050",x"5c5c5c",x"616161",x"5b5b5b",x"545454",x"4c4c4c",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2c190b",x"2c190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"25150a",x"513727",x"4d392c",x"5e432f",x"654732",x"5d4231",x"604634",x"524338",x"4d3323",x"4d3323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"160f07",x"160e07",x"170f07",x"191008",x"1b1108",x"1b1108",x"1a1108",x"191008",x"170f08",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"191008",x"1c1108",x"1c1108",x"5e432d",x"543d28",x"5c432d",x"533c28",x"453220",x"644932",x"6c4f35",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595958",x"474747",x"414141",x"363636",x"434343",x"575757",x"3b3b3b",x"323232",x"312f2e",x"585552",x"434343",x"3e3e3e",x"454544",x"515151",x"4a4a4a",x"3b3a38",x"363434",x"322a26",x"313131",x"323232",x"323232",x"343434",x"000000",x"000000",x"000000",x"4a4a4a",x"434343",x"434343",x"5c5c5c",x"5e5e5e",x"606060",x"636363",x"626262",x"606060",x"606060",x"666665",x"333333",x"323232",x"323232",x"333333",x"545454",x"474747",x"393837",x"363636",x"323232",x"383838",x"333333",x"333333",x"000000",x"000000",x"5a5a5a",x"575757",x"555555",x"606060",x"505050",x"4d4d4d",x"515151",x"5b5b5b",x"555555",x"323232",x"313131",x"313131",x"000000",x"000000",x"000000",x"615343",x"615343",x"5f5343",x"625645",x"615343",x"625443",x"625443",x"625544",x"645646",x"625644",x"615644",x"635645",x"635645",x"635645",x"645746",x"655846",x"655746",x"645645",x"645645",x"655443",x"615444",x"615444",x"615343",x"615443",x"5e5140",x"5f5140",x"5f5140",x"615544",x"645746",x"655846",x"665847",x"665847",x"615343",x"645544",x"625342",x"665443",x"665544",x"675544",x"615141",x"605242",x"625544",x"5e5141",x"5a4e3e",x"5e4d3e",x"5d493a",x"634e3e",x"654e3f",x"514335",x"574235",x"4f3e32",x"544436",x"3c2f26",x"453a2f",x"554538",x"59483a",x"675342",x"65503f",x"625443",x"645746",x"5f5342",x"5f5342",x"645746",x"675948",x"685b49",x"685a49",x"685948",x"665645",x"695645",x"6b5544",x"685847",x"645746",x"625645",x"615443",x"615545",x"5f5343",x"5e5242",x"5b4f40",x"5c5042",x"524638",x"574b3c",x"5b4f41",x"5f5242",x"5d4e3f",x"594a3c",x"655647",x"5d4b3c",x"5c4b3c",x"5e4c3d",x"594a3b",x"57493a",x"5a4a3c",x"5d4e3d",x"5e5040",x"5c4f40",x"5a4d3d",x"5b4e3e",x"574b3c",x"564a3b",x"5e4c3c",x"604d3e",x"624e3e",x"5b4e3f",x"615443",x"675948",x"625344",x"665545",x"635545",x"655544",x"655444",x"675343",x"645545",x"645645",x"655444",x"665646",x"6a5343",x"564639",x"635141",x"635242",x"655443",x"594c3d",x"5d4e3f",x"5d4e3f",x"483d30",x"56493a",x"594d3d",x"5e4e3e",x"574b3c",x"5d5241",x"5e5342",x"5c4f3f",x"594c3d",x"645747",x"635645",x"635645",x"645645",x"645746",x"645647",x"665847",x"655846",x"665847",x"665948",x"665948",x"695a48",x"5c5040",x"695847",x"695746",x"695847",x"655846",x"655847",x"665848",x"655847",x"675948",x"665645",x"695645",x"625344",x"675645",x"675645",x"675645",x"665746",x"665847",x"655847",x"655846",x"645645",x"665544",x"39200e",x"3b210f",x"3c230f",x"3c2210",x"3e230f",x"3f230f",x"40250f",x"3f2410",x"3c220f",x"3d230f",x"39200d",x"331e0c",x"2c190b",x"2c190b",x"000000",x"625e5b",x"625e5b",x"554f4b",x"3b332d",x"625b56",x"5d5753",x"5e5450",x"605a56",x"5d534d",x"4c433c",x"58514c",x"3d3631",x"3d3631",x"5f5e5d",x"505050",x"333333",x"515151",x"545454",x"525252",x"303030",x"323232",x"333333",x"4d4d4d",x"505050",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"333333",x"313131",x"323232",x"313131",x"4a4a4a",x"4e4e4e",x"323232",x"3b3b3b",x"434343",x"575756",x"333333",x"343434",x"323232",x"313131",x"323232",x"323232",x"333333",x"333333",x"333231",x"343434",x"504e4c",x"5c5b5b",x"4c4c4c",x"4e4e4f",x"333333",x"333333",x"333333",x"333333",x"333333",x"000000",x"343434",x"333333",x"454545",x"4e4e4e",x"434343",x"323232",x"333333",x"313131",x"323232",x"323232",x"494745",x"323232",x"333333",x"323232",x"323232",x"4e4e4e",x"313131",x"323232",x"333333",x"3c3c3c",x"4f4f4f",x"333333",x"323232",x"323232",x"333333",x"323232",x"414141",x"565656",x"525151",x"535353",x"5b5b5b",x"454545",x"343434",x"323232",x"313131",x"333333",x"505050",x"5c5c5c",x"676767",x"5d5d5d",x"5e5e5e",x"3f3f3f",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"251509",x"251509",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"4b301f",x"4a372d",x"5a402e",x"624731",x"573f2f",x"564336",x"59493d",x"523928",x"523928",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"170f07",x"160e07",x"160e07",x"180f08",x"1a1008",x"1b1108",x"1a1108",x"191008",x"180f08",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"1a1008",x"1d1108",x"5c422b",x"5e432d",x"543d28",x"5c432d",x"533c28",x"453220",x"644932",x"6c4f35",x"6c4f35",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595958",x"595958",x"595959",x"474747",x"4a4a4a",x"454545",x"4c423c",x"4a4a4a",x"4b4a4a",x"494949",x"434241",x"3f3e3d",x"3e3b39",x"444444",x"494949",x"515151",x"54504d",x"575757",x"3d3d3d",x"333333",x"333333",x"333333",x"313131",x"323232",x"616160",x"545455",x"4a4a4a",x"5a5a5a",x"333333",x"313131",x"323232",x"373433",x"454545",x"3c3c3c",x"4d4d4d",x"4b4a4a",x"616161",x"5f5f5f",x"333333",x"323232",x"5c5c5b",x"5b5b5b",x"616161",x"414141",x"323232",x"383838",x"333333",x"323232",x"3e3e3e",x"484848",x"5c5c5c",x"5a5a5a",x"4a4a4a",x"4e4e4e",x"3b3b3b",x"333333",x"333333",x"4f4f4f",x"5b5b5b",x"595959",x"323232",x"313131",x"313131",x"000000",x"000000",x"605040",x"605040",x"625041",x"5f4f3f",x"6a5242",x"6b5242",x"5f5241",x"6b5242",x"605140",x"5c4e3e",x"665141",x"665040",x"655141",x"675241",x"5f5141",x"625241",x"605140",x"5a4d3c",x"5b4d3d",x"5a4d3c",x"63503f",x"635140",x"665141",x"645040",x"5e5140",x"5d5040",x"5c503f",x"605241",x"615544",x"665747",x"655747",x"605343",x"675645",x"645241",x"665544",x"5d503f",x"60503f",x"5f5140",x"5e5140",x"614f3f",x"5a483a",x"5c4b3c",x"604e3e",x"574637",x"504335",x"4d4032",x"504033",x"5d493a",x"524335",x"544336",x"594a3b",x"42352a",x"42372c",x"483b30",x"584b3c",x"6a5242",x"604e3e",x"665443",x"635443",x"655746",x"665545",x"645443",x"6c5a4a",x"685545",x"695645",x"695747",x"635142",x"635243",x"665545",x"665645",x"635645",x"625545",x"615545",x"5d5141",x"615444",x"655545",x"665645",x"615544",x"625545",x"695645",x"685747",x"5f5242",x"635141",x"685141",x"665343",x"665848",x"594d3d",x"614f3f",x"5b4e3f",x"675141",x"5f5040",x"615444",x"625445",x"645444",x"5f5140",x"5b4c3d",x"5e4d3d",x"5d4d3f",x"605140",x"605342",x"5a4f3f",x"5f5142",x"665745",x"615544",x"635646",x"5a5040",x"6b5e4d",x"675646",x"625645",x"5d5140",x"5e5140",x"615644",x"615644",x"615545",x"5e5141",x"604f40",x"524336",x"645545",x"635645",x"5e5141",x"5c503f",x"5c5040",x"615343",x"615544",x"574b3c",x"615544",x"655343",x"665343",x"675646",x"655544",x"635342",x"645141",x"615141",x"645141",x"665443",x"635241",x"615543",x"5d5140",x"5e5140",x"625141",x"655545",x"665645",x"655645",x"645443",x"665645",x"5f5241",x"615544",x"605343",x"5f5342",x"665847",x"665848",x"645847",x"665948",x"655644",x"665544",x"655544",x"645745",x"685847",x"685a49",x"675a49",x"665948",x"675746",x"685847",x"625645",x"381f0e",x"3a200f",x"3b210f",x"3b210f",x"3d230f",x"3b210f",x"391f0d",x"3b210e",x"3f240f",x"412511",x"3a220e",x"321e0d",x"2b190b",x"2b190b",x"000000",x"615d5b",x"595653",x"514e4c",x"625e5b",x"4e453f",x"48403a",x"4f453d",x"483b30",x"4c4139",x"59514d",x"615c59",x"3f3731",x"3f3731",x"626262",x"4e4e4e",x"555555",x"545454",x"535353",x"565656",x"5c5c5c",x"5f5f5f",x"606060",x"525252",x"4e4e4e",x"343434",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"323232",x"343333",x"3b3b3b",x"333333",x"312f2f",x"333333",x"5e5e5e",x"545353",x"595857",x"383838",x"362e2a",x"333333",x"313131",x"323232",x"333333",x"333333",x"323232",x"333231",x"323232",x"3b3b3b",x"3d3d3d",x"5b5b5b",x"333333",x"333333",x"333333",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"313131",x"323232",x"616161",x"323232",x"323232",x"333333",x"333231",x"696765",x"323232",x"333333",x"323232",x"313131",x"343434",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"333333",x"303030",x"323232",x"313131",x"333333",x"323232",x"323232",x"313131",x"363636",x"323232",x"3d3d3d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"2d190b",x"2d190b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"543a27",x"48352a",x"5f4431",x"583e2d",x"553f30",x"524134",x"544539",x"4c3425",x"4c3425",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"664a32",x"694c33",x"816041",x"7c5b3e",x"7a593d",x"7d5c3f",x"6a4f36",x"745439",x"805f42",x"816043",x"826144",x"876446",x"866345",x"836143",x"8b6848",x"886547",x"8f6c4b",x"825f43",x"8b694a",x"866143",x"835f41",x"815e40",x"805d3f",x"815e41",x"896444",x"8d6948",x"916d4c",x"876446",x"926d4d",x"946f4e",x"946f4e",x"876343",x"8d6948",x"8c6747",x"926d4b",x"8b6646",x"8c6748",x"926c4a",x"926d4c",x"926b49",x"956f4e",x"946e4d",x"946e4d",x"956f4e",x"906b4b",x"916b4a",x"97714f",x"956f4e",x"98724e",x"8f6948",x"936d4c",x"876141",x"876141",x"845f3f",x"7c5a3a",x"896342",x"8d6746",x"916c4a",x"946e4d",x"906948",x"936c4b",x"956f4d",x"946e4d",x"886243",x"8a6545",x"8c6646",x"8d6949",x"7f5d3f",x"846143",x"866243",x"866444",x"8c6846",x"916c4d",x"8a6548",x"8b6849",x"8c6849",x"8b6748",x"805d40",x"906b4b",x"896647",x"8b6747",x"8b6646",x"8a6648",x"815d40",x"825e40",x"7b593b",x"7b593b",x"775639",x"846142",x"856243",x"826043",x"7c5a3f",x"866445",x"836145",x"7b5b3f",x"6e4f35",x"725338",x"694c33",x"5a422d",x"684c33",x"715138",x"6e5036",x"674c32",x"6a4e35",x"6a4e35",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"606060",x"606060",x"4f4f4f",x"454545",x"474747",x"434343",x"434343",x"464646",x"4b4b4b",x"444444",x"483f3a",x"474341",x"4b4744",x"3f3733",x"494441",x"4d4d4d",x"494949",x"505050",x"4d4d4d",x"5b5b5b",x"5a5a5a",x"333333",x"323232",x"333333",x"545353",x"5f5f5f",x"646464",x"313131",x"323232",x"333333",x"333333",x"373433",x"373737",x"3c3c3c",x"4e4e4e",x"4d4947",x"5c5c5c",x"5d5d5c",x"4a4a4a",x"323232",x"323232",x"4e4e4e",x"444444",x"3d3d3d",x"3b3b3b",x"636160",x"323232",x"333333",x"3e3e3e",x"484848",x"525252",x"5b5a5a",x"4a4a4a",x"484848",x"2f2e2d",x"323232",x"323232",x"4f4f4f",x"5c5c5c",x"5f5e5e",x"323232",x"323232",x"323232",x"000000",x"000000",x"615141",x"615141",x"625141",x"614f3f",x"604e3f",x"624f3f",x"625040",x"614d3e",x"625040",x"5e4f40",x"5c4e3d",x"5b4d3d",x"5d4e3e",x"604d3e",x"615040",x"5b4e3e",x"644e3e",x"664f40",x"644f3f",x"664f3f",x"654f3f",x"5c4a3b",x"5c4b3c",x"5b4a3b",x"584a3b",x"5f4c3d",x"634e3e",x"574939",x"564a3b",x"574a3b",x"5d4d3d",x"584a3a",x"5a4b3c",x"625242",x"615141",x"5d5040",x"5b4e3e",x"5e4e3e",x"5d5040",x"5d4d3f",x"5b4c3e",x"58483a",x"584c3d",x"5e4e3f",x"453a2d",x"524437",x"504236",x"514236",x"4c3f33",x"503f32",x"4d3f32",x"554437",x"3e3227",x"463a2e",x"58493a",x"584a3a",x"605241",x"615342",x"605241",x"605343",x"625645",x"615444",x"655343",x"6b5847",x"645747",x"5b4c3c",x"615545",x"625545",x"605444",x"615545",x"5f5242",x"615645",x"625645",x"615545",x"625745",x"645746",x"645746",x"645646",x"635646",x"605345",x"615444",x"605445",x"625645",x"665a49",x"665949",x"665948",x"615343",x"5f5242",x"605344",x"615545",x"5f5243",x"5d5142",x"5f5040",x"5e4e3f",x"5b5040",x"594d3e",x"594c3c",x"564a3b",x"56493a",x"594b3c",x"56493a",x"594d3d",x"5c4e3e",x"5d5040",x"605342",x"685b49",x"6a5c4a",x"675948",x"5e5243",x"5e5140",x"5e5141",x"605242",x"5e5141",x"5d5141",x"594d3d",x"564a3b",x"584b3c",x"5b4d3c",x"5d4d3d",x"5d4f3f",x"5d5040",x"615241",x"605242",x"605342",x"605342",x"665948",x"665a48",x"675948",x"665948",x"5d5040",x"5d5242",x"5c4f3f",x"5d5140",x"5d5140",x"605243",x"5d4d3e",x"58493c",x"625141",x"5d5141",x"564b3c",x"4e4133",x"5c4f40",x"615344",x"5f5343",x"5b4f40",x"5d5141",x"605141",x"625242",x"655445",x"605242",x"615443",x"605344",x"5f5443",x"5f5243",x"5f5242",x"5e5040",x"635141",x"554638",x"6b5242",x"6c5343",x"6a5343",x"695444",x"625645",x"645646",x"3b2210",x"3a210f",x"361e0d",x"371e0d",x"39200e",x"391f0d",x"351d0c",x"361e0d",x"39200d",x"3b230e",x"351f0d",x"2c1a0b",x"25160a",x"25160a",x"000000",x"000000",x"514e4c",x"433f3b",x"403833",x"463a30",x"453a31",x"4f453d",x"483b30",x"4c4139",x"423b36",x"443d38",x"403732",x"403732",x"4e4e4e",x"4d4d4d",x"474747",x"4d4d4d",x"252525",x"323232",x"323232",x"323232",x"3a3a3a",x"5b5b5b",x"616161",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a3a3a",x"3f3f3f",x"333333",x"333333",x"323232",x"5d5d5d",x"403f3e",x"595959",x"373737",x"4a4a4a",x"323232",x"313131",x"353535",x"474747",x"494949",x"4d4d4d",x"636363",x"505050",x"5a5a5a",x"343434",x"333333",x"545454",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"323232",x"323232",x"323232",x"333333",x"343434",x"323232",x"5d5d5d",x"4a4a4a",x"323232",x"323232",x"323232",x"353535",x"323232",x"323232",x"323232",x"3b3b3b",x"3d3d3d",x"323232",x"333333",x"343434",x"323232",x"323232",x"333332",x"323232",x"323232",x"323232",x"353535",x"363130",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"311c0c",x"311c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"543a29",x"4c3b31",x"634733",x"5f4331",x"533d2f",x"584031",x"514135",x"4f3321",x"4f3321",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"78583c",x"78583c",x"73553a",x"75563c",x"79593e",x"74563b",x"5e452f",x"614831",x"684c33",x"6e5136",x"705339",x"77583c",x"75573b",x"7b5a3d",x"7d5d42",x"806043",x"7a5a3e",x"7b5b40",x"825f42",x"805e41",x"825e42",x"7d5a3e",x"715236",x"705136",x"78593b",x"77563b",x"78563a",x"7e5c3f",x"856547",x"876447",x"866546",x"846345",x"856345",x"866447",x"856245",x"896646",x"8e6949",x"8e6949",x"896446",x"876446",x"836143",x"846244",x"805d42",x"846143",x"856143",x"825f41",x"886547",x"876446",x"826040",x"8b6646",x"805c3d",x"825e40",x"805c3d",x"7d5a3b",x"714f33",x"704f34",x"775536",x"7d5a3c",x"7a573a",x"835d40",x"8c6849",x"8a6646",x"866445",x"846245",x"816144",x"866345",x"846145",x"7d5c41",x"8a6748",x"866446",x"846244",x"805f43",x"7f5d41",x"7d5b3e",x"7b5a3d",x"7c5b3f",x"815d40",x"825e40",x"7f5d41",x"805e42",x"74553a",x"75573c",x"77573b",x"7a593c",x"7a583b",x"755539",x"6b4c31",x"67492f",x"705136",x"63472f",x"64482f",x"6e4f35",x"72563b",x"75583d",x"72553a",x"6e5138",x"715339",x"694d35",x"5d442d",x"674c34",x"684d35",x"6c5037",x"6c4f36",x"6a4d34",x"6a4d34",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"606060",x"606060",x"4d4d4d",x"4c4c4c",x"525252",x"505050",x"454545",x"494949",x"4c4c4c",x"535353",x"4c4b4a",x"313130",x"2f2c29",x"32302f",x"323232",x"333333",x"343333",x"363433",x"332f2d",x"333333",x"535353",x"4c4c4c",x"313131",x"333333",x"565656",x"3e3e3e",x"323232",x"323232",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595959",x"565656",x"595654",x"4a4a4a",x"4f4f4f",x"4b4b4b",x"454545",x"444444",x"4a4a4a",x"4c4c4c",x"474747",x"474747",x"606060",x"626262",x"5d5d5d",x"494949",x"4a4a4a",x"454545",x"3c3c3c",x"333333",x"333333",x"333333",x"605f5f",x"5e5d5d",x"5e5e5e",x"323232",x"323232",x"000000",x"000000",x"5d4e3e",x"5d4e3e",x"5b4e3d",x"5b4e3d",x"685141",x"675140",x"5d4b3c",x"604e3e",x"59473b",x"584839",x"534536",x"57493a",x"584a3b",x"5a4d3c",x"5b4e3d",x"584a3b",x"5b4d3d",x"5a4c3c",x"594c3c",x"594c3c",x"574a3a",x"4b3e30",x"4b3e30",x"4e3f32",x"4e3f32",x"524436",x"62503f",x"5f4e3f",x"5b4d3d",x"594b3d",x"5d4e3e",x"62503f",x"5c4e3f",x"574a3c",x"544839",x"5f5141",x"604e3f",x"614f3e",x"614e3e",x"5a493a",x"564638",x"574738",x"584235",x"564336",x"503f33",x"3a2d24",x"4e3f32",x"4e4033",x"4c3e32",x"453a2e",x"4b4033",x"43382d",x"544739",x"594d3d",x"5a4d3d",x"44372b",x"594939",x"665241",x"665443",x"635645",x"625645",x"635544",x"5b4f40",x"625645",x"625645",x"5d5140",x"625645",x"615645",x"615645",x"645746",x"625645",x"645746",x"635645",x"645646",x"625545",x"625745",x"625545",x"615343",x"615142",x"625242",x"615342",x"605343",x"615543",x"625645",x"625645",x"605343",x"5f5242",x"5e5242",x"5f5242",x"5f5242",x"635343",x"645342",x"6a5243",x"5c5041",x"4c4033",x"4c3f32",x"4c3e31",x"615142",x"57483a",x"5c4c3e",x"615141",x"5d5141",x"645645",x"675444",x"665343",x"645647",x"675a49",x"645748",x"605344",x"5c5040",x"5f5141",x"655443",x"625645",x"645646",x"615545",x"5e5142",x"5f5342",x"605343",x"605444",x"5f5242",x"5f5242",x"635645",x"5e5141",x"615343",x"625342",x"5f5041",x"635645",x"635645",x"5d5141",x"655746",x"645746",x"5d5141",x"615544",x"615544",x"5b4f40",x"625644",x"5d5140",x"5d5140",x"534739",x"5b4f40",x"5d5140",x"625443",x"625544",x"5d5040",x"615343",x"645141",x"645243",x"5e5241",x"615141",x"5f5040",x"5f5242",x"5f5142",x"645243",x"6e5445",x"5f5242",x"605343",x"625645",x"635645",x"645645",x"635443",x"635444",x"635545",x"665847",x"685847",x"331c0c",x"331c0c",x"341d0d",x"341d0d",x"351e0d",x"341d0c",x"341d0c",x"351d0d",x"331d0c",x"301c0b",x"2d1a0a",x"241509",x"201409",x"201409",x"000000",x"000000",x"000000",x"353535",x"343434",x"343231",x"333231",x"32251c",x"353230",x"383432",x"373432",x"3a3532",x"3a3532",x"524e4c",x"524e4c",x"464646",x"424242",x"454545",x"464545",x"323232",x"323232",x"323232",x"3a3a3a",x"575757",x"313131",x"343434",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"454545",x"323232",x"323232",x"3a3a3a",x"5e5d5b",x"313131",x"333333",x"343434",x"313131",x"343434",x"343434",x"2e2e2e",x"474747",x"494949",x"4d4d4d",x"636363",x"5b5b5b",x"313131",x"333333",x"313131",x"545454",x"585858",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303131",x"333333",x"323232",x"323232",x"323232",x"333333",x"323232",x"323232",x"5f5f5e",x"5e5d5c",x"33302e",x"323232",x"323232",x"353535",x"323232",x"323232",x"333232",x"3b3b3b",x"3d3d3d",x"323232",x"333333",x"343434",x"323232",x"323232",x"333332",x"323232",x"323232",x"323232",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434343",x"000000",x"000000"),
(x"000000",x"2d1a0b",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"321d0d",x"493324",x"574336",x"604432",x"5f4331",x"533e31",x"523e30",x"5d4738",x"513524",x"513524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"7b5b3e",x"7b5b3e",x"72553a",x"725439",x"79593d",x"6e5137",x"4f3926",x"5b432d",x"604530",x"644931",x"6c4f36",x"6e5139",x"72543a",x"6c4f36",x"6d4f36",x"715439",x"6f5138",x"6e4f37",x"76583d",x"715238",x"725238",x"725236",x"745439",x"75563a",x"745439",x"79583c",x"79593d",x"7b5a3e",x"75563c",x"795a3e",x"75553a",x"76583c",x"7a583d",x"7c5b3f",x"7b5b3f",x"805e43",x"856244",x"805e41",x"805f41",x"7e5d40",x"74553a",x"75563a",x"7a593d",x"7e5c41",x"7f5d41",x"78583c",x"775439",x"79583b",x"7a593c",x"785638",x"79583a",x"765436",x"755336",x"735235",x"795637",x"775637",x"765638",x"78573b",x"7c5b3f",x"7d5b3e",x"7b5a3c",x"7d5a3d",x"79583c",x"7c5a3d",x"78583b",x"77573b",x"77583d",x"795a3f",x"7d5c40",x"795a3e",x"79593e",x"77583d",x"77583b",x"77573b",x"745539",x"78593d",x"77583b",x"745538",x"6e4f35",x"715437",x"6f5135",x"654a30",x"6b4d35",x"654930",x"65482f",x"63472d",x"6f5035",x"6a4d34",x"6e4f35",x"644a31",x"674c33",x"684c34",x"6a4e34",x"6a4d34",x"674b33",x"5f452d",x"5e442e",x"5b432d",x"57412c",x"6f5238",x"6c4f36",x"674c34",x"6a4f36",x"74563b",x"74563b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"606060",x"585858",x"505050",x"4f4f4f",x"414141",x"3c3c3c",x"353535",x"333333",x"323232",x"333333",x"333232",x"323232",x"31302f",x"323231",x"333333",x"333333",x"323131",x"323130",x"312f2e",x"333333",x"3e3e3d",x"4f4e4d",x"4f4f4f",x"333333",x"565555",x"474747",x"313131",x"333333",x"333333",x"3c3c3c",x"333333",x"313131",x"000000",x"000000",x"000000",x"5c5c5c",x"535352",x"4a4a49",x"4f4f4f",x"414141",x"434343",x"444444",x"404040",x"3e3e3e",x"464646",x"464646",x"494948",x"343434",x"333333",x"333333",x"323232",x"474747",x"4f4f4f",x"515151",x"474747",x"313131",x"323232",x"323232",x"696561",x"6e6965",x"606060",x"323232",x"333333",x"333333",x"000000",x"635040",x"635040",x"625040",x"624f3f",x"5f5040",x"5d4f3f",x"5e4f3f",x"594b3c",x"5e503f",x"594d3d",x"594d3d",x"4d4135",x"5c4f3f",x"4f4235",x"5b4f3f",x"524637",x"4d4133",x"4f4334",x"564b3c",x"594c3c",x"5d5041",x"504234",x"604c3c",x"644e3e",x"716151",x"564537",x"564738",x"41352a",x"594c3b",x"584c3c",x"5b4b3c",x"614d3e",x"5d4b3b",x"514436",x"4c3f32",x"5c4d3d",x"624e3f",x"5f4f3e",x"635545",x"635040",x"655141",x"695242",x"6a5242",x"665140",x"6a5141",x"634b3d",x"5a4537",x"6c5443",x"655041",x"6b5848",x"675445",x"6c5746",x"6b5848",x"6d5646",x"6a5343",x"6a5444",x"645141",x"685343",x"5e4f3f",x"5f5040",x"665343",x"695443",x"5e5140",x"605242",x"675645",x"645645",x"5f5141",x"5b4f40",x"5b5040",x"604f3f",x"5c5040",x"5b4f3f",x"5d5040",x"624f3f",x"5f5242",x"5e5040",x"5f5343",x"625645",x"4e4235",x"615243",x"685746",x"625343",x"645544",x"675746",x"685645",x"665646",x"5d5141",x"615444",x"615444",x"5a4d3e",x"645443",x"615343",x"625041",x"645041",x"645041",x"655141",x"635141",x"615041",x"604f41",x"5d4f40",x"5d4e3e",x"605142",x"655444",x"615343",x"625545",x"5d5142",x"615444",x"635445",x"625445",x"57483a",x"564a3b",x"5e4f40",x"615343",x"54483a",x"655443",x"4e4133",x"554739",x"544638",x"504336",x"524335",x"554235",x"5f5041",x"645443",x"534335",x"594739",x"544536",x"625241",x"655545",x"655443",x"615141",x"625142",x"605040",x"625342",x"5e5140",x"5c503f",x"5f4c3d",x"574b3c",x"5e4c3c",x"605040",x"5a4d3d",x"605343",x"635645",x"5e5241",x"5a4c3d",x"56493b",x"554839",x"594d3d",x"594d3e",x"655745",x"5d4f40",x"5e5041",x"675343",x"746657",x"5d5041",x"625142",x"605241",x"615444",x"625544",x"625342",x"635242",x"605141",x"554739",x"594c3c",x"5b4e3f",x"231409",x"2c190b",x"361e0d",x"3c210e",x"3f2310",x"412511",x"402410",x"402410",x"3e230f",x"39200e",x"331d0d",x"2a180b",x"221409",x"221409",x"000000",x"000000",x"3c3c3c",x"3c3c3c",x"353535",x"5c5c5c",x"353433",x"343332",x"353230",x"353333",x"373432",x"5d5a59",x"555250",x"3e3a37",x"3e3a37",x"323232",x"343434",x"363535",x"464545",x"353332",x"363433",x"373432",x"343333",x"4a4a4a",x"5f5f5f",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"595858",x"5e5d5b",x"333333",x"323232",x"313131",x"323232",x"323232",x"313131",x"343434",x"323232",x"343434",x"323232",x"4d4d4d",x"505050",x"555555",x"3d3d3d",x"343434",x"323232",x"5b5a5a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"323232",x"333333",x"333333",x"323232",x"5f5f5e",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"000000",x"000000",x"000000",x"000000",x"414141",x"555555",x"5a5a5a",x"585858",x"565656",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"656565",x"585858",x"5f5f5f",x"525252",x"434343",x"323232",x"323232"),
(x"000000",x"2f1a0b",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"4c3627",x"554032",x"573f30",x"563e2e",x"533c2d",x"5d4434",x"5c493b",x"563a28",x"563a28",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"77573a",x"77573a",x"705137",x"725338",x"6e5037",x"6d5037",x"503a26",x"513a27",x"60452f",x"61462e",x"61452e",x"60472f",x"6c4e35",x"6b4e35",x"715339",x"725339",x"6a4d35",x"684c32",x"725339",x"6d5038",x"6c4e36",x"745539",x"6f5036",x"715238",x"75563a",x"7d5c3f",x"79593e",x"7b5b3f",x"795a3e",x"7b5a3e",x"7e5c41",x"815f43",x"7d5b3f",x"805d42",x"7a5a3d",x"78593c",x"815e41",x"816043",x"7c5b3e",x"7d5b3f",x"76573c",x"76573a",x"715136",x"6e4f34",x"735337",x"77563a",x"7a593c",x"755639",x"755436",x"6c4d31",x"765537",x"755538",x"725236",x"745336",x"725134",x"725236",x"775739",x"78573c",x"7f5c40",x"7c5c40",x"805f3f",x"7a593b",x"7a5a3e",x"7b5b3f",x"7c5b3e",x"75573c",x"715439",x"75573b",x"785a3d",x"7c5c40",x"74563a",x"6e5037",x"745437",x"78583a",x"6d4e34",x"6d4e34",x"715236",x"7a5a3b",x"76573a",x"735437",x"755438",x"6b4d32",x"705136",x"644930",x"64482f",x"64472f",x"684a31",x"644931",x"634830",x"6c5036",x"694d34",x"6f5239",x"6b4e36",x"6a4d35",x"6d5038",x"6a4e36",x"644a32",x"644a31",x"553e29",x"6b4e35",x"664b34",x"664b33",x"664a32",x"705237",x"705237",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c4c4c",x"484848",x"3e3e3e",x"393939",x"393939",x"333333",x"323232",x"323131",x"323232",x"323232",x"31302f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5b5a5a",x"52504f",x"585858",x"515151",x"565656",x"505050",x"404040",x"323232",x"333333",x"3b3b3b",x"3c3c3c",x"333333",x"323232",x"323232",x"000000",x"5e5d5d",x"5e5d5d",x"5c5c5c",x"4f4f4f",x"3b3b3b",x"333333",x"323232",x"434343",x"393939",x"3b3b3b",x"3d3d3d",x"454545",x"4a4a4a",x"404040",x"313131",x"313131",x"323232",x"4f4f4f",x"535353",x"434242",x"323232",x"323232",x"323232",x"545454",x"5b5b5b",x"5f5d5c",x"5f5f5f",x"323232",x"323232",x"000000",x"000000",x"5e4f41",x"5e4f41",x"615244",x"544838",x"564839",x"594c3d",x"5b4e3d",x"5b4e3d",x"5f4f3f",x"5e4d3d",x"5c4d3d",x"564838",x"4c4033",x"5f4a3b",x"4c4032",x"564738",x"534536",x"584b3b",x"534738",x"534638",x"4c4032",x"564a3b",x"584c3c",x"584c3d",x"584b3c",x"554839",x"55493a",x"4a3e31",x"594a3a",x"554738",x"574839",x"574738",x"544537",x"5b4b3b",x"5b4a3b",x"524435",x"5b4a3a",x"574838",x"564939",x"564838",x"594a3a",x"574939",x"5e5142",x"594b3c",x"56493a",x"5e4d3d",x"594a3a",x"57483a",x"564a3a",x"5c4e3e",x"625343",x"635645",x"625343",x"675645",x"5f5342",x"625544",x"655544",x"645544",x"675545",x"6a5443",x"675342",x"5c4e3e",x"504133",x"615242",x"635342",x"635443",x"625342",x"5a4a3c",x"514335",x"4d3f32",x"514235",x"5b4c3c",x"5f4e3e",x"594a3b",x"5c4e3e",x"5b493b",x"584d3e",x"614e3f",x"675544",x"625041",x"625141",x"5c4f40",x"615444",x"5f5242",x"625141",x"615443",x"625241",x"685545",x"645141",x"655141",x"665243",x"665243",x"655141",x"645141",x"665343",x"685645",x"675344",x"645343",x"605143",x"645645",x"655443",x"675343",x"655545",x"615545",x"655646",x"655444",x"5f5142",x"625545",x"615241",x"635141",x"675747",x"5e4e40",x"605344",x"56493a",x"625443",x"614e3e",x"655140",x"635040",x"534335",x"4f4133",x"574a3b",x"5d493b",x"554233",x"58493b",x"4e4033",x"4c4032",x"584c3c",x"605241",x"5e5241",x"645746",x"675948",x"5e4e3f",x"625041",x"635241",x"5d4a3b",x"574a3b",x"59493b",x"564739",x"594a3c",x"5c503f",x"5b4e3e",x"594d3d",x"534838",x"594d3c",x"534637",x"5d5140",x"554839",x"544638",x"54483b",x"5b5041",x"5c5141",x"5d5243",x"5a4e40",x"594d3e",x"574b3c",x"584d3d",x"5d4c3d",x"56483b",x"594c3c",x"5e5040",x"615040",x"5e5040",x"5f5040",x"5d5140",x"221308",x"2d180a",x"381f0d",x"3f230f",x"412410",x"422510",x"40230f",x"422510",x"432611",x"3c220f",x"361f0e",x"2c190b",x"241509",x"241509",x"000000",x"000000",x"434343",x"434343",x"5f5f5f",x"2e2e2e",x"616161",x"5a5858",x"4e4d4d",x"4f4d4d",x"5c5a58",x"54514f",x"42403f",x"30302f",x"30302f",x"4f4f4f",x"323232",x"646464",x"575656",x"494747",x"595756",x"595858",x"5f5f5f",x"525252",x"4e4e4e",x"2e2f2f",x"2e2f2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383838",x"323232",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"373737",x"616161",x"5f5e5e",x"585858",x"4b4745",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"333333",x"5b5b5b",x"515151",x"6b6b6b",x"444343",x"000000",x"000000",x"333333",x"333333",x"313131",x"353535",x"4b4b4b",x"474747",x"3f3f3f",x"414141",x"555555",x"5a5a5a",x"585858",x"565656",x"3e3e3e",x"323232",x"323232",x"383838",x"383838",x"000000",x"000000",x"333333",x"606060",x"636363",x"656565",x"585858",x"5f5f5f",x"565656",x"393939",x"323232",x"323232"),
(x"000000",x"351e0d",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301b0c",x"3f2513",x"5f4331",x"5b4230",x"573f2f",x"573e2f",x"5c4435",x"574539",x"523625",x"523625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"7d5c3f",x"7d5c3f",x"7f5f41",x"76563a",x"705035",x"6a4b32",x"60452e",x"654932",x"694d34",x"71543a",x"76573d",x"7d5d41",x"7a593f",x"75553b",x"75563b",x"755539",x"78583d",x"7b5b3e",x"7c5c3f",x"7e5d41",x"7d5d3f",x"836145",x"825f42",x"7b5a3c",x"785738",x"7a593b",x"7f5f43",x"825f45",x"805d41",x"7c5b3f",x"825f42",x"876547",x"866446",x"876447",x"8b6847",x"7d5c3f",x"7d5b3c",x"7d5b3c",x"815e41",x"815e41",x"815e40",x"876445",x"8c6747",x"8a6646",x"825e41",x"876243",x"856040",x"7e5a3d",x"835e3f",x"7b593a",x"7d5b3b",x"7e5c3d",x"815f3f",x"815f41",x"7e5b3b",x"805b3b",x"775636",x"7b5a39",x"856243",x"886446",x"836040",x"7e5c3e",x"856344",x"856244",x"856444",x"866546",x"846445",x"7b5a3d",x"77563a",x"755439",x"79573c",x"7a583c",x"7d5b3f",x"7e5c40",x"856343",x"846144",x"7d5d3d",x"7b5a3b",x"745438",x"7b5a3c",x"7a5a3c",x"78573a",x"7c5a3d",x"7b5a3c",x"715338",x"79593e",x"76563a",x"6e4f34",x"64492d",x"705134",x"6f5237",x"6e5138",x"74553a",x"705236",x"72553a",x"705239",x"72563b",x"6e5138",x"694e35",x"6d4f35",x"6b4c33",x"6b4d34",x"75553a",x"74553a",x"74553a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"393939",x"393939",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"605f5f",x"605f5f",x"5c5c5c",x"505050",x"313131",x"4f4f4f",x"4d4d4d",x"3b3b3b",x"313131",x"434343",x"494949",x"4b4b4b",x"323232",x"313131",x"313131",x"5e5c5a",x"5e5c5a",x"535353",x"434343",x"3c3c3c",x"323232",x"323232",x"474747",x"515151",x"555555",x"4c4c4c",x"434343",x"3d3d3d",x"434343",x"575757",x"3f3f3f",x"333333",x"323232",x"383838",x"363636",x"333333",x"454545",x"3f3f3f",x"484848",x"5b5b5b",x"585858",x"333333",x"343434",x"323232",x"000000",x"000000",x"5f4d3d",x"5f4d3d",x"634d3e",x"614f3f",x"5c4e3d",x"634f3f",x"5f4d3f",x"5d4d3d",x"5c4c3c",x"5c4b3b",x"483a2d",x"5d5141",x"564939",x"544838",x"554839",x"594a3b",x"604c3d",x"5e4b3c",x"5f4b3b",x"614c3c",x"5b493a",x"5a4a3a",x"594939",x"574838",x"534535",x"554838",x"58493a",x"544637",x"584738",x"5a4739",x"5f4a3a",x"614e3f",x"5d4b3b",x"5d4b3b",x"5e4c3d",x"604e3d",x"5e4c3d",x"624f3f",x"665040",x"695141",x"655041",x"644e3f",x"695241",x"685241",x"685343",x"665141",x"625040",x"645141",x"635040",x"5e4f40",x"625141",x"675343",x"665343",x"614e3e",x"645040",x"655443",x"685342",x"695141",x"695242",x"645342",x"5a4c3c",x"615041",x"5b4b3c",x"594a3b",x"5d4f3f",x"5f5141",x"615041",x"5e4e3f",x"635645",x"655847",x"665948",x"615544",x"665847",x"645747",x"645443",x"685646",x"6b5a49",x"6b5949",x"6a5a49",x"5d4f40",x"685746",x"615444",x"635645",x"6b5b4b",x"6b5b4b",x"534639",x"645444",x"685847",x"665443",x"665747",x"635846",x"675847",x"665746",x"5f5142",x"665646",x"645747",x"635747",x"645948",x"574b3c",x"615645",x"645746",x"665645",x"5e5141",x"5d5040",x"615343",x"615443",x"605242",x"615342",x"605442",x"635645",x"635645",x"635645",x"605443",x"5a4f40",x"5d5040",x"5d5141",x"5e5142",x"605344",x"5e5143",x"655444",x"625645",x"645647",x"635343",x"635343",x"635645",x"645847",x"675645",x"665646",x"665645",x"605443",x"615444",x"635645",x"625644",x"645443",x"625040",x"645443",x"625443",x"5e5140",x"584d3d",x"635343",x"5c4e3d",x"584c3c",x"615443",x"5c4f3f",x"5b4e3e",x"644f3f",x"5d4b3c",x"624e3e",x"614d3e",x"655141",x"655241",x"655242",x"675242",x"615141",x"615242",x"5a4c3d",x"5b4c3c",x"5c4d3d",x"5a4c3d",x"5f4f41",x"5a4c3c",x"5f4f3f",x"5e5140",x"5d5140",x"2f1b0c",x"39200f",x"412511",x"402410",x"422410",x"472813",x"4b2b15",x"4a2b15",x"472a14",x"422612",x"3c2310",x"311c0d",x"28170a",x"28170a",x"000000",x"000000",x"575757",x"575757",x"565555",x"323130",x"3b3938",x"3e3d3d",x"484848",x"413f3f",x"3b3430",x"444444",x"4d4d4d",x"353434",x"353434",x"414141",x"696969",x"3c3c3c",x"3f3c3c",x"575656",x"3b3a3a",x"3a3a3a",x"3b3938",x"323232",x"555555",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"444444",x"444444",x"3d3d3d",x"474747",x"000000",x"000000",x"000000",x"000000",x"333333",x"313131",x"323232",x"323232",x"373737",x"616161",x"333333",x"313131",x"313131",x"353535",x"4b4b4b",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"323232",x"484848",x"626262",x"444343",x"333332",x"4a4a4a",x"000000",x"323232",x"313131",x"333333",x"393939",x"444444",x"474747",x"474747",x"636363",x"535353",x"515151",x"313131",x"323232",x"323232",x"323232",x"323232",x"383838",x"383838",x"303131",x"373737",x"2e2f2f",x"3c3d3d",x"626262",x"444444",x"362d27",x"333333",x"554f47",x"333333",x"313131",x"313131"),
(x"000000",x"321c0c",x"321c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"4b3424",x"593d2b",x"563b29",x"5c3f2d",x"5d4332",x"5d4433",x"5e493a",x"4d3220",x"4d3220",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"705137",x"6d4f35",x"64472f",x"63482f",x"5e432d",x"5d432e",x"583f29",x"553e27",x"62462e",x"664930",x"6e4e32",x"6b4d33",x"705134",x"705033",x"704f32",x"6b4d34",x"735336",x"785639",x"795639",x"7c5a3c",x"7d5b3f",x"7b583b",x"785636",x"7c5939",x"715134",x"775836",x"765637",x"7a593b",x"755638",x"755638",x"79583b",x"7f5b3d",x"805d3f",x"7f5d3f",x"7b5a3b",x"805f40",x"78573a",x"7d5b3f",x"79593b",x"745538",x"7b593b",x"77573b",x"75573c",x"705238",x"76563a",x"75573a",x"7a583b",x"78573a",x"7d5b3d",x"815d3d",x"7d5b3e",x"805d40",x"846142",x"835f40",x"7d5a39",x"7f5c3d",x"755539",x"755638",x"78583c",x"77573c",x"78593b",x"79593c",x"7b593d",x"7f5d3f",x"7f5e42",x"815f41",x"7f5d3f",x"7d5d3e",x"755539",x"836042",x"79593d",x"6c4f35",x"78583a",x"77573a",x"755539",x"755537",x"765639",x"78583a",x"6f5136",x"705036",x"79583b",x"7d5a3d",x"745439",x"7d5b3e",x"7c5b3f",x"735338",x"705034",x"745336",x"67492f",x"6a4c30",x"6a4c32",x"6c4d34",x"6f4f34",x"6d4e33",x"715237",x"6a4d34",x"6b4e36",x"60462f",x"5c412a",x"684c32",x"593f29",x"644831",x"4d3623",x"755942",x"755942",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"5a5a5a",x"636363",x"636363",x"343434",x"616161",x"4e4e4e",x"535353",x"5d5d5d",x"565656",x"505050",x"525252",x"323232",x"333333",x"333333",x"585755",x"585755",x"4a4a4a",x"4c4c4c",x"555555",x"323232",x"31302f",x"000000",x"565656",x"545454",x"555555",x"565656",x"575656",x"444444",x"4b4b4b",x"525252",x"585858",x"5b5b5b",x"4a4a4a",x"3b3b3b",x"3f3f3f",x"454545",x"4d4d4d",x"565656",x"666666",x"363636",x"323232",x"323232",x"323333",x"000000",x"000000",x"614d3d",x"614d3d",x"5d4b3c",x"5f4c3d",x"5e4d3e",x"5f4d3e",x"604c3d",x"564939",x"675040",x"534134",x"5b4739",x"5c483a",x"5b493a",x"554336",x"534335",x"584a3a",x"534436",x"5b4a3a",x"5d4a3b",x"5a493a",x"594739",x"534435",x"534434",x"564637",x"544436",x"4d3d31",x"564637",x"594838",x"574939",x"534636",x"574838",x"58493a",x"564939",x"5c4d3c",x"5a4c3c",x"584b3a",x"5e4e3e",x"5d4d3d",x"584939",x"615140",x"645342",x"655342",x"665343",x"645443",x"5f4f3f",x"5e5141",x"5d5140",x"5e5141",x"604f40",x"605040",x"625141",x"604f40",x"645443",x"5f5242",x"5e5141",x"5e5242",x"615545",x"5d5141",x"5b4f40",x"5d4f41",x"594d3f",x"594d3e",x"55493a",x"5f4f40",x"5f4f40",x"645141",x"645140",x"615140",x"5f4f40",x"645645",x"605343",x"645745",x"625645",x"5b4f3f",x"5d5140",x"635444",x"675645",x"685545",x"655343",x"5f4d3e",x"695242",x"615040",x"625141",x"614d3d",x"695443",x"604e3f",x"695444",x"675442",x"645545",x"625544",x"635745",x"655848",x"6d5c4c",x"5f5141",x"665948",x"685b4a",x"645747",x"6a5c4c",x"605343",x"645546",x"655848",x"645645",x"665948",x"655443",x"655443",x"635545",x"655746",x"665948",x"685a49",x"685a49",x"655746",x"615545",x"615544",x"5e5242",x"5e5040",x"5c4c3d",x"5b4e3f",x"5d4e3e",x"5f5241",x"605141",x"605040",x"635343",x"635444",x"625141",x"635645",x"625444",x"615344",x"615544",x"635545",x"645846",x"625645",x"635746",x"645646",x"695343",x"645141",x"665141",x"655141",x"5a4e3f",x"5d4f40",x"5b4e3e",x"615443",x"615243",x"615443",x"5b4c3c",x"5c4f40",x"5a4d3d",x"42362b",x"5a483a",x"5f4b3d",x"5d483a",x"5b483a",x"544537",x"4e4335",x"544436",x"584738",x"5a4a3b",x"5f4f3f",x"5b4b3c",x"5d4e3e",x"5e4e3f",x"5a4d3e",x"635141",x"685242",x"604f3f",x"2c180a",x"371e0d",x"402410",x"432712",x"462812",x"462812",x"442611",x"432611",x"432611",x"3f2410",x"371f0e",x"2b180b",x"24150a",x"24150a",x"000000",x"000000",x"474645",x"474645",x"5b5959",x"3a3532",x"494644",x"3b3735",x"373433",x"393939",x"363636",x"4b4b4b",x"4f4f4f",x"333333",x"333333",x"484848",x"646464",x"323232",x"292a2a",x"38322e",x"4d4d4d",x"444342",x"3a3735",x"4f4f4f",x"525151",x"262727",x"262727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e3e3e",x"333333",x"444444",x"3a3a3a",x"4e4e4e",x"323232",x"323232",x"323232",x"3e3e3e",x"474747",x"4b4b4b",x"4c4c4c",x"373737",x"464646",x"3a3a3a",x"333333",x"313131",x"333333",x"353535",x"4b4b4b",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"494949",x"333333",x"303030",x"343333",x"343333",x"5d5d5d",x"5b5a5a",x"323232",x"323232",x"323232",x"333333",x"434343",x"343333",x"313131",x"323232",x"323232",x"333333",x"303030",x"333333",x"333333",x"32302f",x"313131",x"323232",x"323232",x"323232",x"303131",x"313131",x"323232",x"323232",x"313131",x"313131",x"323232",x"46423e",x"333333",x"313131",x"313131"),
(x"000000",x"2a170b",x"2a170b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"4a3121",x"5f412e",x"674731",x"61412c",x"5b3f2d",x"5b402f",x"584234",x"523522",x"523522",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"694c33",x"694c33",x"664931",x"654931",x"63462d",x"5c432c",x"5b432c",x"5a412b",x"664a30",x"694c32",x"6e4f34",x"6d4e33",x"6e4e34",x"725137",x"745438",x"6d4f36",x"6e5036",x"78573b",x"765639",x"684b31",x"7b593d",x"78573b",x"7d5a3a",x"7c5a3a",x"7c5939",x"7a5839",x"7a593c",x"7e5b3c",x"755538",x"79583a",x"7e5c3e",x"7d5c3f",x"7d5d3e",x"78563a",x"7b5a3d",x"78583b",x"765739",x"77563a",x"78593c",x"76553a",x"7b5b3d",x"77573a",x"78593c",x"73553a",x"735439",x"75543a",x"735538",x"755438",x"76573a",x"815d3f",x"7e5c3e",x"6f4e33",x"7f5c3f",x"7f5c3f",x"805d3e",x"7c5a3d",x"825f3e",x"7e5c3e",x"7c5a3d",x"765739",x"79583a",x"7d5c3e",x"836143",x"846143",x"826042",x"7e5c40",x"78593c",x"7c5b3e",x"78583c",x"79583c",x"7b5c3f",x"75553a",x"7a593c",x"7d5a3d",x"7c5a3d",x"78573b",x"735337",x"755538",x"785739",x"735437",x"715237",x"75553a",x"77563b",x"6b4c32",x"755539",x"7a583c",x"785638",x"785737",x"775536",x"765638",x"705137",x"705136",x"6a4d33",x"725338",x"715339",x"6f5138",x"6a4e36",x"61452f",x"59402a",x"62472f",x"573e29",x"5a402b",x"563d28",x"513925",x"755942",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"5e5d5d",x"3f3f3f",x"343434",x"323232",x"5a5a5a",x"5d5d5d",x"4a4a4a",x"505050",x"565656",x"383838",x"323232",x"323232",x"323232",x"313131",x"000000",x"585757",x"5d5c5c",x"4e4e4e",x"363636",x"323232",x"323232",x"000000",x"000000",x"000000",x"555555",x"575757",x"505050",x"545454",x"5b5b5b",x"4e4e4e",x"4b4b4b",x"4c4c4c",x"4a4a4a",x"585858",x"5e5e5e",x"505050",x"454545",x"353535",x"323232",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"564738",x"564738",x"524535",x"534536",x"504335",x"5a4a3b",x"544738",x"534537",x"514436",x"504335",x"514436",x"5d4a3c",x"564737",x"584537",x"5c473a",x"5f4c3c",x"564638",x"564737",x"564536",x"524334",x"544537",x"564737",x"514133",x"514233",x"574537",x"524335",x"594837",x"5b4939",x"584737",x"5b4839",x"584839",x"584839",x"634f3f",x"5e4e3e",x"604e3d",x"614f3e",x"564839",x"5d4f3f",x"5f5140",x"615342",x"615443",x"615443",x"635443",x"655443",x"665443",x"56493a",x"655141",x"665241",x"655141",x"665141",x"5e4c3d",x"604f3f",x"5f4e3e",x"605140",x"5e5040",x"5c4f3f",x"5a4d3d",x"5a4e3e",x"544738",x"504335",x"5d4f3f",x"5b4f3e",x"534638",x"5b4e3e",x"5d4f3f",x"534738",x"5c4d3d",x"594d3d",x"5e5141",x"5f5141",x"605040",x"5d5040",x"5f503f",x"604e3f",x"5d5241",x"645544",x"655444",x"615343",x"625141",x"645242",x"655242",x"5f5040",x"634f3f",x"645141",x"514235",x"58483a",x"615140",x"615343",x"655645",x"695545",x"655746",x"625645",x"655443",x"5d5140",x"615242",x"645343",x"665544",x"685847",x"655646",x"57483b",x"6a5c4b",x"665847",x"675444",x"695646",x"675343",x"5c4d3f",x"614f3f",x"5d4d3d",x"594d3d",x"524134",x"45372b",x"564336",x"5b4d3d",x"493b2f",x"514335",x"4e4133",x"5e5140",x"5f5240",x"625242",x"615242",x"615243",x"5c4e3f",x"614f3f",x"5a4a3c",x"5f4d3e",x"635445",x"685747",x"675847",x"655444",x"625344",x"625343",x"615343",x"615242",x"655444",x"645243",x"655343",x"675343",x"635545",x"625443",x"635645",x"675847",x"6a5746",x"695444",x"6a5544",x"604e3f",x"604f3f",x"634f3f",x"644f3f",x"624c3d",x"644f40",x"5b4a3b",x"4e4234",x"524537",x"4a3f31",x"594d3c",x"4d4235",x"524638",x"554a3a",x"584d3d",x"5b5040",x"645342",x"5d5141",x"5e503f",x"5b4d3d",x"29170a",x"331c0c",x"381f0d",x"3d220f",x"3e220f",x"3f230f",x"3d210e",x"381d0c",x"351c0b",x"3a200e",x"351e0d",x"27160a",x"201309",x"201309",x"000000",x"000000",x"4f4d4d",x"444241",x"6d6c6c",x"585553",x"54504e",x"5c5a58",x"5e5e5e",x"555555",x"535353",x"535353",x"505050",x"333333",x"333333",x"444444",x"565656",x"4c4c4c",x"333333",x"555555",x"545353",x"565454",x"595755",x"52504e",x"515151",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"3e3e3e",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"474747",x"4b4b4b",x"4c4c4c",x"333333",x"333333",x"333333",x"323232",x"313131",x"313131",x"4e4e4e",x"4d4d4d",x"333333",x"404040",x"404040",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"434343",x"323232",x"302e2d",x"353434",x"343433",x"323131",x"313130",x"626261",x"5a5959",x"656464",x"323232",x"373737",x"656565",x"555453",x"333333",x"343433",x"333333",x"343434",x"323232",x"333333",x"323232",x"454545",x"333333",x"454545",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"333332",x"323232",x"333333",x"46423e",x"514b45",x"323232",x"000000"),
(x"000000",x"361f0e",x"361f0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2e190b",x"523623",x"63442f",x"65422a",x"593c29",x"5b3c2b",x"5a3e2d",x"5b3f2e",x"563824",x"563824",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"694b32",x"694b32",x"664a30",x"654931",x"694c33",x"644830",x"513a25",x"593f29",x"644a31",x"644830",x"6b4c32",x"6b4c33",x"705036",x"705138",x"6c4f36",x"6f5037",x"6e5037",x"73553a",x"745338",x"664b31",x"6b4e34",x"705034",x"7a593a",x"805d41",x"7c5a3d",x"7d5b3d",x"7b5a3d",x"7d5b3d",x"7c5b3e",x"815f43",x"7b5b3e",x"7d5b3d",x"78573a",x"78583c",x"77563a",x"78573a",x"79593b",x"78573a",x"745439",x"705236",x"77573a",x"715237",x"74543a",x"6e5036",x"735439",x"76573b",x"77573b",x"79583b",x"7a593d",x"7a593c",x"7a593d",x"755638",x"735338",x"765537",x"7d5c3f",x"805f42",x"805f41",x"7e5d40",x"805f40",x"805f40",x"816043",x"846345",x"8a6647",x"7c5c40",x"79593d",x"77583d",x"73543a",x"7d5a3f",x"78573c",x"78583d",x"6d4f35",x"6e5036",x"75553a",x"6d5033",x"765538",x"755539",x"765639",x"75563a",x"78583c",x"735237",x"755639",x"765539",x"755539",x"6f5036",x"705137",x"6a4c32",x"705138",x"79593e",x"75573b",x"75553a",x"73553a",x"77573c",x"76563c",x"75573c",x"6e5138",x"705338",x"5f452f",x"5e442f",x"553d28",x"684a33",x"694c32",x"63472f",x"593f29",x"583f28",x"583f28",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"575757",x"3f3f3f",x"343434",x"323232",x"000000",x"545454",x"474747",x"424242",x"3c3c3c",x"333333",x"333232",x"312f2d",x"323232",x"000000",x"000000",x"585757",x"5d5c5c",x"4e4e4e",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"5b5b5b",x"4e4e4e",x"494949",x"484848",x"4a4a4a",x"585858",x"5e5e5e",x"4b4b4b",x"404040",x"383838",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e4b3c",x"5a493a",x"5a4a3a",x"5b4839",x"5d4a3b",x"5a493a",x"5b4a3a",x"5f4b3c",x"574538",x"5b4839",x"594739",x"5b4a3b",x"5a4738",x"554637",x"57493a",x"5a483a",x"5b493a",x"514234",x"534435",x"564537",x"544436",x"524234",x"504133",x"554336",x"584737",x"5d4a3a",x"564536",x"5b4839",x"5e4b3a",x"5c4a3a",x"5c4c3c",x"604e3d",x"5e4e3e",x"5d4e3d",x"5f4e3e",x"5c4d3d",x"62503f",x"645141",x"645241",x"655443",x"665342",x"645443",x"675343",x"635342",x"5e5141",x"655443",x"675343",x"655443",x"655141",x"614d3f",x"635040",x"604f3f",x"635242",x"625141",x"615140",x"5f5040",x"605040",x"59493a",x"544537",x"615141",x"5d4f3f",x"54493a",x"5e5140",x"5a4d3d",x"55493a",x"5a4d3d",x"5b4f3f",x"5f5241",x"5e5141",x"5b4e3e",x"5a4d3d",x"5c4f3f",x"5a4c3d",x"5e5141",x"615343",x"605342",x"5f5141",x"5d5040",x"5f5141",x"5d4f3f",x"5a4e3d",x"5b4e3e",x"5d503f",x"5a4e3e",x"4d4234",x"5d5040",x"605242",x"635645",x"635645",x"645746",x"615544",x"5d5140",x"5d5040",x"5f5242",x"605343",x"655745",x"665545",x"625445",x"5d5141",x"5d5142",x"645747",x"625645",x"645746",x"615444",x"5b4e3f",x"5a4e3d",x"584a3b",x"4e3f31",x"4e4133",x"524637",x"594a3b",x"624e3e",x"5a493b",x"4c3d30",x"4c3d2f",x"524234",x"604f3e",x"625141",x"5d503f",x"534537",x"605343",x"615544",x"615444",x"645646",x"635647",x"645646",x"645242",x"685242",x"6c5142",x"6a5142",x"695243",x"695242",x"6b5342",x"685343",x"605343",x"655746",x"615545",x"645443",x"665444",x"675949",x"645746",x"615545",x"615544",x"5d4f3f",x"564a3b",x"584b3c",x"5d4d3d",x"5b4c3d",x"594a3c",x"574939",x"524436",x"504033",x"574739",x"594c3c",x"54483a",x"55493a",x"534738",x"5a4e3e",x"5d5142",x"635545",x"5d5041",x"605141",x"27170a",x"2b180b",x"341d0d",x"3b210e",x"3e230f",x"412410",x"422510",x"41240f",x"40230f",x"3c210f",x"381f0e",x"301b0c",x"251509",x"251509",x"251509",x"000000",x"000000",x"363433",x"353332",x"393533",x"454240",x"4b4746",x"3d3632",x"31302f",x"323131",x"343332",x"575656",x"606060",x"343434",x"343434",x"424242",x"444444",x"595959",x"5a5a5a",x"525151",x"454343",x"4c4b4a",x"565452",x"514f4f",x"565656",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"3e3d3d",x"434241",x"595959",x"333333",x"343434",x"333333",x"353535",x"323232",x"323232",x"323232",x"333333",x"333231",x"313131",x"333333",x"313131",x"323232",x"333333",x"333333",x"343434",x"323232",x"505050",x"333333",x"404040",x"404040",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333232",x"353434",x"333232",x"333232",x"333333",x"323232",x"353332",x"383736",x"5b5a59",x"67625d",x"413e3c",x"636262",x"666564",x"5e5d5c",x"595858",x"414141",x"505050",x"3b3b3b",x"343434",x"313131",x"323232",x"545454",x"3e3e3e",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"371f0f",x"371f0f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2b190b",x"4a3323",x"60412d",x"5c3e29",x"5c3e2a",x"5c3d28",x"65432d",x"5f4432",x"553823",x"553823",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"6c5136",x"6c5136",x"6e5036",x"6c5036",x"6d5038",x"5f472f",x"5a422c",x"614730",x"6f5337",x"6d4f35",x"6f5137",x"72553a",x"715439",x"705138",x"725338",x"79593d",x"6f5037",x"78583c",x"76563b",x"705136",x"77563c",x"7b593c",x"7b593c",x"7c5a3c",x"775638",x"755538",x"755539",x"725136",x"735337",x"78573a",x"79583b",x"6f4e36",x"725436",x"77573b",x"7c5a3e",x"7d5d3f",x"7d5c40",x"7f5f40",x"78573c",x"795a3d",x"7f5f41",x"7b5b3e",x"7a5a3c",x"785a3e",x"795a3e",x"7b5b40",x"7b5a3d",x"805d3f",x"76563b",x"7f5e3f",x"7e5d3f",x"77573a",x"7d5c3e",x"79593c",x"7a583b",x"7d5c3e",x"78583b",x"73533a",x"775639",x"7a583a",x"79593b",x"7c5a3e",x"7d5c3f",x"735339",x"715438",x"73553b",x"805e42",x"7d5d40",x"816146",x"795b40",x"7d5d42",x"805f43",x"816043",x"7c5b3e",x"715337",x"836141",x"7c5b3e",x"78583c",x"77563a",x"7c5b3d",x"7b593b",x"7b5b3d",x"78573a",x"76573a",x"79593d",x"75563a",x"75553a",x"715237",x"715237",x"6f4f35",x"684b32",x"6e4e34",x"6b4c34",x"6c4d34",x"6d5037",x"61462f",x"5d432d",x"5e442f",x"59402b",x"624931",x"6c4f37",x"6b4e35",x"61472f",x"60462e",x"6c4e34",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"464646",x"424242",x"3c3c3c",x"333333",x"333333",x"333232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b4b4b",x"404040",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a493a",x"5a4a3a",x"5b4839",x"5d4a3b",x"5a493a",x"5b4a3a",x"5f4b3c",x"574538",x"5b4839",x"594739",x"5b4a3b",x"5a4738",x"554637",x"57493a",x"5a483a",x"5b493a",x"514234",x"534435",x"564537",x"544436",x"524234",x"504133",x"554336",x"584737",x"5d4a3a",x"564536",x"5b4839",x"5e4b3a",x"5c4a3a",x"5c4c3c",x"604e3d",x"5e4e3e",x"5d4e3d",x"5f4e3e",x"5c4d3d",x"62503f",x"645141",x"645241",x"655443",x"665342",x"645443",x"675343",x"635342",x"5e5141",x"655443",x"675343",x"655443",x"655141",x"614d3f",x"635040",x"604f3f",x"635242",x"625141",x"615140",x"5f5040",x"605040",x"59493a",x"544537",x"615141",x"5d4f3f",x"54493a",x"5e5140",x"5a4d3d",x"55493a",x"5a4d3d",x"5b4f3f",x"5f5241",x"5e5141",x"5b4e3e",x"5a4d3d",x"5c4f3f",x"5a4c3d",x"5e5141",x"615343",x"605342",x"5f5141",x"5d5040",x"5f5141",x"5d4f3f",x"5a4e3d",x"5b4e3e",x"5d503f",x"5a4e3e",x"4d4234",x"5d5040",x"605242",x"635645",x"635645",x"645746",x"615544",x"5d5140",x"5d5040",x"5f5242",x"605343",x"655745",x"665545",x"625445",x"5d5141",x"5d5142",x"645747",x"625645",x"645746",x"615444",x"5b4e3f",x"5a4e3d",x"584a3b",x"4e3f31",x"4e4133",x"524637",x"594a3b",x"624e3e",x"5a493b",x"4c3d30",x"4c3d2f",x"524234",x"604f3e",x"625141",x"5d503f",x"534537",x"605343",x"615544",x"615444",x"645646",x"635647",x"645646",x"645242",x"685242",x"6c5142",x"6a5142",x"695243",x"695242",x"6b5342",x"685343",x"605343",x"655746",x"615545",x"645443",x"665444",x"675949",x"645746",x"615545",x"615544",x"5d4f3f",x"564a3b",x"584b3c",x"5d4d3d",x"5b4c3d",x"594a3c",x"574939",x"524436",x"504033",x"574739",x"594c3c",x"54483a",x"55493a",x"534738",x"5a4e3e",x"5d5142",x"635545",x"5d5041",x"241509",x"241509",x"28170a",x"301b0c",x"371e0d",x"3c220f",x"3c210e",x"3d210f",x"3d220f",x"3f2410",x"3c220f",x"351e0d",x"28160a",x"1f1208",x"221409",x"221409",x"000000",x"000000",x"000000",x"363433",x"3b3634",x"454240",x"4e4b49",x"373533",x"31302f",x"323131",x"5a5a5a",x"504e4e",x"3a3938",x"575656",x"575656",x"444444",x"3c3c3c",x"333333",x"372e2a",x"333332",x"3b3a39",x"353433",x"332d28",x"4a4a4a",x"333333",x"3f3f3f",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333232",x"313131",x"323232",x"404040",x"333333",x"333333",x"323232",x"313131",x"353535",x"343434",x"323232",x"313131",x"313131",x"332c29",x"323232",x"434343",x"484848",x"323232",x"333333",x"323232",x"343434",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323131",x"323232",x"343333",x"343433",x"363433",x"373636",x"383331",x"59514a",x"383432",x"3a3533",x"373331",x"343231",x"333130",x"343434",x"313131",x"313131",x"323232",x"323232",x"323232",x"4b4a4a",x"5b5b5b",x"333333",x"323232",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"3a210f",x"3a210f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1a0c",x"422919",x"5e412e",x"62432d",x"6a4831",x"5f412d",x"654731",x"564031",x"51331f",x"51331f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"715238",x"715238",x"6d4f35",x"6e5036",x"61472e",x"61462f",x"5b422b",x"62472f",x"654931",x"6b4c33",x"6e4e35",x"674b31",x"6a4c32",x"694a31",x"6f5035",x"705137",x"6f5037",x"74543a",x"7b5b3e",x"7f5c40",x"7c5a3e",x"7e5c3e",x"7e593b",x"805d3e",x"815f40",x"7e5c3d",x"805e3e",x"735237",x"78573a",x"755538",x"7d5c3d",x"836143",x"7d5c3f",x"7d5c3e",x"7f5d3f",x"805e40",x"7b5a3b",x"78573b",x"79593b",x"7a593c",x"78573b",x"78583b",x"79593c",x"725438",x"715237",x"715138",x"755439",x"76583b",x"76573a",x"7c5a3d",x"7f5e41",x"805e41",x"825f42",x"815e40",x"79573b",x"7e5d3e",x"805f40",x"7e5d3f",x"805f3f",x"765439",x"7d5c3d",x"78573a",x"7e5e40",x"846345",x"836143",x"826042",x"815d41",x"7f5e41",x"7d5c3f",x"78573b",x"7d5c3f",x"7d5a3d",x"785639",x"7b583a",x"755539",x"705136",x"715235",x"735335",x"755538",x"775639",x"755438",x"7d593b",x"7a5a3c",x"7a583d",x"77563b",x"7d5c3e",x"775539",x"775639",x"78573b",x"75563a",x"6e5036",x"684b32",x"705036",x"684b32",x"6e5138",x"78593f",x"6a4f36",x"664b32",x"58402b",x"6c4f36",x"6a4d33",x"64482f",x"62472e",x"6a4d33",x"6a4d33",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25190f",x"25190f",x"24180f",x"2a190e",x"2e1b0e",x"25170e",x"2b1b0f",x"2c1a0d",x"2f1c0e",x"351e0e",x"331d0d",x"2b190b",x"2a170a",x"27160a",x"29170a",x"2d1a0b",x"301b0b",x"2e190b",x"2d190b",x"28160a",x"29170a",x"27160a",x"28170a",x"29170a",x"28170a",x"2b180b",x"311c0d",x"341d0d",x"28160a",x"261509",x"29170a",x"2d1a0b",x"2e1a0b",x"2d190b",x"2c180b",x"2e1a0b",x"2c190b",x"2d1a0b",x"2b190b",x"29170a",x"241509",x"271709",x"2a180b",x"27160a",x"25160a",x"231409",x"26160a",x"231409",x"23150a",x"25150a",x"24150a",x"26160a",x"28170b",x"2a180b",x"2e1a0c",x"27170b",x"2a180b",x"2a180a",x"29170a",x"26160a",x"28170a",x"231409",x"221409",x"231409",x"24150a",x"27170a",x"28170a",x"28170a",x"28160a",x"27170a",x"26160a",x"26150a",x"25150a",x"241509",x"221509",x"27160a",x"221409",x"251509",x"24150a",x"28170a",x"27160a",x"2c1a0a",x"26170a",x"231509",x"221409",x"1f1209",x"241509",x"231409",x"1a1008",x"1a1008",x"301a0b",x"341d0c",x"2e1a0b",x"26160a",x"2a180a",x"301b0b",x"2b180a",x"2d1a0a",x"2d190b",x"2d190b",x"25150a",x"160e07",x"160f07",x"170f07",x"180f08",x"191008",x"1e1309",x"27180a",x"221509",x"271709",x"291909",x"281909",x"2b1a0b",x"221408",x"261709",x"241509",x"221509",x"241609",x"2a1a0a",x"201308",x"1e1208",x"201208",x"211309",x"221409",x"231409",x"211409",x"211309",x"221409",x"221409",x"221409",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"201308",x"201309",x"201309",x"201309",x"201309",x"221409",x"23150a",x"201309",x"211409",x"221309",x"23150a",x"221409",x"221409",x"221409",x"221409",x"23150a",x"231409",x"231509",x"241509",x"231409",x"25150a",x"231409",x"221409",x"231409",x"241409",x"201309",x"211309",x"1f1208",x"201208",x"201309",x"201309",x"201309",x"211409",x"201309",x"211309",x"1f1309",x"201309",x"1f1309",x"1f1309",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"191008",x"190f08",x"190f08",x"1b1108",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"1b1108",x"1c1108",x"1f1408",x"201408",x"201308",x"211409",x"211409",x"211409",x"201409",x"261709",x"2d1c0a",x"38230c",x"472a10",x"472a10",x"000000",x"000000",x"000000",x"1f1208",x"1f1208",x"221409",x"2b180b",x"311b0c",x"381f0e",x"381f0e",x"39200e",x"3a200e",x"38200e",x"331d0d",x"2b190b",x"231509",x"1a1008",x"28170a",x"28170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5b5a5a",x"504e4e",x"3a3938",x"575656",x"000000",x"000000",x"000000",x"323232",x"372e2a",x"333332",x"3b3a39",x"353433",x"332d28",x"333333",x"333333",x"3f3f3f",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333231",x"323232",x"333333",x"323232",x"333333",x"333333",x"424242",x"323232",x"333333",x"383838",x"525252",x"5f5f5f",x"393939",x"515151",x"545454",x"323232",x"333333",x"323232",x"3a3a3a",x"313131",x"313131",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343333",x"333231",x"363433",x"373636",x"3a3634",x"554d46",x"393532",x"383533",x"383533",x"36302d",x"353332",x"333333",x"323232",x"323232",x"313131",x"323232",x"323232",x"4b4a4a",x"5b5b5b",x"3c3c3c",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"331d0d",x"331d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"4c382a",x"594131",x"553e30",x"5c4232",x"5c4231",x"624634",x"504033",x"543725",x"543725",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"73553b",x"73553b",x"76573c",x"886951",x"85664b",x"7c6049",x"795d45",x"7f6149",x"8c6d54",x"85654b",x"85664c",x"88694e",x"89694c",x"88694d",x"816147",x"816145",x"836248",x"816045",x"846348",x"87664a",x"8a694c",x"8b694d",x"866448",x"8c6a4c",x"8c6949",x"8b694a",x"8a684a",x"866447",x"846345",x"815f43",x"826043",x"836143",x"856346",x"856346",x"856347",x"856245",x"896649",x"836143",x"846245",x"846143",x"846144",x"886546",x"826042",x"836244",x"866345",x"856345",x"856244",x"846143",x"846244",x"886445",x"896545",x"8d6a4b",x"8e6a4b",x"886445",x"846144",x"866243",x"876446",x"866346",x"846244",x"8a6648",x"886446",x"8b6849",x"8a6748",x"8c694b",x"926e50",x"8d6a4c",x"8d6b4c",x"89674a",x"856448",x"846348",x"836246",x"866649",x"896549",x"876547",x"88684b",x"856346",x"8b694a",x"8b694c",x"886649",x"8a674a",x"856346",x"8a694b",x"8a694e",x"89684b",x"8f6d50",x"89694e",x"85654a",x"88694e",x"86664b",x"88694f",x"816348",x"846448",x"8e6d51",x"806147",x"806147",x"826349",x"7d5f46",x"81634a",x"745a44",x"82644b",x"82664d",x"7e6148",x"7b624d",x"795d44",x"795d44",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"25190f",x"25190f",x"24180f",x"2a190e",x"2e1b0e",x"25170e",x"2b1b0f",x"2c1a0d",x"2f1c0e",x"351e0e",x"331d0d",x"2b190b",x"2a170a",x"27160a",x"29170a",x"2d1a0b",x"301b0b",x"2e190b",x"2d190b",x"28160a",x"29170a",x"27160a",x"28170a",x"29170a",x"28170a",x"2b180b",x"311c0d",x"341d0d",x"28160a",x"261509",x"29170a",x"2d1a0b",x"2e1a0b",x"2d190b",x"2c180b",x"2e1a0b",x"2c190b",x"2d1a0b",x"2b190b",x"29170a",x"241509",x"271709",x"2a180b",x"27160a",x"25160a",x"231409",x"26160a",x"231409",x"23150a",x"25150a",x"24150a",x"26160a",x"28170b",x"2a180b",x"2e1a0c",x"27170b",x"2a180b",x"2a180a",x"29170a",x"26160a",x"28170a",x"231409",x"221409",x"231409",x"24150a",x"27170a",x"28170a",x"28170a",x"28160a",x"27170a",x"26160a",x"26150a",x"25150a",x"241509",x"221509",x"27160a",x"221409",x"251509",x"24150a",x"28170a",x"27160a",x"2c1a0a",x"26170a",x"231509",x"221409",x"1f1209",x"241509",x"231409",x"1a1008",x"1a1008",x"301a0b",x"341d0c",x"2e1a0b",x"26160a",x"2a180a",x"301b0b",x"2b180a",x"2d1a0a",x"2d190b",x"2d190b",x"25150a",x"160e07",x"160f07",x"170f07",x"180f08",x"191008",x"1e1309",x"27180a",x"221509",x"271709",x"291909",x"281909",x"2b1a0b",x"221408",x"261709",x"241509",x"221509",x"241609",x"2a1a0a",x"201308",x"1e1208",x"201208",x"211309",x"221409",x"231409",x"211409",x"211309",x"221409",x"221409",x"221409",x"201309",x"201309",x"1f1208",x"1f1208",x"1e1208",x"201308",x"201309",x"201309",x"201309",x"201309",x"221409",x"23150a",x"201309",x"211409",x"221309",x"23150a",x"221409",x"221409",x"221409",x"221409",x"23150a",x"231409",x"231509",x"241509",x"231409",x"25150a",x"231409",x"221409",x"231409",x"241409",x"201309",x"211309",x"1f1208",x"201208",x"201309",x"201309",x"201309",x"211409",x"201309",x"211309",x"1f1309",x"201309",x"1f1309",x"1f1309",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"191008",x"190f08",x"190f08",x"1b1108",x"170f07",x"170f07",x"160f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"160e07",x"160e07",x"160e07",x"160f07",x"170f07",x"1b1108",x"1c1108",x"1f1408",x"201408",x"201308",x"211409",x"211409",x"211409",x"201409",x"261709",x"2d1c0a",x"38230c",x"472a10",x"472a10",x"000000",x"000000",x"000000",x"37200e",x"37200e",x"452912",x"482a13",x"482913",x"462912",x"472913",x"4a2b14",x"482a12",x"4b2c14",x"4a2b14",x"4b2c14",x"4c2d14",x"4c2d15",x"432511",x"432511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"323131",x"303030",x"606060",x"333333",x"333333",x"333333",x"323232",x"333333",x"585858",x"474544",x"494949",x"323232",x"333232",x"323232",x"373636",x"313131",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a3634",x"554d46",x"393532",x"383533",x"383533",x"36302d",x"353332",x"333333",x"323232",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"351f0f",x"351f0f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0c",x"463123",x"5f493a",x"5f4738",x"594132",x"5d4230",x"594132",x"4b3c31",x"513623",x"513623",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"73553b",x"73553b",x"76573c",x"886951",x"85664b",x"7c6049",x"795d45",x"7f6149",x"8c6d54",x"85654b",x"85664c",x"88694e",x"89694c",x"88694d",x"816147",x"816145",x"836248",x"816045",x"846348",x"87664a",x"8a694c",x"8b694d",x"866448",x"8c6a4c",x"8c6949",x"8b694a",x"8a684a",x"866447",x"846345",x"815f43",x"826043",x"836143",x"856346",x"856346",x"856347",x"856245",x"896649",x"836143",x"846245",x"846143",x"846144",x"886546",x"826042",x"836244",x"866345",x"856345",x"856244",x"846143",x"846244",x"886445",x"896545",x"8d6a4b",x"8e6a4b",x"886445",x"846144",x"866243",x"876446",x"866346",x"846244",x"8a6648",x"886446",x"8b6849",x"8a6748",x"8c694b",x"926e50",x"8d6a4c",x"8d6b4c",x"89674a",x"856448",x"846348",x"836246",x"866649",x"896549",x"876547",x"88684b",x"856346",x"8b694a",x"8b694c",x"886649",x"8a674a",x"856346",x"8a694b",x"8a694e",x"89684b",x"8f6d50",x"89694e",x"85654a",x"88694e",x"86664b",x"88694f",x"816348",x"846448",x"8e6d51",x"806147",x"806147",x"826349",x"7d5f46",x"81634a",x"745a44",x"82644b",x"82664d",x"7e6148",x"7b624d",x"795d44",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"23180f",x"23180f",x"1f160f",x"1e160f",x"1e140d",x"22160d",x"20160d",x"20140b",x"21150b",x"241509",x"231409",x"1f1208",x"1f1208",x"201309",x"221409",x"221409",x"201208",x"201208",x"1d1108",x"1e1108",x"1d1108",x"201308",x"231409",x"211409",x"201309",x"1f1208",x"1c1108",x"1d1108",x"1c1108",x"1e1208",x"211409",x"28170a",x"2b1a09",x"291809",x"281809",x"231508",x"221409",x"211309",x"201309",x"201309",x"211408",x"271809",x"251609",x"1f1308",x"1e1208",x"1e1208",x"1f1209",x"1f1209",x"1f1309",x"1f1208",x"1f1209",x"1f1309",x"201309",x"211309",x"211409",x"211409",x"211409",x"211409",x"211409",x"201309",x"201309",x"201309",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"190f08",x"170f07",x"160e07",x"150e07",x"150e07",x"241508",x"301c0b",x"271609",x"2c1a0a",x"2d190b",x"2a170a",x"2d190a",x"2d190b",x"2b180b",x"2e1a0b",x"2d190b",x"2d190b",x"2e1a0b",x"301b0c",x"28160a",x"261509",x"251509",x"28160a",x"241509",x"2b180b",x"160e07",x"160e07",x"160f07",x"170f07",x"180f07",x"190f07",x"1c1208",x"221509",x"1f1308",x"231509",x"241609",x"281809",x"221509",x"1f1308",x"261709",x"211409",x"221409",x"1f1308",x"231509",x"1e1108",x"1c1108",x"1e1108",x"1f1208",x"211309",x"231409",x"231509",x"231509",x"231409",x"221409",x"211309",x"201208",x"201208",x"211309",x"1f1208",x"1d1108",x"1d1108",x"1c1108",x"1d1108",x"201309",x"211309",x"221409",x"231509",x"221409",x"24150a",x"221409",x"221409",x"221409",x"221409",x"231509",x"231509",x"24150a",x"231409",x"231409",x"231409",x"231409",x"231409",x"221409",x"221409",x"221409",x"221409",x"221409",x"211309",x"211309",x"211409",x"211309",x"201309",x"201309",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"1d1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"180f07",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"160f07",x"160e07",x"170f07",x"180f07",x"1a1108",x"1c1108",x"1f1308",x"1f1308",x"201308",x"201408",x"1f1308",x"1c1208",x"1d1108",x"1f1308",x"2c1c09",x"35210b",x"3d250d",x"3e260d",x"3e260d",x"000000",x"000000",x"37200e",x"37200e",x"452912",x"482a13",x"482913",x"462912",x"472913",x"4a2b14",x"482a12",x"4b2c14",x"4a2b14",x"4b2c14",x"4c2d14",x"4c2d15",x"432511",x"432511",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"313131",x"5d5d5d",x"323232",x"323232",x"323231",x"333333",x"323232",x"343535",x"3e3b38",x"404040",x"363636",x"323232",x"333232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"351e0d",x"351e0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29170a",x"543c2c",x"5f4839",x"5d4333",x"593e2c",x"5a402e",x"4f3929",x"4a3a2e",x"513421",x"513421",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"271a0f",x"271a0f",x"21170f",x"1f170f",x"291c12",x"29190e",x"20160c",x"22160d",x"20140b",x"201308",x"201208",x"27160a",x"2a180b",x"241509",x"26170a",x"261609",x"261609",x"231409",x"201309",x"1f1208",x"241509",x"211408",x"231508",x"251609",x"231508",x"1f1208",x"1e1108",x"1d1108",x"1e1208",x"201308",x"27170a",x"2e1c0b",x"341f0b",x"301c0b",x"27170a",x"251509",x"241509",x"231509",x"221408",x"211408",x"28190a",x"27170a",x"231409",x"201308",x"1f1208",x"201309",x"201309",x"201309",x"1f1209",x"1f1309",x"201409",x"201309",x"201309",x"211309",x"211409",x"221409",x"231409",x"24150a",x"24150a",x"23150a",x"221409",x"211409",x"211409",x"201309",x"201309",x"201309",x"1f1309",x"201309",x"1f1309",x"1f1309",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"1a1008",x"191008",x"170f07",x"170f07",x"160e07",x"150e07",x"2b1a0a",x"341e0d",x"351f0d",x"331e0c",x"311c0c",x"2f1c0c",x"2d1a0b",x"2e1a0b",x"2f1b0c",x"331d0d",x"2c180b",x"2d190b",x"2f1a0b",x"331d0d",x"311b0c",x"2c190b",x"2b190b",x"29170a",x"28170a",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"190f08",x"1a1008",x"1c1108",x"1c1108",x"1d1108",x"1f1308",x"1f1208",x"221408",x"1e1208",x"1f1208",x"1e1208",x"201209",x"1f1208",x"201208",x"211409",x"221309",x"211309",x"201308",x"201308",x"211308",x"221309",x"221409",x"221409",x"221309",x"211309",x"211309",x"211308",x"221409",x"201309",x"201308",x"201208",x"1f1208",x"1f1208",x"1f1208",x"201309",x"201309",x"201308",x"221409",x"221409",x"25160a",x"25150a",x"241509",x"241509",x"241509",x"25150a",x"26160a",x"25150a",x"241509",x"26160a",x"25160a",x"241509",x"241509",x"231409",x"241509",x"24150a",x"25160a",x"26160a",x"25160a",x"25150a",x"24150a",x"24150a",x"24150a",x"231509",x"231409",x"221409",x"221409",x"211409",x"221409",x"211309",x"201309",x"201309",x"1f1208",x"1e1208",x"1d1208",x"1c1108",x"1b1108",x"1a1008",x"191008",x"180f07",x"180f08",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"190f08",x"1b1008",x"1d1208",x"1f1308",x"1e1208",x"1f1308",x"1f1308",x"1f1308",x"1e1308",x"1c1108",x"1b1107",x"281a09",x"33200a",x"38220c",x"39220c",x"39220c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"313131",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"2e2e2e",x"313131",x"2c2c2c",x"323232",x"313131",x"5d5d5d",x"333333",x"323232",x"333333",x"333333",x"323232",x"343535",x"44403d",x"393837",x"3b3b3b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"2f2f2f",x"323232",x"323232",x"333333",x"323232",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"341e0e",x"341e0e",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"574030",x"624d3e",x"5d4737",x"5a4333",x"573f2f",x"563f30",x"4e3e32",x"553622",x"553622",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e4136",x"483d34",x"5d4736",x"624b39",x"67513f",x"69513e",x"695240",x"695340",x"655140",x"695240",x"69523e",x"785c45",x"6b543f",x"6c5440",x"67513e",x"644e3d",x"644f3d",x"664f3d",x"624c3b",x"66513f",x"67503e",x"69513d",x"765941",x"634b38",x"664e3a",x"634d3a",x"5e4a38",x"644d39",x"6e523b",x"604936",x"684e39",x"674e3a",x"6b523d",x"745741",x"715641",x"715743",x"6e5540",x"6b5340",x"6b5441",x"6b5544",x"685443",x"705844",x"6f5743",x"735640",x"6c513a",x"604935",x"624935",x"56412e",x"553f2d",x"604833",x"58412f",x"4b3829",x"533d2b",x"58402d",x"5e4732",x"6d5139",x"654a35",x"5a4331",x"614a36",x"5f4734",x"674e39",x"604b38",x"5c4939",x"65503e",x"6c533e",x"67513f",x"6c513b",x"654e3b",x"69503c",x"624c3a",x"66503e",x"6b523f",x"6a523e",x"674f3b",x"6e5643",x"6f5642",x"6b5442",x"735741",x"6a5240",x"6e5643",x"695241",x"745a45",x"765b46",x"6e5644",x"715a47",x"745c47",x"6f5845",x"635141",x"000000",x"000000",x"000000",x"291a11",x"291a11",x"23180f",x"1f160f",x"2a1f17",x"20150d",x"22160d",x"23160d",x"26170b",x"231309",x"231409",x"29170a",x"221409",x"2a180a",x"2a180b",x"29170a",x"2a180a",x"27160a",x"27160a",x"211409",x"29160a",x"271609",x"271609",x"211309",x"271509",x"241409",x"201308",x"231409",x"211309",x"2d1a0b",x"2b180a",x"331d0b",x"311d0b",x"331e0b",x"2d190b",x"2a170a",x"27160a",x"241509",x"221409",x"231509",x"231508",x"231509",x"1e1208",x"201309",x"1f1309",x"1f1209",x"241509",x"2d190b",x"27160a",x"2b180b",x"2d190b",x"2f1b0c",x"321d0d",x"301b0c",x"311c0c",x"321c0d",x"331d0d",x"2f1b0c",x"301b0c",x"301b0c",x"2f1a0b",x"2f1a0b",x"2f1b0c",x"321c0d",x"311c0c",x"2e190b",x"2d190b",x"2d1a0b",x"2f1a0b",x"301b0c",x"2c190a",x"331e0c",x"2e1b0b",x"311c0c",x"2c190b",x"2f1b0c",x"2d190b",x"331d0d",x"2e1a0c",x"331d0d",x"311c0c",x"331d0c",x"301b0c",x"321c0c",x"2f1a0b",x"2c190b",x"301b0c",x"301c0c",x"341e0d",x"311c0d",x"2d190b",x"301a0b",x"2c190b",x"301b0c",x"2a180b",x"301b0c",x"311b0c",x"301b0c",x"2f1a0b",x"311c0c",x"331c0c",x"301b0c",x"2b180a",x"2a170a",x"261609",x"1b1008",x"1c1108",x"1d1108",x"1d1108",x"201308",x"221409",x"241409",x"201308",x"251509",x"2a180a",x"28170a",x"26160a",x"2a180a",x"2b180b",x"2c190b",x"2c190b",x"2d190b",x"29170a",x"281609",x"271609",x"29170a",x"281609",x"271509",x"28160a",x"271609",x"2c190b",x"2b190b",x"2a170a",x"29170a",x"29170a",x"2b180a",x"2c180a",x"2b180a",x"2b180a",x"2b180a",x"2c190b",x"2e1a0b",x"2f1b0c",x"331d0d",x"2c180b",x"2d190b",x"2d190b",x"2e1a0c",x"301b0c",x"2f1b0c",x"2d190b",x"2d190b",x"2c190b",x"2f1b0c",x"2e1b0c",x"2e1b0c",x"2b190b",x"2e1a0b",x"2f1b0c",x"301c0c",x"2f1b0c",x"2c190b",x"2b180a",x"2b170a",x"2d190b",x"2d190b",x"2b190b",x"2c190b",x"29170a",x"2c190b",x"2c190b",x"2e1a0b",x"29170a",x"2b180b",x"2a180b",x"2b190b",x"2a170a",x"2b180b",x"2a180b",x"28170a",x"28170a",x"26160a",x"231409",x"2d190b",x"2c190b",x"2c190b",x"2d190b",x"2b180b",x"2e1a0b",x"2f1b0c",x"301c0d",x"351e0e",x"301b0c",x"2b180b",x"2c190b",x"2d190b",x"321c0d",x"2f1b0c",x"1a1008",x"1a1008",x"1b1008",x"1c1108",x"1f1308",x"221409",x"231409",x"251509",x"241509",x"28160a",x"201308",x"281609",x"2d1b0a",x"2f1c0a",x"221508",x"201308",x"201308",x"000000",x"000000",x"000000",x"000000",x"515151",x"313131",x"333333",x"484848",x"333333",x"313131",x"343434",x"373737",x"383838",x"323232",x"323232",x"313131",x"313131",x"313131",x"323232",x"333333",x"323232",x"323232",x"333333",x"373737",x"444444",x"494949",x"484848",x"484848",x"424242",x"3c3c3c",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"313131",x"333333",x"323232",x"333232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f3030",x"303030",x"323232",x"313131",x"2e2e2e",x"313131",x"2c2c2c",x"323232",x"2b2b2b",x"323232",x"303030",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"313131",x"282828",x"313131",x"323232",x"323232",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"331d0d",x"331d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1b0c",x"625144",x"5f4c3d",x"5d4a3d",x"5c483a",x"5c4738",x"604b3c",x"4e4237",x"543d2d",x"543d2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e321f",x"4e321f",x"4e4136",x"483d34",x"5d4736",x"624b39",x"67513f",x"69513e",x"695240",x"695340",x"655140",x"695240",x"69523e",x"785c45",x"6b543f",x"6c5440",x"67513e",x"644e3d",x"644f3d",x"664f3d",x"624c3b",x"66513f",x"67503e",x"69513d",x"765941",x"634b38",x"664e3a",x"634d3a",x"5e4a38",x"644d39",x"6e523b",x"604936",x"684e39",x"674e3a",x"6b523d",x"745741",x"715641",x"715743",x"6e5540",x"6b5340",x"6b5441",x"6b5544",x"685443",x"705844",x"6f5743",x"735640",x"6c513a",x"604935",x"624935",x"56412e",x"553f2d",x"604833",x"58412f",x"4b3829",x"533d2b",x"58402d",x"5e4732",x"6d5139",x"654a35",x"5a4331",x"614a36",x"5f4734",x"674e39",x"604b38",x"5c4939",x"65503e",x"6c533e",x"67513f",x"6c513b",x"654e3b",x"69503c",x"624c3a",x"66503e",x"6b523f",x"6a523e",x"674f3b",x"6e5643",x"6f5642",x"6b5442",x"735741",x"6a5240",x"6e5643",x"695241",x"745a45",x"765b46",x"6e5644",x"715a47",x"745c47",x"6f5845",x"635141",x"634e3d",x"634e3d",x"000000",x"2f1e13",x"2f1e13",x"271b11",x"271e17",x"261a10",x"291a0f",x"24160d",x"28180d",x"26170b",x"2a180b",x"29160a",x"251409",x"231409",x"251509",x"2a170a",x"2c190b",x"2d190b",x"2a180b",x"301b0c",x"2e1a0b",x"27170a",x"241509",x"2c180b",x"29170a",x"271609",x"271509",x"261509",x"2a170a",x"2b180b",x"241509",x"261609",x"2b180a",x"2d190a",x"2d190a",x"2b180a",x"2c190a",x"29170a",x"231509",x"201309",x"1f1208",x"1d1108",x"1d1108",x"1e1208",x"211409",x"1f1309",x"1f1209",x"211309",x"25150a",x"27160a",x"2c190b",x"2e1a0c",x"2c190b",x"331d0d",x"361f0e",x"311c0d",x"331d0d",x"331d0d",x"2d1a0b",x"301b0c",x"301b0c",x"2f1b0c",x"2f1a0c",x"311b0c",x"2f1b0c",x"2e1a0b",x"2d190b",x"301b0c",x"2f1b0c",x"2e1a0c",x"301b0c",x"301b0b",x"2e1a0b",x"301b0b",x"2e1a0b",x"2f1c0c",x"301b0c",x"2a180b",x"2c190b",x"2a180b",x"2e190b",x"2b180b",x"2d190b",x"2d190b",x"2c180a",x"2c180a",x"2b160a",x"2a170a",x"2a170a",x"2e1a0b",x"321c0c",x"2f1a0b",x"311b0c",x"2d190b",x"28170a",x"2c190b",x"321c0d",x"321c0c",x"2d1a0b",x"2f1a0b",x"2b180a",x"2b170a",x"2f1a0b",x"2d1a0b",x"2b180b",x"2e1a0c",x"1d1108",x"1f1208",x"201309",x"201309",x"201308",x"201208",x"27160a",x"26160a",x"201208",x"241409",x"251509",x"28170a",x"28170a",x"2a180b",x"29170a",x"2f1b0c",x"2c190b",x"2c190b",x"2d190b",x"2b180b",x"2b180a",x"27160a",x"271509",x"261509",x"251509",x"29170a",x"2a180a",x"29170a",x"27160a",x"29170a",x"2b180a",x"291609",x"2a170a",x"2a180a",x"29170a",x"2c190b",x"2d190b",x"2d1a0b",x"2c190b",x"2d190b",x"2f1b0d",x"301c0d",x"2f1b0c",x"2c190b",x"2d190b",x"2d190b",x"2e1a0b",x"2f1b0c",x"2f1b0c",x"2e1b0c",x"2f1b0d",x"2d1a0c",x"2f1c0d",x"2f1b0c",x"2f1b0c",x"2d190b",x"2c190b",x"2b180a",x"2b180b",x"2b180b",x"2c190b",x"2b180b",x"2d190b",x"2b180b",x"2d190b",x"2a180b",x"28170a",x"29170a",x"28170a",x"26160a",x"26160a",x"2c190b",x"2c190b",x"29180b",x"27160a",x"2b190b",x"26160a",x"231409",x"26160a",x"251509",x"29170a",x"29170a",x"251409",x"281509",x"241409",x"28160a",x"2a180b",x"29170a",x"2a180b",x"2f1a0b",x"2d1a0b",x"311c0c",x"331d0d",x"1c1108",x"1c1108",x"1c1108",x"1b1008",x"1a1008",x"1d1208",x"221509",x"25150a",x"1f1309",x"24150a",x"231509",x"201309",x"2e1b0b",x"311c0b",x"1a1107",x"191007",x"191007",x"000000",x"000000",x"000000",x"515151",x"515151",x"313131",x"333333",x"505050",x"393939",x"383838",x"343434",x"373737",x"383838",x"323232",x"313131",x"2e2e2e",x"313131",x"2f3030",x"2f2f2f",x"333333",x"323232",x"323232",x"333333",x"3f3f3f",x"444444",x"494949",x"484848",x"484848",x"424242",x"3a3a3a",x"313131",x"323232",x"000000",x"333333",x"323232",x"323232",x"313131",x"333333",x"333333",x"333232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"323232",x"323232",x"2e2e2e",x"303030",x"2d2d2d",x"333333",x"343434",x"303030",x"323232",x"2e2e2e",x"333333",x"2e2e2e",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333232",x"313131",x"313131",x"303030",x"323232",x"313131",x"343434",x"353535",x"3b3b3b",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"2d2d2d",x"333333",x"313131",x"2e2e2e",x"343333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"452611",x"452611",x"4e2c14",x"4f2d15",x"4c2b14",x"452610",x"42230f",x"462610",x"3f220f",x"432410",x"4f3423",x"4b2a13",x"4a2912",x"452611",x"482913",x"4b2a13",x"4b2912",x"4b2f1d",x"4b2f1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"532f16",x"532f16",x"4f4238",x"493d34",x"4e3f34",x"4f4136",x"58493d",x"5b4a3d",x"5c4d41",x"594a3e",x"594c41",x"56493e",x"534439",x"56483d",x"56463a",x"59483b",x"57493e",x"55473c",x"53463c",x"56473a",x"57483c",x"57493d",x"58483d",x"5a493b",x"574539",x"564235",x"503e32",x"43392f",x"4b3e33",x"4b3e33",x"5e4534",x"483a2f",x"523f32",x"554437",x"5a4537",x"5d4a3d",x"654e3e",x"5c4b3f",x"644d3c",x"5d4c3e",x"5a4d41",x"594c42",x"574c41",x"5f4f42",x"58483c",x"604838",x"41352b",x"3d3127",x"3c2e25",x"362d26",x"3e2f25",x"403125",x"332921",x"312a22",x"332a21",x"403024",x"3c2f26",x"403228",x"48372b",x"3a3028",x"44352a",x"47382d",x"4f3d30",x"433931",x"484037",x"55483d",x"5b483a",x"56493e",x"524033",x"57483c",x"5d4a3d",x"524338",x"54453a",x"5a493c",x"54463b",x"574537",x"5c4b3e",x"5d4d41",x"5f4e43",x"5a4a3f",x"604d40",x"5a4b3f",x"5f4f42",x"6b5647",x"675344",x"5e4f42",x"615043",x"665447",x"5b4d41",x"5b4f43",x"4c3b2f",x"4c3b2f",x"000000",x"301e12",x"301e12",x"281b11",x"20160f",x"20160e",x"291a10",x"26180e",x"25170b",x"27180c",x"251509",x"281609",x"271509",x"241409",x"231409",x"28170a",x"2d190b",x"2d1a0b",x"2b190b",x"2b180b",x"2a170a",x"221409",x"241409",x"29170a",x"271509",x"291609",x"261509",x"2a180a",x"28160a",x"29170a",x"231409",x"221409",x"28160a",x"2c180a",x"2d190b",x"2c180a",x"2b180a",x"271609",x"231409",x"1e1208",x"1d1108",x"1b1008",x"1c1108",x"1c1108",x"221409",x"1e1208",x"1f1309",x"25160a",x"27170a",x"2a170a",x"27160a",x"2b190b",x"311c0d",x"2e1a0c",x"311c0d",x"301b0c",x"2f1a0c",x"301b0c",x"331c0d",x"341c0d",x"301b0c",x"341d0d",x"341e0d",x"311c0c",x"341d0e",x"331e0e",x"351f0e",x"37200f",x"351e0e",x"331e0e",x"331d0e",x"2e1a0c",x"311c0d",x"311c0c",x"331d0d",x"2f1b0c",x"321d0d",x"2f1b0c",x"321c0d",x"311b0c",x"2f1b0c",x"2d1a0b",x"311c0c",x"2f1a0b",x"2e1a0b",x"2b180a",x"2b180a",x"2b180a",x"2b170a",x"29170a",x"2c180b",x"2f1a0b",x"331d0d",x"301b0c",x"311c0d",x"2f1b0c",x"321d0d",x"28170a",x"301b0c",x"2c180b",x"28160a",x"2d1a0b",x"261609",x"221409",x"2b180b",x"2d1a0b",x"1c1108",x"1d1208",x"201309",x"211309",x"221409",x"241509",x"221409",x"221409",x"241409",x"261609",x"261509",x"27160a",x"28170a",x"27160a",x"2b180b",x"2c190b",x"29170a",x"271609",x"28160a",x"261509",x"261509",x"261509",x"261509",x"28160a",x"28160a",x"29170a",x"28170a",x"29170a",x"261509",x"271609",x"29170a",x"29170a",x"28170a",x"29170a",x"29170a",x"2c190b",x"2e1a0b",x"2c190b",x"2b180b",x"2e1a0c",x"311c0c",x"2f1b0c",x"2f1b0c",x"2d1a0c",x"2f1a0c",x"2c190b",x"2c180b",x"2e1a0b",x"2f1b0c",x"2f1a0c",x"2d1a0c",x"2f1b0c",x"2b190b",x"2b180b",x"2c190b",x"2a180b",x"2c190b",x"2f1a0b",x"2c190b",x"2e1a0c",x"2e1b0c",x"311c0d",x"2f1b0c",x"2f1b0c",x"2e1a0c",x"2e1a0c",x"2e1b0c",x"301b0d",x"29180b",x"27170a",x"2b190b",x"2f1b0c",x"29180b",x"29180a",x"2d1a0b",x"2a180b",x"29170a",x"241509",x"2e1a0b",x"2b180b",x"29170a",x"2a170a",x"261509",x"281609",x"251409",x"261509",x"261509",x"2a170a",x"2d190b",x"2c190b",x"311c0d",x"2e1b0c",x"2f1b0c",x"1d1208",x"1d1108",x"1c1108",x"1b1108",x"1c1108",x"1d1208",x"231409",x"28160a",x"241509",x"29170a",x"27160a",x"26160a",x"2b190a",x"2d190b",x"1a1107",x"191007",x"191007",x"000000",x"000000",x"000000",x"514f4e",x"514f4e",x"4e4d4d",x"545454",x"454545",x"4b4b4b",x"494949",x"515151",x"616161",x"595959",x"2c2d2d",x"333333",x"313131",x"2b2b2b",x"2f2f2f",x"303030",x"313131",x"3a3a3a",x"3d3d3d",x"373737",x"373737",x"353535",x"3b3b3b",x"3b3b3b",x"3e3f3f",x"383838",x"323232",x"313131",x"323232",x"333333",x"333333",x"333333",x"4e4e4e",x"353535",x"404040",x"3e3e3e",x"2e2e2e",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"333333",x"323232",x"3d3d3d",x"464646",x"414141",x"3e3e3e",x"353535",x"333333",x"414141",x"3d3d3d",x"333333",x"343434",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"414141",x"414141",x"535353",x"434343",x"494949",x"333333",x"3d3d3d",x"4f4f4f",x"323232",x"333333",x"333333",x"323130",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"2d2d2d",x"333333",x"313131",x"2e2e2e",x"343333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"452611",x"4e2c14",x"4f2d15",x"4c2b14",x"452610",x"42230f",x"462610",x"3f220f",x"432410",x"000000",x"4b2a13",x"4a2912",x"452611",x"482913",x"4b2a13",x"4b2912",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2b14",x"4b2b14",x"473c33",x"403329",x"4e3526",x"443125",x"4a3526",x"48362a",x"4f3b2d",x"4a3b30",x"4b3a2e",x"463429",x"473427",x"3f2e22",x"473528",x"593e2c",x"483528",x"4b3627",x"4e392b",x"4e392b",x"4e3b2c",x"51392b",x"4e382a",x"503625",x"583a26",x"4e3523",x"513321",x"4d3323",x"463224",x"4a3528",x"4f3727",x"3c2a1e",x"432e20",x"503727",x"573c2a",x"543a29",x"4d3626",x"5a3e2b",x"553a28",x"62422d",x"4d3829",x"4c382b",x"503b2c",x"553f2f",x"574031",x"453529",x"433125",x"3b2b20",x"35271d",x"37281e",x"2e231a",x"39281c",x"33241a",x"34241b",x"442c1d",x"533621",x"3b281c",x"3d281a",x"432c1d",x"482f1f",x"462f20",x"412d20",x"412d1f",x"3d2c21",x"3f3026",x"423226",x"4a3a2e",x"4c3a2e",x"543e2d",x"534033",x"513c2e",x"4c3c31",x"4e3c30",x"4f3a2b",x"533f31",x"5d4231",x"573f31",x"574336",x"544134",x"574235",x"503a2b",x"50392b",x"523a2b",x"563e2e",x"4f3d30",x"544236",x"56483c",x"685547",x"605044",x"5f4d3f",x"563c2c",x"563c2c",x"000000",x"2e1d12",x"2e1d12",x"271a11",x"20160e",x"22170f",x"24170d",x"26180e",x"23150b",x"20140a",x"211308",x"251509",x"241409",x"221409",x"28170a",x"281609",x"2d190b",x"28160a",x"2a180a",x"2b180a",x"271609",x"221409",x"241409",x"301b0b",x"2f1a0b",x"2f1a0b",x"2c190b",x"2b190b",x"26160a",x"29170a",x"221309",x"231408",x"29160a",x"2e190b",x"2f1a0b",x"2e1a0b",x"2a180b",x"29170a",x"241509",x"1a1008",x"190f07",x"1a1008",x"1a1008",x"1b1108",x"1e1208",x"1d1208",x"201309",x"24150a",x"25160a",x"2b180b",x"2e1a0b",x"2c190b",x"2a170a",x"28160a",x"2a170a",x"2d190b",x"2e1a0b",x"2e1a0b",x"2c190b",x"2f1a0b",x"301b0b",x"301b0c",x"2b180b",x"2b180b",x"2e1a0b",x"2e1a0b",x"311b0c",x"2f1a0c",x"2b180b",x"2f1a0c",x"2d190b",x"2e1a0c",x"2e1b0c",x"2f1b0c",x"2d190b",x"311c0c",x"2e1a0b",x"2c180b",x"2f1a0b",x"2d190b",x"2d190b",x"2f1a0b",x"2d180b",x"2c190b",x"2d190b",x"2e190b",x"2d190b",x"2d190b",x"311b0c",x"2c180a",x"2a180a",x"29170a",x"2d190b",x"2c190b",x"2e1a0b",x"2a180a",x"2a180b",x"2f1b0c",x"311c0c",x"28160a",x"29170a",x"2e1a0b",x"2e1a0b",x"28160a",x"2c180b",x"241509",x"1a1008",x"1d1108",x"1d1108",x"1f1208",x"1f1208",x"1f1208",x"211309",x"201308",x"231409",x"221309",x"29170a",x"29170a",x"29170a",x"28160a",x"28160a",x"2a170a",x"261509",x"281609",x"271509",x"29170a",x"2b180a",x"27160a",x"29170a",x"2b180b",x"2c190b",x"2c190b",x"29170a",x"251509",x"251509",x"261509",x"2b180a",x"2b180a",x"2a180a",x"2d190b",x"2e1a0b",x"2b180b",x"29170a",x"2c190b",x"301c0d",x"301c0d",x"321d0d",x"321d0d",x"301c0d",x"2d1a0b",x"2e1b0c",x"2c190b",x"2e1a0b",x"2d190b",x"29170a",x"271609",x"28160a",x"27160a",x"2a170a",x"2a180a",x"28170a",x"28170a",x"2a180a",x"2b180b",x"28160a",x"2a180a",x"2a180b",x"28170a",x"2c180b",x"27160a",x"28170a",x"29170a",x"2a170a",x"2a180b",x"25160a",x"29170b",x"25150a",x"29170a",x"29180b",x"27160a",x"27160a",x"26160a",x"27160a",x"221409",x"2a180a",x"28170a",x"29170a",x"2a180a",x"2d190b",x"2a170a",x"251509",x"28160a",x"28160a",x"251509",x"2d190b",x"2b180b",x"2a180a",x"2c190b",x"2b190b",x"1c1108",x"1d1108",x"1c1108",x"1b1108",x"1c1108",x"1c1108",x"1e1208",x"25150a",x"221409",x"231409",x"221309",x"241409",x"2a180a",x"2a180a",x"1d1208",x"1c1208",x"1c1208",x"000000",x"000000",x"000000",x"525252",x"4c4c4c",x"4b4b4b",x"454545",x"3a3a3a",x"444444",x"494949",x"525252",x"5a5a5a",x"5d5d5d",x"323232",x"333333",x"323232",x"313131",x"2f2f2f",x"2f2f2f",x"2f2f2f",x"383838",x"313131",x"2f2f2f",x"353535",x"2f2f2f",x"363636",x"353535",x"3c3c3c",x"3b3b3b",x"3d3d3d",x"323232",x"333333",x"333333",x"323232",x"2e2e2e",x"424242",x"505050",x"4d4d4d",x"4c4c4c",x"333333",x"323232",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"373737",x"373737",x"5e5e5e",x"606060",x"565656",x"575757",x"565656",x"515151",x"515151",x"484848",x"4d4d4d",x"505050",x"575757",x"565656",x"363636",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"565656",x"565656",x"333333",x"323232",x"434343",x"4c4c4c",x"484848",x"454545",x"545454",x"515151",x"333333",x"323232",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"565656",x"4a4a4a",x"323232",x"313131",x"2a2a2a",x"323232",x"323232",x"2e2e2e",x"000000",x"000000",x"000000",x"313131",x"313131",x"323232",x"333333",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"53321b",x"53321b",x"594537",x"4c392c",x"5c3e2a",x"463123",x"3f2e22",x"463020",x"473122",x"3c2b20",x"482f20",x"412c1e",x"492e1d",x"39251a",x"3c2517",x"472b19",x"3c2616",x"3f2818",x"3d281a",x"402c1e",x"4a3322",x"4c3221",x"432e1f",x"483020",x"4c3220",x"50331f",x"452d1d",x"482f1f",x"462f1f",x"472f1f",x"4a301e",x"3b271b",x"4a2f1c",x"452c1c",x"583821",x"4c321f",x"4b301d",x"472c1b",x"523420",x"523420",x"482e1c",x"442d1d",x"4d3221",x"483122",x"483324",x"443226",x"4a3324",x"3d2c20",x"392a1f",x"3d2b1e",x"3d291c",x"402819",x"352215",x"2f1e15",x"312115",x"3c2717",x"332015",x"3b2517",x"352216",x"412919",x"402919",x"3f281b",x"40291a",x"312016",x"362317",x"3c281a",x"402c1d",x"3d2c20",x"513522",x"513421",x"3c281c",x"422d1e",x"4b3220",x"422c1e",x"533622",x"503525",x"4e3526",x"513726",x"4e3524",x"4f3323",x"472e1f",x"4e311e",x"4d311f",x"472e1e",x"4a301f",x"4e3423",x"4c3629",x"594436",x"5a473a",x"655548",x"523b2d",x"523b2d",x"000000",x"311f13",x"311f13",x"2b1c11",x"241a12",x"23180e",x"24180d",x"29190f",x"21160b",x"20140a",x"1f1208",x"211409",x"201309",x"2a180b",x"251509",x"27160a",x"27160a",x"241509",x"201309",x"201309",x"201309",x"25150a",x"291709",x"2c1a0a",x"2c1a0a",x"2b190b",x"241609",x"231509",x"1f1208",x"1f1208",x"211308",x"261609",x"2e1b0a",x"2c190a",x"2b190a",x"2e190a",x"251508",x"1b1008",x"180f07",x"170f07",x"160e07",x"170f07",x"170f07",x"180f07",x"191008",x"1b1108",x"201309",x"28170a",x"221409",x"28160a",x"271509",x"261509",x"2a160a",x"2a170a",x"2c180a",x"2c180a",x"2a170a",x"2f1a0b",x"301b0c",x"301b0c",x"351d0d",x"331d0d",x"311c0d",x"321c0d",x"311c0d",x"2d1a0b",x"301b0c",x"311c0c",x"2f1a0b",x"2d190b",x"2e1a0b",x"2e190b",x"2a180a",x"2b180b",x"2c190b",x"2d190b",x"2c180a",x"2b180a",x"2d190b",x"2c190b",x"2c190a",x"2c180a",x"2d1a0a",x"2c190a",x"2d190b",x"301b0c",x"2e1a0b",x"2d190b",x"2c190b",x"2d190b",x"2a180a",x"2d190b",x"2e1a0b",x"2b180b",x"28160a",x"2f1b0c",x"331d0c",x"301b0c",x"2f1a0b",x"2e190b",x"321d0d",x"351e0e",x"2f1b0c",x"311c0c",x"26160a",x"26160a",x"1c1108",x"1e1208",x"211409",x"26170a",x"26170a",x"25160a",x"231409",x"28170a",x"2a180b",x"2c190b",x"29170b",x"26160a",x"2a190b",x"2a180b",x"2b180b",x"2a170a",x"2a180b",x"2b190b",x"2e1a0b",x"2d190b",x"28160a",x"29170a",x"2c190b",x"2a180b",x"2a180a",x"2a170a",x"261609",x"261509",x"251509",x"251509",x"231309",x"251409",x"261409",x"241308",x"241308",x"251409",x"271609",x"2b180a",x"2b180b",x"2d190b",x"2e1a0c",x"2f1b0c",x"2d1a0b",x"2d190b",x"2e1a0c",x"2a180b",x"261509",x"261509",x"241409",x"241409",x"251409",x"251409",x"251509",x"271609",x"28160a",x"27160a",x"2c190b",x"2c190b",x"2d190b",x"2c190b",x"2d1a0b",x"2e1a0c",x"2d190b",x"2b180b",x"2a180b",x"27160a",x"2b180b",x"29170a",x"2a180b",x"27160a",x"28160a",x"28170a",x"28160a",x"251509",x"251509",x"261509",x"281709",x"241509",x"2d190b",x"2c190a",x"2a180a",x"2c180b",x"2d190b",x"29170a",x"2b180a",x"2a170a",x"29170a",x"261509",x"2f1b0c",x"2b180b",x"2d190b",x"2c180b",x"2d1a0b",x"1d1108",x"1c1108",x"1b1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1a1008",x"1e1208",x"160e07",x"1b1108",x"201308",x"2c1a0a",x"301d0b",x"1f1309",x"201409",x"201409",x"000000",x"000000",x"000000",x"4a4a4a",x"414040",x"3f3f3f",x"434343",x"343434",x"3c3c3c",x"434343",x"4f4f4f",x"5e5e5e",x"626262",x"383838",x"313131",x"323232",x"323232",x"333333",x"362b26",x"323232",x"373737",x"363636",x"323232",x"323232",x"484848",x"2b2b2b",x"393939",x"363636",x"393939",x"3f3f3f",x"434343",x"454545",x"4a4a4a",x"343434",x"393939",x"404040",x"444444",x"424242",x"404040",x"4f4f4f",x"3a3a3a",x"343434",x"323232",x"323232",x"323232",x"313131",x"000000",x"000000",x"444444",x"3e3d3d",x"403e3d",x"3d3c3b",x"313131",x"4e4e4e",x"494949",x"525252",x"534a43",x"4b4b4b",x"585858",x"535353",x"444444",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"333333",x"313131",x"323232",x"323232",x"545454",x"424242",x"4c4c4c",x"505050",x"484848",x"535353",x"646464",x"646464",x"545454",x"545454",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"323232",x"323232",x"333333",x"515151",x"323232",x"4e4e4e",x"404040",x"353535",x"2e2e2e",x"2e2e2e",x"000000",x"000000",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"313131",x"323232",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2c190b",x"2c190b",x"4b2a13",x"482711",x"472711",x"462813",x"512f16",x"4f2d15",x"492a14",x"462913",x"4d2c15",x"4e2c14",x"4d2b14",x"4f2c15",x"4f2c14",x"4d2b14",x"523016",x"502e15",x"4c2a13",x"4f2d15",x"472711",x"502d15",x"4a2a13",x"513117",x"522f17",x"502e16",x"502e16",x"4d2d15",x"533117",x"533118",x"543218",x"523117",x"553319",x"533117",x"553218",x"583419",x"533117",x"4c2c15",x"4d2b14",x"573219",x"4c2b14",x"4e2c14",x"4e2b12",x"4a2912",x"472711",x"482812",x"4e2b14",x"4c2b14",x"4f2c15",x"4e2c15",x"4c2b14",x"4e2c15",x"4e2c14",x"502d15",x"522f16",x"482711",x"512f16",x"4e2d14",x"502e15",x"512e16",x"502e16",x"512e16",x"4f2d15",x"4d2c14",x"4f2d14",x"4d2b13",x"4e2d14",x"512e15",x"502d15",x"4b2a13",x"655041",x"56483d",x"493e34",x"533f32",x"403329",x"3b3027",x"332a23",x"3b2d23",x"3f2d21",x"3f2c1f",x"412b1d",x"462d1c",x"302217",x"462b19",x"291d15",x"362317",x"3a2518",x"412d1f",x"402e21",x"513828",x"49372b",x"4c392b",x"523b2b",x"483528",x"4c3729",x"4a372a",x"3e3229",x"4b3a2e",x"423226",x"352b23",x"382a21",x"402c1f",x"4e3524",x"453021",x"523521",x"482f1e",x"4a2f1e",x"4b3120",x"412c1e",x"412c1e",x"412f21",x"473325",x"443428",x"5a3d2b",x"392f27",x"3e3127",x"352d26",x"382d24",x"35281d",x"3d291c",x"382519",x"302016",x"2f2017",x"302115",x"352317",x"342316",x"2f2016",x"3c2719",x"322318",x"3f291b",x"2d2117",x"231b15",x"2b1e14",x"291d14",x"362519",x"2b2118",x"3a271a",x"352418",x"2b1e14",x"2d2016",x"302218",x"472d1a",x"4d3221",x"493224",x"442f23",x"473023",x"3a2a1f",x"3d2a1d",x"261e17",x"3c281a",x"412a1b",x"412a1b",x"34241a",x"3b291c",x"35281f",x"4b3a2e",x"5e493a",x"645243",x"4e3a2c",x"4e3a2c",x"000000",x"342114",x"342114",x"2d1d12",x"251a11",x"20170f",x"23170e",x"20160d",x"1f130b",x"1d1108",x"1f1309",x"24150a",x"241509",x"201309",x"201309",x"201309",x"211308",x"1f1208",x"1f1208",x"1c1108",x"1f1208",x"1f1208",x"251609",x"2b1a0a",x"2b190a",x"2d1b0b",x"231509",x"221408",x"1d1108",x"1d1108",x"211408",x"2a1909",x"2c1b0a",x"2c1b0a",x"29190a",x"29180a",x"201409",x"190f07",x"160e07",x"181007",x"180f07",x"180f07",x"150e07",x"160e07",x"170f07",x"191008",x"1a1008",x"1a1008",x"1b1008",x"1d1108",x"1f1309",x"201309",x"201309",x"211409",x"211409",x"221409",x"221409",x"221409",x"221409",x"221409",x"241509",x"25150a",x"25160a",x"26160a",x"27170a",x"26160a",x"24150a",x"231509",x"221409",x"211309",x"201309",x"1f1208",x"1e1208",x"1e1208",x"1f1208",x"201309",x"201309",x"201208",x"211309",x"201309",x"221408",x"2e1a0b",x"2e1a0b",x"2d190b",x"2b180a",x"2c180a",x"2a170a",x"28160a",x"2a180a",x"2c190b",x"2f1a0b",x"2b180b",x"2c190b",x"2b180b",x"2f1a0b",x"2d190b",x"341d0d",x"351d0d",x"321c0c",x"331d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"180f08",x"1b1108",x"1c1108",x"1e1308",x"24150a",x"211408",x"1f1208",x"1f1208",x"221409",x"221409",x"231509",x"221409",x"221409",x"231409",x"1f1208",x"221309",x"201308",x"211309",x"231409",x"201208",x"221409",x"221409",x"211309",x"1f1208",x"1f1208",x"1e1108",x"1e1208",x"201309",x"201309",x"211409",x"221409",x"221409",x"211309",x"221409",x"231409",x"231409",x"231409",x"241509",x"201208",x"201208",x"1f1108",x"211308",x"221409",x"211309",x"201208",x"1f1208",x"1f1208",x"221409",x"221409",x"221409",x"221409",x"231509",x"23150a",x"231509",x"231409",x"211409",x"201309",x"1f1309",x"1f1309",x"1e1208",x"1e1208",x"1e1208",x"1d1208",x"1d1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"1b1008",x"1b1108",x"1b1108",x"1d1108",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"201209",x"201308",x"271809",x"251609",x"231609",x"231509",x"1c1107",x"1c1107",x"170f07",x"1a1007",x"160e07",x"170f07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1b1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1b1108",x"191008",x"180f08",x"170f07",x"160e07",x"150e07",x"150e07",x"1f1408",x"2d1d0a",x"2d1c0a",x"311d0b",x"321e0b",x"321e0b",x"000000",x"000000",x"000000",x"3d3d3d",x"383838",x"3b3b3b",x"3f3f3f",x"303030",x"363636",x"3b3b3b",x"434343",x"595959",x"5d5d5d",x"4e4e4e",x"323232",x"323232",x"313131",x"333333",x"313131",x"303030",x"323232",x"343434",x"3d3d3d",x"323232",x"454545",x"3f3f3f",x"3b3b3b",x"373737",x"3a3a3a",x"3d3d3d",x"3d3d3d",x"3c3c3c",x"424242",x"3a3a3a",x"353535",x"3d3d3d",x"3c3c3c",x"3b3b3b",x"363636",x"424242",x"444444",x"4b4b4b",x"4a4a4a",x"343434",x"303030",x"323232",x"323232",x"323232",x"333333",x"333333",x"2e2e2e",x"393836",x"323232",x"303030",x"464646",x"404040",x"493d38",x"4c4c4c",x"474747",x"323232",x"323130",x"343434",x"313131",x"333333",x"323131",x"333333",x"323232",x"323232",x"303030",x"333333",x"323232",x"323232",x"323232",x"323232",x"313131",x"313131",x"333333",x"333333",x"323232",x"313131",x"313131",x"353535",x"575757",x"4d4d4d",x"4c4c4c",x"4a4a4a",x"454545",x"404040",x"454340",x"494643",x"514f4c",x"585858",x"323232",x"323232",x"2d2d2d",x"2f2f2f",x"313131",x"323232",x"313131",x"313131",x"303030",x"323232",x"3d3d3d",x"4b4b4b",x"585858",x"3b3b3b",x"474747",x"525252",x"282828",x"282828",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"343434",x"343434",x"323232",x"333333",x"313131",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2c190b",x"2c190b",x"4b2a13",x"482711",x"472711",x"462813",x"512f16",x"4f2d15",x"492a14",x"462913",x"4d2c15",x"4e2c14",x"4d2b14",x"4f2c15",x"4f2c14",x"4d2b14",x"523016",x"502e15",x"4c2a13",x"4f2d15",x"472711",x"502d15",x"4a2a13",x"513117",x"522f17",x"502e16",x"502e16",x"4d2d15",x"533117",x"533118",x"543218",x"523117",x"553319",x"533117",x"553218",x"583419",x"533117",x"4c2c15",x"4d2b14",x"573219",x"4c2b14",x"4e2c14",x"4e2b12",x"4a2912",x"472711",x"482812",x"4e2b14",x"4c2b14",x"4f2c15",x"4e2c15",x"4c2b14",x"4e2c15",x"4e2c14",x"502d15",x"522f16",x"482711",x"512f16",x"4e2d14",x"502e15",x"512e16",x"502e16",x"512e16",x"4f2d15",x"4d2c14",x"4f2d14",x"4d2b13",x"4e2d14",x"512e15",x"502d15",x"4e2c14",x"4b2913",x"502e15",x"3e220e",x"3e210d",x"4a2911",x"43240f",x"46260f",x"4e2b12",x"492810",x"452610",x"482913",x"482812",x"4a2a13",x"4a2b14",x"4b2a14",x"482913",x"4f2e15",x"4a2a13",x"432c1d",x"412d20",x"442f22",x"493324",x"4a3324",x"4b3424",x"4d3423",x"4e3524",x"4a3425",x"4d3424",x"4a3323",x"482f1f",x"4f3320",x"4e3220",x"4d311e",x"3f291b",x"3f291a",x"4b2e1b",x"412818",x"3d2718",x"392517",x"3b2719",x"3d291b",x"442d1d",x"4b3120",x"452e1d",x"412f22",x"432e1f",x"432d1e",x"422c1c",x"3e2819",x"3f2717",x"3e2616",x"362214",x"321f12",x"2b1b11",x"382214",x"322013",x"321f12",x"3d2616",x"352013",x"3a2415",x"412717",x"422817",x"412815",x"362112",x"372214",x"3c2617",x"432917",x"342012",x"281a10",x"311f12",x"372213",x"3a2415",x"3d2718",x"3c271a",x"3c281a",x"492e1c",x"462b1a",x"3d2617",x"3f2717",x"452b19",x"432816",x"3b2414",x"3a2214",x"3a2415",x"3f291a",x"4c3b2f",x"5a483b",x"604f42",x"442f21",x"442f21",x"000000",x"311f13",x"311f13",x"2c1d11",x"22180f",x"21170f",x"23160d",x"21140a",x"1f130b",x"241509",x"2b180b",x"29180a",x"1e1208",x"231409",x"221409",x"1f1208",x"201308",x"1f1208",x"29170a",x"221409",x"1b1008",x"241509",x"28170a",x"221409",x"251609",x"2b180b",x"29170a",x"2c190b",x"241509",x"1c1108",x"1e1208",x"29180a",x"301c0c",x"241609",x"1f1308",x"221409",x"261609",x"241509",x"1d1108",x"1d1208",x"1a1008",x"160e07",x"160e07",x"160f07",x"1c1108",x"1a1008",x"1b1108",x"1b1008",x"1e1208",x"201309",x"24150a",x"23150a",x"231409",x"221409",x"2a190b",x"27170a",x"2a180b",x"28170b",x"28180b",x"2c1a0c",x"2c190b",x"27160a",x"29170a",x"29170a",x"231409",x"28170a",x"27160a",x"29170a",x"231509",x"241509",x"231409",x"241509",x"25150a",x"231509",x"251509",x"241509",x"221409",x"201308",x"231409",x"251509",x"211408",x"2c190a",x"301a0b",x"2d180a",x"2f1a0b",x"321c0c",x"2d190b",x"2e190b",x"301b0c",x"321b0c",x"321c0c",x"361f0e",x"38200e",x"321d0d",x"3c2311",x"3c2312",x"371f0e",x"371f0d",x"381f0e",x"3b210f",x"2f1b0c",x"23150a",x"150e07",x"150e07",x"160e07",x"170f07",x"180f08",x"1a1008",x"1a1008",x"1b1008",x"1d1108",x"1e1208",x"1f1209",x"201309",x"211409",x"211409",x"221409",x"221409",x"211308",x"1e1208",x"221409",x"221409",x"201308",x"221409",x"211309",x"1e1208",x"1f1208",x"201309",x"1f1208",x"1f1208",x"1f1208",x"1e1208",x"1e1208",x"201309",x"221409",x"221409",x"231409",x"231409",x"231409",x"241509",x"241509",x"25150a",x"25160a",x"25160a",x"241509",x"231409",x"241509",x"241509",x"241509",x"221409",x"211309",x"24150a",x"23150a",x"23150a",x"211309",x"1f1208",x"221409",x"221409",x"221409",x"221409",x"221409",x"211409",x"201309",x"1e1208",x"1d1208",x"1c1108",x"1b1008",x"1b1108",x"1b1108",x"1b1108",x"1b1108",x"1b1008",x"1a1008",x"1a1008",x"1b1108",x"1c1108",x"1d1108",x"1d1208",x"1e1208",x"1f1208",x"1f1208",x"1f1208",x"231509",x"2a1a0a",x"2a1a0a",x"271709",x"291a0a",x"221509",x"271808",x"291a09",x"241608",x"1a1007",x"191007",x"160e07",x"170f07",x"191008",x"1a1108",x"1c1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1b1108",x"1a1008",x"191008",x"180f07",x"160f07",x"150e07",x"160f07",x"1a1107",x"211508",x"311f0a",x"2d1c0a",x"3c230e",x"3c230d",x"3c230d",x"000000",x"000000",x"000000",x"363636",x"4c4c4c",x"4b4b4b",x"313131",x"333333",x"333333",x"333333",x"323232",x"302d2a",x"313131",x"323232",x"323232",x"343433",x"313131",x"333333",x"323232",x"323232",x"333333",x"353535",x"363636",x"363636",x"313131",x"323232",x"343434",x"323232",x"383838",x"3c3c3c",x"3a3a3a",x"3c3c3c",x"3c3c3c",x"3d3d3d",x"3d3937",x"3f3f3f",x"363636",x"363636",x"3a3a3a",x"363636",x"3f3f3f",x"3c3c3c",x"434343",x"4a4a4a",x"515151",x"323232",x"323232",x"303030",x"323232",x"333333",x"323232",x"2c2c2c",x"4b4b4b",x"3f3f3f",x"393939",x"373737",x"3b3b3b",x"333333",x"323232",x"323232",x"323232",x"343434",x"313131",x"333333",x"323131",x"333333",x"323232",x"323232",x"303030",x"323232",x"434343",x"474747",x"2e2e2e",x"313131",x"313131",x"313131",x"333333",x"333333",x"323232",x"404040",x"4b4b4b",x"474747",x"434343",x"3c3c3c",x"383838",x"363636",x"2f2f2f",x"323232",x"313131",x"333333",x"323232",x"333333",x"323232",x"323232",x"2d2d2d",x"2f2f2f",x"313131",x"323232",x"323232",x"303030",x"494949",x"4d4d4d",x"4a4a4a",x"474747",x"414141",x"474747",x"484848",x"414141",x"323232",x"323232",x"323232",x"323232",x"323232",x"383838",x"383838",x"3c3c3c",x"383838",x"323232",x"36312d",x"333333",x"323232",x"323232",x"333333",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"5e4c3f",x"5e4c3f",x"3b200e",x"26160a",x"3b200e",x"3a200e",x"381f0d",x"361e0d",x"2f1a0c",x"38200e",x"150e07",x"2e1b0c",x"3a210f",x"3c210f",x"432511",x"3e220f",x"3d2310",x"3d220f",x"3e230f",x"3f2310",x"391f0e",x"381f0e",x"3c2210",x"422611",x"412410",x"3a200e",x"3a200e",x"3b200e",x"3c210e",x"3c210e",x"3b200e",x"412410",x"412410",x"412410",x"3b200e",x"381e0d",x"381e0c",x"351c0c",x"3c210e",x"412511",x"412511",x"422511",x"3f220f",x"3f230f",x"3f220f",x"391e0c",x"371d0d",x"3f230f",x"3d2310",x"402410",x"432611",x"402410",x"3d220f",x"3d210f",x"402310",x"422611",x"412511",x"432611",x"432611",x"3f230f",x"3b200e",x"3b200e",x"3a1f0d",x"3b200e",x"3a1f0d",x"391f0d",x"381e0c",x"371d0c",x"361c0c",x"3b200e",x"3d220f",x"3d210f",x"3e220f",x"381f0c",x"361e0c",x"40230f",x"331c0b",x"301a0a",x"351d0c",x"3a1f0d",x"381f0c",x"341c0c",x"341e0d",x"2d190b",x"301b0c",x"150e07",x"2a170a",x"150e07",x"150e07",x"412d20",x"442f22",x"493324",x"4a3324",x"4b3424",x"4d3423",x"4e3524",x"4a3425",x"4d3424",x"4a3323",x"482f1f",x"4f3320",x"4e3220",x"4d311e",x"3f291b",x"3f291a",x"4b2e1b",x"412818",x"3d2718",x"392517",x"3b2719",x"3d291b",x"442d1d",x"4b3120",x"452e1d",x"412f22",x"432e1f",x"432d1e",x"422c1c",x"3e2819",x"3f2717",x"3e2616",x"362214",x"321f12",x"2b1b11",x"382214",x"322013",x"321f12",x"3d2616",x"352013",x"3a2415",x"412717",x"422817",x"412815",x"362112",x"372214",x"3c2617",x"432917",x"342012",x"281a10",x"311f12",x"372213",x"3a2415",x"3d2718",x"3c271a",x"3c281a",x"492e1c",x"462b1a",x"3d2617",x"3f2717",x"452b19",x"432816",x"3b2414",x"3a2214",x"3a2415",x"3f291a",x"4c3b2f",x"5a483b",x"604f42",x"442f21",x"000000",x"000000",x"1f1710",x"1f1710",x"211811",x"22170f",x"24180f",x"21160d",x"1e130a",x"1a110a",x"160e07",x"2c190b",x"201309",x"1f1209",x"1f1209",x"4a2c16",x"211409",x"201309",x"201309",x"201309",x"311b0b",x"361e0c",x"201208",x"221409",x"241509",x"26160a",x"29170a",x"29170a",x"27160a",x"211409",x"211309",x"26160a",x"251509",x"251509",x"25150a",x"211309",x"1d1108",x"1f1208",x"201308",x"221409",x"201208",x"211308",x"201308",x"1c1108",x"1d1108",x"201308",x"1f1208",x"201308",x"241509",x"201208",x"1d1108",x"1f1208",x"25160a",x"26160a",x"27170a",x"26160a",x"25160a",x"211409",x"221409",x"25150a",x"26160a",x"28170a",x"27160a",x"26160a",x"241509",x"241509",x"261609",x"27160a",x"24150a",x"26160a",x"231509",x"201309",x"201309",x"211309",x"231409",x"231409",x"241509",x"251509",x"241409",x"221309",x"251509",x"28170a",x"241509",x"261609",x"241409",x"211309",x"201209",x"201309",x"231409",x"221409",x"201308",x"1f1208",x"1b1108",x"191007",x"1c120a",x"21150b",x"20140b",x"201409",x"201209",x"1f1208",x"1d1208",x"1c1108",x"170f07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1a1008",x"1c1108",x"1d1108",x"201309",x"201309",x"201208",x"201309",x"211309",x"211309",x"211309",x"221409",x"221408",x"221309",x"221409",x"231409",x"251509",x"251509",x"251509",x"251609",x"251509",x"241409",x"24150a",x"24150a",x"231409",x"221409",x"231409",x"221409",x"221309",x"241509",x"251609",x"241509",x"251609",x"241409",x"231509",x"231409",x"231409",x"241409",x"231409",x"211308",x"211308",x"211308",x"211308",x"221409",x"241509",x"241509",x"261609",x"26160a",x"25150a",x"241509",x"241509",x"26150a",x"27170a",x"251509",x"25150a",x"231509",x"211309",x"201309",x"211309",x"201309",x"221409",x"211409",x"1f1209",x"1c1108",x"1d1209",x"1f1209",x"1f1209",x"1f1209",x"1e1209",x"1d1108",x"1c1008",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"211408",x"231509",x"281909",x"2b1b0a",x"291a0a",x"301e0a",x"2b1b09",x"2e1d0a",x"221508",x"1e1308",x"1a1107",x"191007",x"160e07",x"170f07",x"180f07",x"190f08",x"1a1008",x"1c1008",x"201309",x"201209",x"211409",x"1e1108",x"1b1008",x"170f07",x"191008",x"1f1208",x"211309",x"221409",x"1f1308",x"271809",x"2d1c0a",x"2d1c0a",x"2e1a0b",x"432510",x"000000",x"000000",x"000000",x"000000",x"505050",x"505050",x"494949",x"333333",x"343434",x"323232",x"323131",x"323232",x"302d2b",x"313131",x"323232",x"323232",x"333333",x"2a2a2a",x"313131",x"333333",x"333333",x"313131",x"323232",x"393939",x"3a3a3a",x"3c3c3c",x"383838",x"393939",x"323232",x"393939",x"3b3b3b",x"3a3a3a",x"3a3a3a",x"3a3a3a",x"3a3a3a",x"3a3a3a",x"3a3a3a",x"3b3b3b",x"3c3c3c",x"3a3a3a",x"353535",x"404040",x"3d3d3d",x"414141",x"434242",x"444444",x"3d3d3d",x"4c4c4c",x"4f4f4f",x"505050",x"424242",x"4d4d4d",x"3c3c3c",x"3e3e3e",x"3f3f3f",x"3c3c3c",x"3e3e3e",x"3b3b3b",x"3d3d3d",x"46423f",x"4d4d4d",x"555555",x"4c4c4c",x"4d4d4d",x"505050",x"515151",x"505050",x"4e4e4e",x"4c4c4c",x"4a4a4a",x"484848",x"444444",x"444444",x"3c3c3c",x"474747",x"515151",x"565656",x"525252",x"494949",x"4b4b4b",x"3c3c3c",x"343434",x"282828",x"343434",x"393939",x"3c3c3c",x"3d3d3d",x"3a3a3a",x"444444",x"434343",x"464646",x"4a4a4a",x"515151",x"4f4f4f",x"535353",x"525252",x"505050",x"4f4f4f",x"505050",x"494949",x"484848",x"414141",x"3e3e3e",x"383838",x"343434",x"323232",x"323232",x"323232",x"373737",x"404040",x"4a4a4a",x"4a4a4a",x"434343",x"3b3b3b",x"343434",x"393939",x"383838",x"3f3f3f",x"343434",x"323232",x"323232",x"313131",x"323232",x"3d3d3d",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d3c30",x"4d3c30",x"351d0d",x"1b1008",x"371e0d",x"371e0d",x"28160a",x"2c180b",x"2f1a0b",x"301a0b",x"150e07",x"241308",x"2b1609",x"2c1609",x"211006",x"221006",x"221006",x"221006",x"251207",x"321a0b",x"351c0c",x"311b0b",x"311b0b",x"341c0c",x"361e0d",x"371e0d",x"381f0d",x"371f0d",x"3a210e",x"3f2310",x"402410",x"402410",x"3f240f",x"3c210e",x"371e0d",x"381e0d",x"391f0d",x"361d0c",x"361d0c",x"391f0d",x"422510",x"3e230f",x"432711",x"422611",x"482a14",x"422511",x"3e220f",x"3d220f",x"432611",x"432712",x"412611",x"422611",x"432611",x"432612",x"442712",x"402511",x"432611",x"452812",x"472914",x"432612",x"462813",x"472913",x"432612",x"422611",x"412410",x"402410",x"3c220f",x"3d210f",x"3e220f",x"3c210e",x"3a1f0d",x"3a200e",x"3c210e",x"3d220f",x"381f0c",x"351c0b",x"3a200d",x"3b200d",x"341d0c",x"341c0b",x"321b0b",x"29170a",x"29170a",x"2c180a",x"2a1609",x"150e07",x"261509",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211811",x"211811",x"241911",x"24180f",x"25180f",x"25180d",x"21150b",x"23150a",x"160f07",x"341e0d",x"221409",x"1f1209",x"51301a",x"452915",x"191008",x"412410",x"201309",x"201309",x"311b0b",x"361e0c",x"201208",x"221409",x"241509",x"26160a",x"29170a",x"29170a",x"27160a",x"211409",x"211309",x"26160a",x"251509",x"251509",x"25150a",x"211309",x"1d1108",x"1f1208",x"201308",x"221409",x"201208",x"211308",x"201308",x"1c1108",x"1d1108",x"201308",x"1f1208",x"201308",x"241509",x"201208",x"1d1108",x"1f1208",x"25160a",x"26160a",x"27170a",x"26160a",x"25160a",x"211409",x"221409",x"25150a",x"26160a",x"28170a",x"27160a",x"26160a",x"241509",x"241509",x"261609",x"27160a",x"24150a",x"26160a",x"231509",x"201309",x"201309",x"211309",x"231409",x"231409",x"241509",x"251509",x"241409",x"221309",x"251509",x"28170a",x"241509",x"261609",x"241409",x"211309",x"201209",x"201309",x"231409",x"221409",x"201308",x"1f1208",x"1b1108",x"191007",x"1c120a",x"21150b",x"20140b",x"201409",x"201209",x"1f1208",x"1d1208",x"1c1108",x"170f07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1a1008",x"1c1108",x"1d1108",x"201309",x"201309",x"201208",x"201309",x"211309",x"211309",x"211309",x"221409",x"221408",x"221309",x"221409",x"231409",x"251509",x"251509",x"251509",x"251609",x"251509",x"241409",x"24150a",x"24150a",x"231409",x"221409",x"231409",x"221409",x"221309",x"241509",x"251609",x"241509",x"251609",x"241409",x"231509",x"231409",x"231409",x"241409",x"231409",x"211308",x"211308",x"211308",x"211308",x"221409",x"241509",x"241509",x"261609",x"26160a",x"25150a",x"241509",x"241509",x"26150a",x"27170a",x"251509",x"25150a",x"231509",x"211309",x"201309",x"211309",x"201309",x"221409",x"211409",x"1f1209",x"1c1108",x"1d1209",x"1f1209",x"1f1209",x"1f1209",x"1e1209",x"1d1108",x"1c1008",x"1e1208",x"1e1208",x"1f1208",x"1f1208",x"211408",x"231509",x"281909",x"2b1b0a",x"291a0a",x"301e0a",x"2b1b09",x"2e1d0a",x"221508",x"1e1308",x"1a1107",x"191007",x"160e07",x"170f07",x"180f07",x"190f08",x"1a1008",x"1c1008",x"201309",x"201209",x"211409",x"1e1108",x"1b1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"433a32",x"463d34",x"4a4137",x"4a4137",x"2e1a0b",x"432510",x"000000",x"000000",x"000000",x"000000",x"000000",x"505050",x"494949",x"333333",x"343434",x"333333",x"323131",x"323232",x"302d2b",x"000000",x"000000",x"323232",x"323232",x"323232",x"333333",x"313131",x"524c49",x"323232",x"353535",x"343434",x"383838",x"333333",x"333333",x"353535",x"323232",x"393939",x"3a3a3a",x"383838",x"3b3b3b",x"373737",x"3d3d3d",x"3a3a3a",x"393939",x"373737",x"3a3a3a",x"3c3c3c",x"3b3b3b",x"3a3a3a",x"3e3e3e",x"414141",x"3f3f3f",x"404040",x"414141",x"414141",x"404040",x"444444",x"3d3d3d",x"3e3e3e",x"434343",x"3e3e3e",x"3d3d3d",x"3f3f3f",x"3c3c3c",x"353535",x"3f3f3f",x"3d3d3d",x"444444",x"434343",x"434343",x"454545",x"434343",x"464646",x"434343",x"474747",x"484848",x"494949",x"434343",x"414141",x"3a3a3a",x"434343",x"434343",x"414141",x"454545",x"424242",x"3a3a3a",x"3f3f3f",x"424242",x"2e2e2e",x"515151",x"373737",x"4b4b4b",x"3e3e3e",x"383838",x"3d3d3d",x"414141",x"424242",x"414141",x"464646",x"444444",x"484848",x"454545",x"464646",x"424242",x"414141",x"434343",x"454545",x"3f3f3f",x"3e3e3e",x"3b3b3b",x"3e3e3e",x"383838",x"4b4b4b",x"4c4c4c",x"3b3b3b",x"3f3f3f",x"414141",x"414141",x"454545",x"3f3f3f",x"3c3c3c",x"3e3e3e",x"444444",x"4b4b4b",x"454545",x"3b3b3b",x"323232",x"474747",x"444444",x"363636",x"3b3b3b",x"464646",x"3c3c3c",x"3c3c3c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3f2f24",x"3f2f24",x"39200e",x"2c190b",x"381f0e",x"341c0c",x"180f08",x"150e07",x"27160a",x"321c0c",x"150e07",x"311c0c",x"371f0e",x"3d220f",x"3e220f",x"402410",x"3c210e",x"371d0c",x"3b200e",x"3e230f",x"402410",x"3c210f",x"3f230f",x"3f2410",x"402410",x"3c210f",x"391f0d",x"371e0d",x"3f2310",x"402410",x"432611",x"412511",x"402310",x"3c210e",x"3e220f",x"3f240f",x"3e220f",x"422611",x"3f2310",x"412511",x"3f2310",x"3f2410",x"412411",x"3f2310",x"402510",x"422510",x"402411",x"3f2410",x"3b200e",x"3a200e",x"412511",x"432611",x"452812",x"402410",x"3c210e",x"371d0c",x"3c210f",x"3f230f",x"3a1f0d",x"3a1f0d",x"402310",x"3f2310",x"422611",x"412410",x"3f230f",x"391f0d",x"3f220f",x"40230f",x"3c210f",x"3f230f",x"3b200e",x"3b200e",x"3d210f",x"391f0d",x"402510",x"3e230e",x"3a200d",x"3c210e",x"351d0c",x"3c210e",x"361e0c",x"241509",x"150e07",x"211409",x"321c0c",x"150e07",x"321c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221911",x"221911",x"251911",x"26190f",x"281a10",x"29190e",x"26190e",x"21140b",x"170f07",x"38200e",x"2a180a",x"51321b",x"2f1d10",x"412614",x"422613",x"27170b",x"3b2212",x"311c0c",x"3b2211",x"402411",x"412411",x"422613",x"432511",x"442610",x"462711",x"422510",x"442611",x"482812",x"452712",x"472912",x"4a2a13",x"452711",x"432511",x"3f230f",x"422410",x"412410",x"412410",x"432511",x"482913",x"4c2c14",x"4c2c15",x"4e2e15",x"472913",x"482913",x"492914",x"4a2a13",x"4d2c15",x"4d2d15",x"4d2d15",x"4a2a14",x"452712",x"452611",x"462712",x"432511",x"4a2a14",x"472812",x"502f17",x"523118",x"4c2d15",x"492913",x"452711",x"4c2c14",x"4a2a14",x"482914",x"4b2b14",x"482812",x"482812",x"4a2a14",x"462712",x"452712",x"482812",x"442711",x"462812",x"4f2e16",x"512f17",x"502f16",x"4d2c14",x"4c2b15",x"4b2b14",x"4e2d15",x"4d2c15",x"472712",x"452711",x"472812",x"492812",x"492812",x"472711",x"492812",x"4b2b14",x"4c2b14",x"492a13",x"4c2b14",x"4d2c15",x"492912",x"462711",x"402411",x"3f2410",x"422511",x"452712",x"482812",x"4a2913",x"4a2913",x"482812",x"492812",x"4c2a14",x"4c2b14",x"492913",x"432410",x"40220e",x"3d220f",x"452611",x"452610",x"40230f",x"40230f",x"452711",x"41230f",x"41230f",x"43240f",x"472711",x"442610",x"422410",x"492811",x"462711",x"492812",x"452711",x"412510",x"482812",x"4a2913",x"4c2b14",x"4c2c14",x"482812",x"482712",x"462711",x"452610",x"472711",x"482812",x"4b2b14",x"4d2c15",x"4e2d15",x"4c2c14",x"4c2b14",x"492913",x"4c2c14",x"4c2c15",x"4b2c15",x"4a2a13",x"4f2e15",x"502f16",x"4a2a14",x"4b2a13",x"472812",x"4b2b15",x"482812",x"4c2b14",x"4a2a13",x"502f16",x"512f16",x"502f17",x"4a2913",x"462711",x"4b2b14",x"4f2d16",x"4c2c15",x"4b2b14",x"462711",x"482812",x"4a2a14",x"4a2a13",x"482913",x"482812",x"492913",x"4b2b14",x"4f2d15",x"4e2d16",x"4d2d15",x"4a2a14",x"4d2c15",x"502e16",x"492a14",x"4e2d15",x"472711",x"462711",x"452610",x"462711",x"472811",x"462811",x"4b2c12",x"512f15",x"42250f",x"000000",x"000000",x"000000",x"000000",x"000000",x"665143",x"665143",x"5e4c3f",x"4d433a",x"55473a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"190f08",x"3f362e",x"453c34",x"4d443a",x"4d443a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"2d2d2d",x"323232",x"333333",x"313131",x"333333",x"313131",x"323232",x"000000",x"000000",x"333333",x"333333",x"2f2f2f",x"343434",x"323232",x"484848",x"323232",x"363636",x"363636",x"373737",x"373737",x"363636",x"383838",x"373737",x"393939",x"3a3a3a",x"3d3d3d",x"3c3c3c",x"3c3c3c",x"3a3a3a",x"3b3b3b",x"383838",x"393939",x"3b3b3b",x"3a3a3a",x"3b3b3b",x"3c3c3c",x"3d3d3d",x"404040",x"414141",x"434343",x"434343",x"444444",x"454545",x"434343",x"404141",x"3f3f3f",x"3f3f3f",x"3c3c3c",x"3c3c3c",x"3a3a3a",x"3e3e3e",x"383838",x"3c3c3c",x"3d3d3d",x"404040",x"454545",x"434343",x"404040",x"444444",x"434343",x"484848",x"4a4a4a",x"454545",x"424242",x"4e4e4e",x"414141",x"444444",x"4a4a4a",x"414141",x"323232",x"444444",x"444444",x"424242",x"3f3f3f",x"4a4a4a",x"313131",x"545454",x"292929",x"575757",x"3c3c3c",x"343434",x"3d3d3d",x"434343",x"464646",x"424242",x"434343",x"464646",x"474747",x"474747",x"3b3b3b",x"414141",x"464646",x"454545",x"464646",x"454545",x"3f3f3f",x"3d3d3d",x"3e3e3e",x"303030",x"3f3f3f",x"313131",x"414141",x"3f3f3f",x"444444",x"4a4a4a",x"4b4b4b",x"494949",x"464646",x"4e4e4e",x"4d4d4d",x"545454",x"4d4d4d",x"595959",x"565656",x"555555",x"585858",x"464646",x"494949",x"535353",x"4b4b4b",x"4b4b4b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3c281b",x"3c281b",x"361e0c",x"331c0c",x"3a200e",x"301a0b",x"251509",x"201208",x"2f1a0b",x"341e0d",x"150e07",x"3a210f",x"412611",x"442712",x"432712",x"452813",x"452813",x"432712",x"422612",x"452812",x"432612",x"422511",x"3f2411",x"3a200e",x"3f2310",x"412612",x"402411",x"3e2310",x"442712",x"432712",x"452813",x"482913",x"432711",x"402410",x"422611",x"452712",x"432611",x"402511",x"412511",x"3f230f",x"3c210e",x"3b200e",x"3d220f",x"3e220f",x"412411",x"412411",x"412511",x"3f2511",x"402410",x"3c210f",x"3a200e",x"3a200e",x"432611",x"432611",x"442711",x"462813",x"442712",x"462913",x"432611",x"3f230f",x"3e230f",x"3b200e",x"3d210e",x"3b210e",x"391f0d",x"3c210f",x"462812",x"462913",x"442711",x"422410",x"3a1f0d",x"3e230f",x"3d210e",x"3a200d",x"3b200e",x"3c220f",x"3a200e",x"3f2310",x"3a210f",x"3c210f",x"341d0c",x"2b180a",x"2b180a",x"2a180a",x"2d190b",x"150e07",x"331c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"221810",x"221810",x"261a11",x"291b10",x"2c1b11",x"2a190d",x"28190e",x"1d130a",x"180f08",x"361e0d",x"382111",x"482a15",x"472a15",x"412714",x"3c2211",x"442714",x"3b2212",x"160f07",x"3b2211",x"402411",x"412411",x"422613",x"432511",x"442610",x"462711",x"422510",x"442611",x"482812",x"452712",x"472912",x"4a2a13",x"452711",x"432511",x"3f230f",x"422410",x"412410",x"412410",x"432511",x"482913",x"4c2c14",x"4c2c15",x"4e2e15",x"472913",x"482913",x"492914",x"4a2a13",x"4d2c15",x"4d2d15",x"4d2d15",x"4a2a14",x"452712",x"452611",x"462712",x"432511",x"4a2a14",x"472812",x"502f17",x"523118",x"4c2d15",x"492913",x"452711",x"4c2c14",x"4a2a14",x"482914",x"4b2b14",x"482812",x"482812",x"4a2a14",x"462712",x"452712",x"482812",x"442711",x"462812",x"4f2e16",x"512f17",x"502f16",x"4d2c14",x"4c2b15",x"4b2b14",x"4e2d15",x"4d2c15",x"472712",x"452711",x"472812",x"492812",x"492812",x"472711",x"492812",x"4b2b14",x"4c2b14",x"492a13",x"4c2b14",x"4d2c15",x"492912",x"462711",x"402411",x"3f2410",x"422511",x"452712",x"482812",x"4a2913",x"4a2913",x"482812",x"492812",x"4c2a14",x"4c2b14",x"492913",x"432410",x"40220e",x"3d220f",x"452611",x"452610",x"40230f",x"40230f",x"452711",x"41230f",x"41230f",x"43240f",x"472711",x"442610",x"422410",x"492811",x"462711",x"492812",x"452711",x"412510",x"482812",x"4a2913",x"4c2b14",x"4c2c14",x"482812",x"482712",x"462711",x"452610",x"472711",x"482812",x"4b2b14",x"4d2c15",x"4e2d15",x"4c2c14",x"4c2b14",x"492913",x"4c2c14",x"4c2c15",x"4b2c15",x"4a2a13",x"4f2e15",x"502f16",x"4a2a14",x"4b2a13",x"472812",x"4b2b15",x"482812",x"4c2b14",x"4a2a13",x"502f16",x"512f16",x"502f17",x"4a2913",x"462711",x"4b2b14",x"4f2d16",x"4c2c15",x"4b2b14",x"462711",x"482812",x"4a2a14",x"4a2a13",x"482913",x"482812",x"492913",x"4b2b14",x"4f2d15",x"4e2d16",x"4d2d15",x"4a2a14",x"4d2c15",x"502e16",x"492a14",x"4e2d15",x"472711",x"462711",x"452610",x"462711",x"472811",x"462811",x"4b2c12",x"512f15",x"42250f",x"42250f",x"000000",x"000000",x"000000",x"000000",x"5f4b3e",x"5f4b3e",x"594538",x"484037",x"4d4339",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3b322a",x"413931",x"4a4037",x"4a4037",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"2f2f2f",x"2d2d2d",x"323232",x"333333",x"313131",x"333333",x"313131",x"323232",x"2b2b2b",x"333333",x"2f2f2f",x"2e2e2e",x"3a3a3a",x"313131",x"343434",x"2f2f2f",x"3a3a3a",x"383838",x"343434",x"353535",x"333333",x"3b3b3b",x"393939",x"2a2a2a",x"3e3e3e",x"3b3b3b",x"3e3e3e",x"3b3b3b",x"3b3b3b",x"3d3d3d",x"373737",x"393939",x"3a3a3b",x"3b3b3b",x"393939",x"383838",x"3e3e3e",x"3b3b3b",x"414141",x"464646",x"454545",x"535353",x"5a5a5a",x"5d5d5d",x"5e5e5e",x"5b5b5b",x"545454",x"4a4a4a",x"424242",x"45362d",x"333333",x"323232",x"373737",x"3b3b3b",x"4e4e4e",x"565656",x"5d5d5d",x"646464",x"636262",x"676767",x"636363",x"686868",x"5d5d5c",x"616161",x"5d5d5d",x"555555",x"4f4f4f",x"4b4b4b",x"525252",x"595959",x"5e5e5e",x"616161",x"686868",x"5e5e5e",x"5b5b5b",x"4b4b4b",x"414141",x"212121",x"444444",x"454545",x"383838",x"414141",x"494949",x"565656",x"585858",x"5b5b5b",x"5e5e5e",x"616161",x"5a5a5a",x"616160",x"666665",x"626262",x"595858",x"666666",x"5c5c5c",x"4c4c4c",x"3d3d3d",x"3c3c3c",x"383838",x"3d3d3d",x"3a3a3a",x"373737",x"404040",x"383838",x"424242",x"4f4f4f",x"565656",x"585858",x"525252",x"565656",x"565656",x"575757",x"575757",x"5b5a5a",x"5c5c5c",x"595959",x"555555",x"5c5c5c",x"5e5e5e",x"515151",x"4e4e4e",x"4e4e4e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3b281b",x"3b281b",x"3d220f",x"2d190b",x"3b210e",x"2e1a0b",x"2f1a0b",x"2f1b0b",x"2d190b",x"2a180a",x"150e07",x"341c0c",x"331c0b",x"361d0c",x"381e0d",x"3b200d",x"3b200e",x"3d220f",x"412510",x"3f2410",x"3e230f",x"3a200e",x"371e0d",x"351d0c",x"321b0b",x"3f2310",x"39200e",x"39200e",x"3e230f",x"3b210e",x"3d220f",x"412410",x"3e230f",x"3e230f",x"3c210f",x"3b200e",x"3a200e",x"3e220f",x"3e220f",x"3e230f",x"3d220f",x"3d210f",x"3d210e",x"3d220f",x"3d220f",x"3e220f",x"391f0e",x"3a200e",x"3b200e",x"3d230f",x"412511",x"3e230f",x"3f230f",x"3d220f",x"432611",x"3e230f",x"412410",x"412410",x"3f230f",x"412310",x"402410",x"402510",x"412410",x"3f220f",x"3c210f",x"412410",x"412511",x"402410",x"3f2410",x"40230f",x"3e230f",x"381e0d",x"391f0d",x"3b200e",x"3f2310",x"3c210f",x"3a1f0d",x"3c210e",x"361e0d",x"3d220f",x"2f1a0b",x"2c180a",x"2e1a0b",x"241509",x"251509",x"150e07",x"361d0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1108",x"1b1108",x"1e1308",x"1e1308",x"1d1308",x"1c1208",x"221608",x"191007",x"1f1408",x"1e1308",x"191007",x"181007",x"150e07",x"1a1107",x"1b1108",x"160f07",x"191007",x"1c1208",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"000000",x"000000",x"000000",x"231911",x"231911",x"271a11",x"2c1b10",x"2d1c0f",x"2e1b0f",x"29190e",x"22140b",x"191008",x"361e0d",x"4e3f35",x"1a130c",x"19120b",x"19130c",x"1a130c",x"1a130c",x"1a130c",x"4b2b14",x"492813",x"4d2b15",x"482712",x"4e2c14",x"4c2a12",x"472711",x"4b2912",x"4b2911",x"482711",x"4f2c13",x"462611",x"482811",x"482812",x"482811",x"4b2913",x"432510",x"4e2c14",x"4c2a13",x"482812",x"432410",x"442510",x"43240f",x"452712",x"4a2a13",x"4c2b13",x"4c2b13",x"4a2913",x"442611",x"4c2913",x"422511",x"422511",x"40230f",x"432510",x"472811",x"452611",x"482811",x"43250f",x"42240f",x"40230f",x"452610",x"43250f",x"482710",x"452610",x"462711",x"4b2913",x"4e2b14",x"4c2b13",x"40230f",x"422410",x"3e210f",x"41230f",x"492813",x"472710",x"482811",x"462712",x"482811",x"482812",x"4a2913",x"4a2912",x"4a2912",x"492912",x"452610",x"43240f",x"4b2a13",x"4c2b13",x"4d2b13",x"4c2a13",x"4a2911",x"492811",x"4c2a13",x"472811",x"482812",x"422510",x"482811",x"472711",x"4f2d14",x"482812",x"4c2b14",x"472712",x"4a2913",x"4e2d15",x"4e2b13",x"4d2b14",x"4c2a12",x"4f2d14",x"4d2a12",x"4e2c13",x"522e15",x"522e15",x"4a2912",x"4c2913",x"482912",x"563116",x"512d15",x"4d2b14",x"4c2a13",x"4e2c14",x"45250f",x"452610",x"4a2811",x"502d14",x"492812",x"40230f",x"4e2b13",x"462610",x"502c14",x"472811",x"45250f",x"4b2811",x"4b2912",x"4a2812",x"482711",x"452510",x"492811",x"482811",x"4b2912",x"472711",x"502d14",x"4f2d15",x"532f16",x"4c2b13",x"452610",x"472711",x"452510",x"4e2d14",x"4c2b13",x"492912",x"4f2d14",x"4c2b13",x"512d14",x"4e2b14",x"512d15",x"4f2d15",x"502c14",x"4d2b14",x"4f2c13",x"4c2a13",x"4e2b12",x"4b2811",x"482711",x"43250f",x"44250f",x"452610",x"432410",x"452610",x"4b2912",x"4a2913",x"4b2b13",x"4e2c14",x"472711",x"3f230f",x"442510",x"42220f",x"4c2a13",x"4a2911",x"4a2913",x"522e14",x"482812",x"472811",x"4a2913",x"482812",x"4b2a12",x"4a2912",x"4c2a12",x"482811",x"472811",x"4c2a13",x"4d2b13",x"4b2a12",x"502d14",x"462711",x"462711",x"000000",x"000000",x"000000",x"000000",x"381d0d",x"381d0d",x"513b2d",x"2e2720",x"4d433a",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"150e07",x"150e07",x"150e07",x"150e07",x"292019",x"3e362e",x"4b4238",x"4b4238",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"2f2f2f",x"313131",x"333333",x"333333",x"313131",x"323232",x"323232",x"323232",x"303030",x"333333",x"313131",x"2f2f2f",x"313131",x"303030",x"313030",x"303030",x"323232",x"353535",x"303030",x"313131",x"414141",x"333333",x"3b3b3b",x"353535",x"3b3b3b",x"3b3b3c",x"3f3f3f",x"424343",x"3d3d3d",x"3a3a3a",x"3d3d3d",x"383838",x"3a3a3a",x"323232",x"383838",x"3a3a3a",x"3c3c3c",x"404040",x"4b4b4b",x"5d5d5d",x"545454",x"555454",x"484645",x"4e4945",x"635d58",x"6d6761",x"625e5a",x"5a5653",x"3f3f3f",x"3a3a3a",x"333333",x"333333",x"313131",x"333333",x"2c2c2c",x"655f59",x"65605b",x"676059",x"655f59",x"65605a",x"69635d",x"68615b",x"6a645f",x"6b655f",x"716b66",x"6c6761",x"6f6a64",x"746e68",x"65605c",x"67635e",x"65605b",x"635f5a",x"65605a",x"69635d",x"5c5c5b",x"5a5a5a",x"575757",x"4f4f4f",x"343434",x"393939",x"323232",x"343434",x"323232",x"534e4a",x"625c56",x"635e59",x"635f5a",x"645f5a",x"6a655f",x"6b6661",x"696460",x"67635e",x"67615c",x"6a635e",x"65605b",x"535353",x"676767",x"4e4e4e",x"3a3a3a",x"313131",x"373737",x"363636",x"343434",x"3e3e3e",x"2f2f2f",x"625c56",x"58534e",x"3c3a38",x"424241",x"4c4c4c",x"595959",x"575757",x"565656",x"656565",x"5a5a5a",x"434241",x"67625e",x"635f5c",x"585756",x"525252",x"535353",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482e1d",x"482e1d",x"412410",x"321c0c",x"3b220f",x"150e07",x"38200f",x"3a210f",x"150e07",x"2c180a",x"150e07",x"3a200e",x"3b200e",x"3c210f",x"3c210e",x"3f230f",x"422510",x"422510",x"3f230f",x"3c210e",x"3d210e",x"3c210f",x"3a200e",x"341c0c",x"341c0c",x"3d210e",x"452811",x"452712",x"3f240f",x"40240f",x"3e230f",x"422511",x"412410",x"412510",x"432712",x"452812",x"432612",x"422611",x"402410",x"3c210e",x"3d2310",x"3f230f",x"402510",x"402410",x"412410",x"41240f",x"3e230f",x"422510",x"432712",x"412510",x"432711",x"442813",x"472913",x"432712",x"412511",x"432711",x"432611",x"412410",x"402410",x"412611",x"462813",x"462812",x"432510",x"3d210e",x"3a200d",x"3c210e",x"412410",x"442711",x"452712",x"462812",x"442711",x"422510",x"3d220f",x"432611",x"3b200e",x"3b200d",x"361d0c",x"351c0c",x"2f1a0b",x"371e0d",x"150e07",x"2b180a",x"301a0b",x"150e07",x"221409",x"150e07",x"3a200e",x"150e07",x"4b2b13",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1108",x"1b1108",x"1e1308",x"1e1308",x"1d1308",x"1c1208",x"221608",x"191007",x"1f1408",x"1e1308",x"191007",x"181007",x"150e07",x"1a1107",x"1b1108",x"160f07",x"191007",x"1c1208",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"29180b",x"000000",x"000000",x"221810",x"221810",x"281b11",x"2e1d11",x"2f1d11",x"2e1c0f",x"2a1a0e",x"24160b",x"1a1008",x"371f0e",x"463a30",x"482a15",x"472a15",x"3d2413",x"412613",x"422613",x"422613",x"3e2210",x"3a1f0f",x"3a1f0e",x"3b200f",x"3c210f",x"3d220f",x"391e0d",x"381e0c",x"381e0d",x"3b200e",x"3d220f",x"432511",x"3e230f",x"3e2310",x"3f2310",x"40230f",x"40230f",x"402410",x"3f240f",x"402410",x"40230f",x"422611",x"3d220f",x"3b220f",x"3c220f",x"3b210f",x"3d2310",x"3b210f",x"38200e",x"3b210f",x"3d220f",x"3c220f",x"3e2310",x"412511",x"3e2310",x"381f0e",x"351d0d",x"371e0d",x"3a200e",x"40240f",x"3f230f",x"3e220f",x"3e220f",x"3e230f",x"3e220f",x"3d210e",x"3b200e",x"3a200e",x"3a200e",x"381f0d",x"331b0b",x"351d0c",x"371e0d",x"402510",x"3e2310",x"3b210f",x"3b210f",x"3d220f",x"402410",x"412410",x"3c220f",x"442712",x"432712",x"402511",x"432611",x"402310",x"3f230f",x"462812",x"412410",x"442711",x"432611",x"402310",x"41240f",x"412510",x"442711",x"452712",x"422511",x"452813",x"422611",x"412511",x"432712",x"402410",x"432711",x"412510",x"422410",x"432611",x"472913",x"452812",x"432611",x"432510",x"3d210e",x"3e210e",x"3a200e",x"422510",x"452712",x"462812",x"442611",x"452712",x"412410",x"3f2310",x"3f2410",x"3c210e",x"381e0d",x"391f0c",x"3b1f0d",x"3c200d",x"3b200d",x"422611",x"391f0d",x"3a1f0d",x"381d0c",x"3a1f0e",x"3e220f",x"3f240f",x"402410",x"3e220f",x"402410",x"3d220f",x"381f0d",x"3d220f",x"3f2410",x"3e220f",x"3e220f",x"442611",x"3c210f",x"462813",x"432712",x"412411",x"432611",x"422511",x"452711",x"412410",x"412411",x"412411",x"452712",x"472913",x"432611",x"422611",x"3f230f",x"3e220e",x"41230f",x"40240f",x"40230f",x"40230f",x"40230f",x"402410",x"422510",x"412410",x"3f230f",x"3f220f",x"3a200e",x"41240f",x"391e0d",x"391f0d",x"3b200e",x"412510",x"412511",x"402410",x"412410",x"412410",x"412411",x"402410",x"422511",x"452812",x"472913",x"422711",x"442712",x"412411",x"432510",x"422511",x"422511",x"4a2913",x"4a2913",x"000000",x"000000",x"000000",x"000000",x"371c0c",x"371c0c",x"4f3728",x"272019",x"4d433a",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"150e07",x"150e07",x"150e07",x"170f07",x"22170e",x"3a3129",x"4c4338",x"4c4338",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"333333",x"343434",x"313131",x"343434",x"323232",x"3c3c3c",x"454546",x"5a5a5a",x"3c3c3c",x"323232",x"333333",x"2f2f2f",x"303030",x"313131",x"2f2f2f",x"343434",x"333333",x"434343",x"323232",x"545454",x"444444",x"3f3f40",x"393939",x"404040",x"434343",x"424242",x"454545",x"3f3f3f",x"414141",x"393939",x"373737",x"313131",x"313131",x"383838",x"3d3d3d",x"424242",x"525252",x"60605f",x"4a4a4a",x"4e4e4e",x"4b4b4a",x"484645",x"4e4945",x"635d58",x"323232",x"2f2f2f",x"333333",x"313131",x"313131",x"333333",x"2f2f2f",x"303030",x"313131",x"333333",x"2f2f2f",x"323232",x"333333",x"655f59",x"65605a",x"69635d",x"68615b",x"6a645f",x"6b655f",x"706a64",x"706b65",x"6f6a64",x"746e68",x"6d6862",x"66615b",x"635e58",x"645e59",x"65605a",x"69635d",x"5c5c5b",x"545353",x"515050",x"4a4a4a",x"4f4f4f",x"323232",x"3f3f3f",x"373737",x"404040",x"333333",x"2d2d2d",x"323232",x"333333",x"3f3f3f",x"6a655f",x"6b6661",x"696460",x"67635e",x"67615c",x"6a635e",x"575654",x"4d4d4d",x"3f3f3f",x"3a3a3a",x"636362",x"4b4b4b",x"424242",x"404040",x"595959",x"565656",x"373737",x"313131",x"524d49",x"41403f",x"434342",x"494949",x"4b4a4a",x"585858",x"656565",x"515050",x"3f3f3e",x"383838",x"67625e",x"65615b",x"5c5956",x"525252",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3e291b",x"3e291b",x"3e230f",x"38200e",x"3f2310",x"351e0e",x"371e0d",x"30190a",x"2f1a0b",x"371f0d",x"231409",x"361d0c",x"331c0b",x"321a0a",x"31190a",x"341b0b",x"371d0b",x"361c0b",x"381e0d",x"3f220f",x"40230f",x"3b200e",x"371e0d",x"341c0b",x"341c0c",x"381e0c",x"371d0c",x"371e0d",x"371e0c",x"3a1f0d",x"3b200d",x"361d0c",x"361d0c",x"341c0c",x"381e0c",x"371e0c",x"371d0c",x"391f0d",x"351c0c",x"331c0c",x"381f0d",x"3b200e",x"391f0d",x"391f0d",x"381e0c",x"361d0c",x"3a200e",x"3c210e",x"3b200e",x"3f220f",x"3c210e",x"3b200e",x"3b200e",x"3e220f",x"391f0d",x"381e0d",x"371e0c",x"351b0b",x"341c0b",x"361d0c",x"381e0c",x"361d0c",x"361d0c",x"341b0b",x"351c0b",x"361c0c",x"331a0b",x"321a0b",x"33190a",x"321a0b",x"30190a",x"361d0c",x"371d0c",x"351b0b",x"331b0b",x"3a200e",x"3d220f",x"3b210f",x"371f0d",x"3e220f",x"311b0c",x"371f0e",x"3b210f",x"341d0d",x"361e0d",x"150e07",x"3c210f",x"3b200e",x"492812",x"452711",x"432712",x"432711",x"432611",x"432611",x"452812",x"3e220f",x"3e220f",x"432611",x"422510",x"402310",x"3e220e",x"3f230f",x"3b210f",x"412511",x"3e220f",x"3f2310",x"412411",x"422511",x"3d220f",x"351c0c",x"371d0d",x"351d0d",x"3b200e",x"391f0d",x"341c0b",x"351c0b",x"321a0a",x"341b0b",x"341b0b",x"361c0b",x"371d0c",x"3c210e",x"40230f",x"3f230f",x"3c220e",x"3b200d",x"391f0c",x"381e0c",x"381e0c",x"39200c",x"3a200d",x"381f0c",x"39200d",x"381e0c",x"3a200d",x"39200d",x"391f0c",x"3b200d",x"361d0c",x"371e0d",x"331c0c",x"351c0c",x"341c0c",x"351d0d",x"371e0d",x"371e0d",x"371e0c",x"381e0c",x"3b200d",x"3a200e",x"3a200e",x"3b210e",x"391f0e",x"3f220f",x"391f0d",x"422410",x"150e07",x"170f07",x"170f07",x"000000",x"000000",x"241911",x"241911",x"291b12",x"2f1e11",x"311e10",x"301c0f",x"2d1c0f",x"2b190c",x"1b1108",x"371f0d",x"483f36",x"392011",x"361f0f",x"3a2011",x"361f0f",x"321c0f",x"3e2311",x"3f2512",x"3e2311",x"402411",x"422612",x"3b200e",x"3f230f",x"422511",x"3d220f",x"402410",x"3b210e",x"3e230f",x"3d220f",x"3e230f",x"3f230f",x"3e230f",x"3c210e",x"422611",x"412510",x"422511",x"3d220f",x"3b200e",x"422611",x"3f2410",x"381f0e",x"3b200e",x"391f0d",x"3f2410",x"402410",x"38200e",x"381f0e",x"3a200f",x"3c210f",x"3c210f",x"381f0d",x"311a0b",x"351d0c",x"3a200e",x"351d0c",x"351c0b",x"351c0c",x"331a0b",x"321a0a",x"321a0b",x"30190b",x"341a0b",x"361e0c",x"3c210e",x"381f0e",x"361e0d",x"351d0c",x"341c0b",x"331b0b",x"321b0b",x"341c0c",x"361d0c",x"341c0c",x"351d0c",x"361d0c",x"351c0c",x"351d0c",x"381e0d",x"371d0c",x"341c0c",x"371e0c",x"331c0c",x"391e0d",x"3a1f0d",x"3d210e",x"3a200e",x"3a200e",x"3b200d",x"381d0c",x"3a1f0d",x"3d210e",x"3d210e",x"3e220f",x"3d220f",x"3e220f",x"3e220f",x"3f220f",x"3e220f",x"3b200e",x"3a1f0d",x"351c0b",x"331a0b",x"341b0b",x"381e0d",x"371e0c",x"371d0c",x"381d0c",x"361c0b",x"371c0c",x"351c0c",x"351b0b",x"371c0b",x"331a0b",x"341b0b",x"371c0c",x"3b200d",x"371d0c",x"321a0b",x"371d0c",x"3a200e",x"422510",x"40240f",x"3e230f",x"3e220f",x"3f230f",x"422510",x"3f230f",x"3e220f",x"3a200e",x"3f220f",x"3e220f",x"3d220f",x"3f220f",x"3c210f",x"371e0d",x"432611",x"422611",x"412510",x"422511",x"391f0d",x"3d220f",x"412410",x"3e220f",x"3d210f",x"3e220f",x"40230f",x"3f2310",x"412410",x"3f230f",x"432611",x"432611",x"422611",x"3f230f",x"361c0c",x"3a1f0d",x"3e220f",x"3c210e",x"3a1f0d",x"361c0c",x"341c0b",x"351b0b",x"331a0a",x"351c0b",x"371d0c",x"371d0c",x"3b210e",x"3d210e",x"3d210e",x"3c210e",x"371d0c",x"371d0c",x"381e0c",x"371d0c",x"381f0d",x"3b200d",x"3a1f0d",x"3b200e",x"381e0d",x"3a1f0d",x"3b200d",x"3a1f0d",x"391f0d",x"331c0c",x"381f0d",x"391f0d",x"381e0d",x"3b200e",x"3c210e",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"391e0d",x"391e0d",x"513423",x"2a2119",x"4f463d",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"160e07",x"150e07",x"150e07",x"150e07",x"27180d",x"2d261f",x"4b4238",x"4b4238",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"3c3c3c",x"3a3a3a",x"3f3f3f",x"383838",x"3e3e3e",x"4a4a4a",x"4e4e4e",x"535353",x"5f5f5f",x"3e3e3e",x"313131",x"303030",x"323232",x"323232",x"333333",x"333333",x"3a3a3a",x"393939",x"3e3f3f",x"323232",x"4e4e4e",x"2e2e2e",x"424242",x"3e3e3e",x"404040",x"4b4b4b",x"535353",x"5e5e5e",x"5f5f5f",x"5b5b5b",x"515151",x"484848",x"424242",x"3d3d3d",x"474747",x"505050",x"5b5b5b",x"5e5e5e",x"414141",x"4c4c4c",x"4a4a4a",x"4a4a49",x"000000",x"4c4c4c",x"303030",x"313131",x"303030",x"343434",x"333333",x"313131",x"454545",x"4b4b4b",x"454545",x"4a4a4a",x"4d4d4d",x"424242",x"313131",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"555555",x"515050",x"414141",x"373737",x"4a4a4a",x"3a3a3a",x"3a3a3a",x"434343",x"4b4b4b",x"494949",x"5b5b5b",x"5b5b5b",x"4e4e4e",x"4e4e4e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"484848",x"393939",x"323232",x"303030",x"4f4f4f",x"565656",x"595959",x"696868",x"5f5f5f",x"333333",x"323232",x"000000",x"000000",x"434242",x"4a4a4a",x"4a4949",x"5e5a58",x"696560",x"565453",x"484747",x"3f3f3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452d1e",x"452d1e",x"3e230f",x"3e230f",x"402410",x"412511",x"3e220f",x"3c210f",x"381e0d",x"2c180a",x"2c180a",x"331b0b",x"381e0d",x"3b200e",x"39200e",x"3a200e",x"3b200e",x"3d220f",x"3d220f",x"3d220f",x"40240f",x"3c210e",x"3d210e",x"3b200e",x"3a200e",x"3e220f",x"402410",x"3f230f",x"3c210f",x"3e220f",x"391f0d",x"391f0d",x"3a200e",x"412510",x"422611",x"432711",x"422611",x"442712",x"422611",x"3d220f",x"3c210f",x"422511",x"3f2310",x"381e0d",x"3c210e",x"391f0d",x"3d220f",x"381f0d",x"3c210f",x"3c210e",x"3d210e",x"3a200d",x"371d0c",x"381e0c",x"3a1f0d",x"361c0c",x"361c0c",x"2e1609",x"30180a",x"381e0c",x"3e220f",x"3b200e",x"3b200d",x"3b200e",x"3a1f0d",x"3c210e",x"3d220f",x"3d210f",x"3b200e",x"3a200e",x"3b200e",x"3a200e",x"381f0e",x"3f2410",x"3e220f",x"3c210f",x"3b210f",x"3c220f",x"3a210e",x"402410",x"3f2310",x"3f2310",x"3c210f",x"371e0d",x"391f0d",x"2b180a",x"3d210e",x"3f230f",x"4b2b13",x"432611",x"412410",x"3f230f",x"472813",x"442611",x"432611",x"462812",x"452813",x"452712",x"432611",x"452812",x"452812",x"462913",x"402511",x"2c190b",x"1a1008",x"201309",x"24150a",x"26160a",x"26160a",x"26160a",x"27160a",x"241409",x"251509",x"251509",x"231409",x"251509",x"251509",x"221409",x"211309",x"241509",x"1d1108",x"29170a",x"241509",x"261609",x"2b190b",x"2a190a",x"2f1c0b",x"2c1a0a",x"2f1c0b",x"241509",x"211309",x"241509",x"231409",x"231409",x"1f1208",x"25150a",x"25160a",x"24150a",x"211409",x"241609",x"24150a",x"231409",x"211309",x"331c0c",x"3e230f",x"3b200e",x"3a200e",x"3a200e",x"3c210e",x"371d0c",x"3e220f",x"3d210f",x"3a200e",x"3a200d",x"371e0d",x"3c200d",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"241910",x"241910",x"2a1c11",x"311e12",x"341f11",x"321e0f",x"321e10",x"2a190c",x"1c1108",x"3a210f",x"4d4034",x"3f2412",x"3d2312",x"412613",x"3d2412",x"3d2312",x"412614",x"422512",x"412511",x"3c2210",x"412410",x"3d230f",x"422611",x"3e220f",x"391f0e",x"361e0d",x"391f0d",x"391f0e",x"3e220f",x"40230f",x"422511",x"422511",x"3f2410",x"432611",x"412511",x"3f230f",x"3e2310",x"432711",x"442712",x"3e2310",x"452711",x"432712",x"432712",x"422712",x"3f2411",x"39200e",x"3e230f",x"3a210f",x"3d230f",x"3c210f",x"3e230f",x"3c210e",x"391f0d",x"391f0d",x"361c0c",x"381d0d",x"391f0d",x"3b200e",x"361e0d",x"3a200e",x"3b200e",x"39200e",x"3a200e",x"39200e",x"351d0d",x"381f0d",x"381f0d",x"381f0d",x"3b200e",x"3b210e",x"3d230f",x"3d220f",x"3b210e",x"3d210f",x"381f0d",x"391f0d",x"3b210e",x"412510",x"402511",x"412511",x"402511",x"452712",x"432611",x"3e220f",x"3e220f",x"3d220f",x"412510",x"39200e",x"3d220e",x"3c210e",x"391f0d",x"3c210e",x"3c210e",x"3b200e",x"3c210e",x"3b200d",x"391f0d",x"361d0c",x"381e0d",x"361c0c",x"331a0b",x"2e1709",x"31190a",x"3b200e",x"3b210e",x"3c200e",x"3b200e",x"3b200d",x"3b200d",x"381f0d",x"3a200d",x"3a200e",x"3e220f",x"3d210e",x"3c210f",x"402310",x"3e230f",x"432611",x"3e230f",x"3a210f",x"3f240f",x"3f240f",x"3f2410",x"412511",x"432611",x"412411",x"3e220f",x"3b200e",x"3d210e",x"3b200e",x"3c210e",x"3f230f",x"412410",x"412411",x"3f2410",x"3e230f",x"452813",x"3f230f",x"412511",x"412611",x"422612",x"432611",x"432611",x"452812",x"472913",x"492a14",x"452812",x"412410",x"412410",x"452712",x"432611",x"442711",x"422510",x"422410",x"3e210e",x"3c200d",x"3b200d",x"3a1f0d",x"3b1f0d",x"3c210e",x"432510",x"412410",x"3d210e",x"3e220f",x"3d220f",x"3f230f",x"3c210e",x"381f0d",x"3d210e",x"3b200e",x"3c210e",x"3e220f",x"3f230f",x"3f2310",x"412410",x"3e220f",x"3e220f",x"3d210e",x"3c210e",x"452711",x"472913",x"472913",x"452712",x"432611",x"432611",x"3e230f",x"3e230f",x"422510",x"4a2913",x"4a2913",x"000000",x"000000",x"000000",x"000000",x"381e0d",x"381e0d",x"4f321f",x"2d221a",x"4d443b",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"150e07",x"150e07",x"150e07",x"190f08",x"2a190c",x"2c2118",x"494037",x"494037",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"545454",x"484848",x"4b4b4b",x"414141",x"494949",x"575757",x"545454",x"5b5b5b",x"626262",x"484848",x"313131",x"313131",x"333333",x"323232",x"383838",x"3d3d3d",x"434343",x"434343",x"474747",x"454545",x"4e4e4e",x"4c4c4c",x"474747",x"464646",x"555555",x"666666",x"5c5c5c",x"565656",x"63615e",x"504f4e",x"494949",x"515151",x"585858",x"4c4c4c",x"575656",x"5e5e5e",x"424242",x"393939",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"565656",x"565656",x"636363",x"646464",x"535353",x"595959",x"575757",x"535353",x"525252",x"5f5f5f",x"565656",x"5c5b5b",x"5f5f5e",x"606060",x"3a3a3a",x"3a3a3a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434343",x"434343",x"313131",x"303030",x"3b3b3b",x"313131",x"383838",x"4c4c4c",x"565656",x"555555",x"414141",x"464646",x"464646",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4a4a",x"4a4a4a",x"626261",x"60605f",x"606060",x"666666",x"5f5f5f",x"545454",x"373737",x"363636",x"000000",x"000000",x"000000",x"000000",x"535251",x"5e5a58",x"696560",x"565453",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"463020",x"463020",x"462813",x"432712",x"27160a",x"442712",x"3f2410",x"422611",x"3f2310",x"150e07",x"351d0c",x"39200d",x"3a1f0d",x"3e220e",x"3c210e",x"391f0e",x"3a200e",x"391f0e",x"3d210f",x"3f2410",x"412511",x"422511",x"412511",x"3f2310",x"3a200e",x"371e0d",x"351c0b",x"351c0c",x"391e0d",x"391f0d",x"361d0c",x"351c0c",x"361d0c",x"381e0d",x"351c0c",x"371e0c",x"361e0d",x"3f230f",x"422611",x"3c220f",x"402510",x"412511",x"442712",x"412511",x"3f240f",x"3f230f",x"3f230f",x"3f230f",x"3c210e",x"432611",x"412511",x"40230f",x"40240f",x"402410",x"432611",x"412411",x"402410",x"412510",x"412410",x"462711",x"3f230f",x"3e220f",x"3b200e",x"381f0d",x"371e0d",x"391f0d",x"3a1f0d",x"371e0d",x"391f0d",x"3c210e",x"3a200e",x"3a200e",x"3e220f",x"3f230f",x"412510",x"3f240f",x"402310",x"3b210e",x"371e0d",x"2c190b",x"381f0d",x"3d220f",x"402511",x"412511",x"150e07",x"2d1a0b",x"422511",x"512e15",x"321d0c",x"361e0d",x"351e0e",x"36200e",x"3a2210",x"37200f",x"351e0e",x"341d0d",x"341d0d",x"371f0e",x"2f1a0b",x"301b0c",x"331d0d",x"37200f",x"38200f",x"361f0e",x"341e0e",x"36200f",x"2f1b0c",x"2a190b",x"211309",x"231509",x"191008",x"1e1208",x"27160a",x"150e07",x"150e07",x"1e1108",x"211309",x"221409",x"221409",x"1a1008",x"150e07",x"150e07",x"25170a",x"251809",x"251809",x"241708",x"2a1a09",x"261809",x"281809",x"150e07",x"150e07",x"191008",x"201208",x"221309",x"150e07",x"1f1208",x"150e07",x"150e07",x"150e07",x"1e1208",x"27160a",x"25160a",x"231509",x"24150a",x"24150a",x"2e1a0b",x"311c0c",x"311b0c",x"2e1a0b",x"2f1b0b",x"2f1a0b",x"311b0c",x"2f1b0c",x"26160a",x"211409",x"301b0c",x"331d0d",x"150e07",x"150e07",x"000000",x"000000",x"241910",x"241910",x"2b1b10",x"322012",x"352011",x"321e10",x"331e10",x"2a190c",x"1d1108",x"371e0d",x"4f4136",x"402413",x"3c2211",x"3d2313",x"3c2312",x"3b2211",x"402613",x"3f2412",x"3f2411",x"3d2210",x"361d0d",x"331c0c",x"3b210e",x"3c220f",x"402410",x"402410",x"462812",x"412511",x"412411",x"432611",x"3f240f",x"422611",x"412511",x"432712",x"422612",x"422611",x"432611",x"3e230f",x"3c230f",x"412511",x"3e220f",x"412410",x"432612",x"452913",x"432712",x"402511",x"412611",x"3a2210",x"3b210f",x"3e2310",x"412511",x"3e2310",x"39200e",x"3b210f",x"3b200e",x"321c0c",x"351d0c",x"3a200d",x"391f0e",x"3c210e",x"331c0c",x"381f0e",x"3a200e",x"3f2410",x"3d2310",x"3b210f",x"3d2310",x"402410",x"3a200e",x"361d0c",x"351c0c",x"361d0c",x"351d0c",x"381f0d",x"341c0b",x"351c0c",x"351c0c",x"351d0c",x"331b0b",x"351c0c",x"3a200e",x"3d220f",x"432611",x"432611",x"3f2410",x"422611",x"3f2411",x"412511",x"402410",x"3f240f",x"402410",x"3f230f",x"3e220f",x"402511",x"422510",x"3e220f",x"3f240f",x"432611",x"422611",x"402410",x"432611",x"432611",x"412410",x"402410",x"3d210f",x"3d210e",x"3d220f",x"3b200e",x"3d210e",x"3a1f0d",x"381f0d",x"391f0d",x"391f0d",x"391f0d",x"391f0d",x"3b200e",x"3f230f",x"402410",x"3d220f",x"3c220f",x"3b210f",x"391f0e",x"391f0d",x"3a1f0d",x"3a200e",x"3e230f",x"422511",x"412511",x"412511",x"412511",x"422611",x"3d2310",x"422510",x"432611",x"3f2410",x"432712",x"442712",x"452813",x"432611",x"402310",x"402410",x"422510",x"3e230f",x"3f230f",x"462813",x"452813",x"482a14",x"462813",x"442712",x"4a2b14",x"422510",x"432611",x"432611",x"442812",x"482912",x"432711",x"40230f",x"3d220e",x"3b200e",x"3b200e",x"3d210e",x"3f230f",x"3a200e",x"3f220f",x"40230f",x"422611",x"412511",x"422611",x"432611",x"452712",x"412410",x"3a200d",x"391e0c",x"381e0c",x"371d0d",x"381f0d",x"381e0c",x"371d0c",x"381e0c",x"361d0c",x"341c0b",x"391f0d",x"3c200e",x"3c210e",x"402410",x"3f2410",x"422611",x"452712",x"482813",x"482813",x"000000",x"000000",x"000000",x"000000",x"3b200d",x"3b200d",x"563721",x"2f2118",x"494037",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"27180c",x"221a13",x"40372f",x"40372f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5d5d5d",x"5d5d5d",x"5b5b5b",x"5e5e5e",x"4c4c4c",x"5c5c5c",x"626262",x"5f5e5e",x"636363",x"626261",x"4d4d4d",x"3d3d3d",x"313131",x"353535",x"434343",x"4c4c4c",x"515151",x"5a5a5a",x"585858",x"595959",x"5a5a5a",x"626262",x"5a5a5a",x"5f5f5f",x"626262",x"6d6d6d",x"5a5a5b",x"575757",x"5a5959",x"63615e",x"464646",x"585858",x"515151",x"616261",x"656565",x"636362",x"626262",x"333333",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"676767",x"676767",x"5a5a5a",x"504f4f",x"656565",x"5d5c5c",x"646363",x"616161",x"606060",x"5c5c5c",x"5f5f5f",x"565655",x"64605d",x"4a4a4a",x"3c3c3c",x"3d3d3d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"585858",x"585858",x"555555",x"525151",x"525252",x"5b5b5b",x"5a5a5a",x"5f5f5f",x"565656",x"323232",x"333232",x"414141",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"616161",x"616161",x"656260",x"605a56",x"67615c",x"6f6c68",x"64615f",x"474645",x"545454",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"453225",x"453225",x"402410",x"3a200e",x"150e07",x"412411",x"412410",x"422611",x"3f2310",x"150e07",x"321c0c",x"39200e",x"381f0d",x"3a200d",x"3d210e",x"3b200d",x"2f1b0c",x"311c0d",x"311c0d",x"321d0e",x"361e0d",x"3f2410",x"3e2310",x"3f2410",x"381f0d",x"38200f",x"3c210f",x"391f0d",x"402410",x"3b200e",x"3a1f0e",x"381f0d",x"371d0c",x"351c0c",x"331b0c",x"391f0d",x"422611",x"3c200e",x"432511",x"3d220f",x"402410",x"412510",x"381e0d",x"3d210e",x"3c210e",x"3b200e",x"3b200e",x"3d210e",x"412410",x"3b200e",x"3f230f",x"3a200e",x"3d210f",x"3f230f",x"3a200e",x"3d210f",x"41240f",x"442611",x"412410",x"442712",x"3f2410",x"412410",x"432511",x"3f2410",x"39200e",x"3a200e",x"3d230f",x"3e230f",x"452712",x"432611",x"3f230f",x"38200e",x"492a14",x"402410",x"402410",x"412411",x"442712",x"3f2410",x"412612",x"150e07",x"432612",x"452914",x"402512",x"432712",x"150e07",x"27170a",x"3b210f",x"522f16",x"412511",x"412511",x"402511",x"3d2310",x"3c210f",x"3f2511",x"402511",x"422611",x"402410",x"402511",x"412511",x"402512",x"3d2411",x"3d230f",x"412511",x"3e230f",x"3c220f",x"361e0d",x"180f07",x"150e07",x"38200e",x"3a210f",x"150e07",x"150e07",x"321c0c",x"150e07",x"150e07",x"2e190b",x"29170a",x"150e07",x"150e07",x"28160a",x"150e07",x"251509",x"281709",x"261709",x"301c0a",x"311c0b",x"2f1c0a",x"1b1108",x"281609",x"150e07",x"150e07",x"1c1108",x"28160a",x"150e07",x"261409",x"1c1108",x"271509",x"29170a",x"2a170a",x"150e07",x"1b1008",x"1f1208",x"1a1008",x"150e07",x"2b180b",x"311b0b",x"331c0c",x"371e0d",x"38200e",x"391f0e",x"39200e",x"3c220f",x"361e0d",x"38200e",x"3a210f",x"321d0d",x"402511",x"150e07",x"150e07",x"000000",x"000000",x"24180f",x"24180f",x"2a1b10",x"331f11",x"341f11",x"331e0f",x"331e10",x"321d0e",x"1f1208",x"341d0c",x"4a3b30",x"4b2c16",x"452915",x"462a16",x"442815",x"3b2312",x"412512",x"432813",x"402513",x"432712",x"442813",x"3b2210",x"422612",x"442713",x"412612",x"442813",x"442813",x"432611",x"422511",x"452812",x"452712",x"462913",x"412511",x"3f2310",x"422611",x"432712",x"452813",x"462812",x"432711",x"412510",x"452913",x"442713",x"432712",x"402410",x"3e2310",x"3b210f",x"3a200e",x"39200e",x"422510",x"3b210f",x"3f2310",x"3d230f",x"3c220f",x"3a210e",x"361f0d",x"381f0e",x"381f0d",x"391f0d",x"351d0c",x"341c0b",x"361d0c",x"341c0c",x"361e0c",x"351d0c",x"371e0d",x"321b0b",x"341c0c",x"341c0c",x"331c0b",x"351c0c",x"321a0b",x"31190a",x"321a0b",x"341c0c",x"361d0c",x"311a0a",x"321a0a",x"331c0b",x"331c0c",x"331b0b",x"331b0b",x"2f1709",x"31190a",x"3c210e",x"3d220f",x"3a200e",x"3c210e",x"381f0d",x"3d210e",x"3d220f",x"3e230f",x"422511",x"412510",x"422511",x"432611",x"452712",x"442712",x"452812",x"432711",x"422510",x"412410",x"3c210e",x"402310",x"432711",x"422611",x"452711",x"422511",x"422611",x"432511",x"432611",x"452712",x"462812",x"462813",x"432712",x"442813",x"452813",x"442712",x"422511",x"402410",x"3f2410",x"402511",x"422612",x"452813",x"462913",x"452813",x"472a14",x"442813",x"472914",x"442813",x"3f2411",x"402410",x"432712",x"432712",x"452812",x"3f2410",x"432611",x"402410",x"452813",x"472913",x"452812",x"452712",x"452712",x"462913",x"472914",x"472913",x"452712",x"3f2310",x"402410",x"3f2410",x"3d220f",x"3f2310",x"412511",x"412511",x"402510",x"422511",x"422510",x"412510",x"402410",x"381f0d",x"3b200d",x"3c210e",x"351d0c",x"391f0d",x"391e0d",x"3c210e",x"341c0c",x"381e0d",x"381f0d",x"361d0c",x"391f0d",x"381e0d",x"361d0c",x"341b0b",x"321a0b",x"341b0b",x"381f0c",x"3a1f0d",x"331b0b",x"32190a",x"351c0c",x"331b0b",x"361d0c",x"361c0c",x"31190a",x"31190a",x"391f0d",x"3b210e",x"3f230f",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"3a200d",x"3a200d",x"53331e",x"302016",x"50473e",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"23180f",x"3c342c",x"3c342c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5b5651",x"5b5651",x"5f5954",x"625b53",x"6c6965",x"6f6a64",x"6e6862",x"69635e",x"605a53",x"645d57",x"76726d",x"6f6a65",x"6f6a64",x"77726d",x"6f6a65",x"76716d",x"79746f",x"6d6966",x"6e6a67",x"6c6864",x"6f6a67",x"76716c",x"6f6c6a",x"6f6c6a",x"6f6c69",x"636363",x"5a5a5a",x"575757",x"000000",x"000000",x"5c5c5c",x"616161",x"636363",x"6c6b69",x"6a6662",x"65615e",x"4a4a4a",x"494949",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"656565",x"4e4e4e",x"4b4a4a",x"4c4b4a",x"565351",x"5d5a58",x"635e59",x"66615c",x"635f5b",x"605c59",x"595653",x"595754",x"4f4e4e",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"5f5f5f",x"626161",x"595856",x"565656",x"5d5c5c",x"4e4d4d",x"5a5a5a",x"5a5a5a",x"464646",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5f5f5e",x"656260",x"605a56",x"746e68",x"6f6c68",x"706a66",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"443226",x"443226",x"402511",x"3c2310",x"412511",x"3f2410",x"3f2411",x"3e220f",x"432612",x"402511",x"1d1108",x"3d220f",x"170f07",x"371e0d",x"311c0c",x"24150a",x"2f1b0c",x"311c0d",x"311c0d",x"321d0e",x"361e0d",x"5f5f5f",x"575757",x"555555",x"636363",x"38200f",x"3c210f",x"391f0d",x"402410",x"3b200e",x"3a1f0e",x"381f0d",x"371d0c",x"351c0c",x"331b0c",x"391f0d",x"422611",x"3c200e",x"432511",x"3d220f",x"402410",x"412510",x"381e0d",x"3d210e",x"3c210e",x"3b200e",x"3b200e",x"3d210e",x"412410",x"3b200e",x"3f230f",x"3a200e",x"3d210f",x"3f230f",x"3a200e",x"3d210f",x"41240f",x"442611",x"412410",x"442712",x"3f2410",x"412410",x"432511",x"3f2410",x"39200e",x"3a200e",x"3d230f",x"3e230f",x"452712",x"432611",x"3f230f",x"311c0c",x"361f0e",x"4d2b14",x"3e2411",x"482711",x"150e07",x"211409",x"3b2311",x"3b210f",x"3e2311",x"38200f",x"3f2411",x"391f0e",x"3d2411",x"150e07",x"3b2210",x"563219",x"472a14",x"442813",x"422612",x"402410",x"3f2410",x"3f2310",x"3c210f",x"39200e",x"3a200e",x"3c210f",x"3d2310",x"3b210f",x"3e230f",x"3f2410",x"402410",x"3d220f",x"3a200e",x"331d0d",x"351d0d",x"391f0e",x"3c220f",x"231409",x"231409",x"39200e",x"2a180b",x"150e07",x"261409",x"2a170a",x"2f1a0b",x"3c210f",x"150e07",x"241509",x"150e07",x"311b0b",x"311b0b",x"150e07",x"150e07",x"150e07",x"5d5449",x"150e07",x"150e07",x"150e07",x"2e1a0b",x"28170a",x"261509",x"311b0b",x"150e07",x"150e07",x"180f07",x"2f1a0b",x"28170a",x"2d190b",x"351d0c",x"381f0d",x"341d0c",x"351d0d",x"2a170a",x"341d0d",x"321c0c",x"331c0c",x"331c0c",x"361e0d",x"361e0d",x"3b210f",x"39200e",x"351e0e",x"3b210f",x"3a210f",x"412511",x"150e07",x"150e07",x"000000",x"000000",x"22180f",x"22180f",x"291a0f",x"342011",x"321d0f",x"311d0f",x"311c0d",x"2f1c0d",x"201309",x"341c0c",x"4a3b2f",x"462915",x"412613",x"3f2412",x"402511",x"3a200f",x"402412",x"442814",x"412613",x"422612",x"402411",x"3f2411",x"442712",x"3f2411",x"422712",x"442813",x"452914",x"412612",x"452813",x"492c15",x"462914",x"482a14",x"402410",x"402410",x"402511",x"3f2410",x"3e220f",x"381f0d",x"3d220f",x"3c210f",x"3e2310",x"402410",x"3e230f",x"3c220f",x"3f2310",x"3f240f",x"3a200e",x"341c0c",x"381f0e",x"3c210f",x"381f0e",x"3e220f",x"391f0e",x"3b210f",x"311b0b",x"301a0b",x"2d170a",x"361d0c",x"3a200e",x"3c220f",x"3d220f",x"341c0c",x"351d0c",x"391f0d",x"3c210f",x"3b210f",x"3a200e",x"3d220f",x"3d220f",x"3c210e",x"3c210e",x"381f0d",x"371f0d",x"351d0c",x"371e0d",x"381f0d",x"391f0d",x"391f0d",x"3c210e",x"3c210e",x"3a200e",x"381e0d",x"391f0d",x"3d210e",x"3a200e",x"371e0d",x"391f0d",x"39200e",x"391f0e",x"3b200e",x"3a200e",x"3d220f",x"3f2310",x"3c210f",x"412411",x"422511",x"432712",x"452812",x"432611",x"422511",x"432712",x"432611",x"3d210e",x"452712",x"472914",x"422511",x"422611",x"452712",x"422611",x"432611",x"432611",x"402410",x"442712",x"422611",x"402410",x"3f2310",x"3e220f",x"3c210f",x"3c210f",x"412611",x"3f2411",x"452812",x"422611",x"452812",x"412511",x"452812",x"402511",x"462914",x"462914",x"442713",x"442713",x"442813",x"462914",x"422712",x"3f2411",x"3f2410",x"402410",x"3b210f",x"412510",x"3f230f",x"3b210e",x"3c210f",x"3f2310",x"422511",x"412511",x"412511",x"3e230f",x"3f2410",x"40240f",x"3f220f",x"422510",x"3b210f",x"3f230f",x"3b200e",x"3a200e",x"3f230f",x"3e220f",x"371d0c",x"331b0b",x"331b0b",x"381f0d",x"422510",x"412511",x"3f230f",x"371d0d",x"351d0c",x"3c210e",x"40240f",x"3d220f",x"402410",x"402310",x"3e220f",x"3e220e",x"3d210e",x"3c210e",x"3b200e",x"361e0d",x"3a200d",x"3c210e",x"3b210e",x"391f0d",x"3b210e",x"3b200e",x"3a200e",x"3c210e",x"3f230f",x"3f220f",x"3d220e",x"40230e",x"40230e",x"000000",x"000000",x"000000",x"000000",x"391f0d",x"391f0d",x"492c18",x"2c1e14",x"4d443b",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"160e07",x"150e07",x"150e07",x"150e07",x"26160a",x"24180e",x"372f27",x"372f27",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"525252",x"525252",x"383838",x"343434",x"484848",x"353535",x"333333",x"323232",x"323232",x"333333",x"323232",x"323232",x"313131",x"313131",x"303030",x"323232",x"333333",x"303030",x"313232",x"363636",x"303030",x"303030",x"343434",x"333333",x"404040",x"3a3a3a",x"313131",x"2f2f2f",x"000000",x"000000",x"323232",x"323232",x"333333",x"343434",x"313131",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"323232",x"323232",x"323232",x"333333",x"333333",x"303030",x"313131",x"323232",x"343434",x"323232",x"313131",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"2f2f2f",x"333333",x"323232",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"2f2f2f",x"292929",x"313131",x"303030",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"432f21",x"432f21",x"452813",x"38200f",x"412411",x"412511",x"412411",x"3d220f",x"432712",x"3f2410",x"2b180b",x"3c210f",x"29180b",x"26160a",x"26160a",x"343434",x"343434",x"323232",x"323232",x"323232",x"5a5a5a",x"5f5f5f",x"575757",x"555555",x"636363",x"5b5b5b",x"666666",x"616161",x"5b5b5b",x"404040",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d220f",x"27160a",x"675345",x"43240f",x"24150a",x"26160a",x"3e2411",x"3a200f",x"3f2411",x"3d2411",x"3e2310",x"3f2411",x"3f2411",x"191008",x"3a210f",x"512f16",x"422612",x"3d2310",x"462913",x"412611",x"452813",x"422611",x"452914",x"462914",x"3f230f",x"402410",x"422611",x"412511",x"412611",x"402511",x"412511",x"402410",x"3a210e",x"3b210e",x"371f0d",x"331d0d",x"39200f",x"3a220f",x"311b0c",x"1f1208",x"371f0d",x"341d0c",x"301b0b",x"381f0d",x"2a180a",x"29170a",x"351e0d",x"321b0c",x"311b0b",x"201308",x"2f1a0b",x"361e0d",x"150e07",x"331c0c",x"301a0b",x"150e07",x"201208",x"2c170a",x"150e07",x"28170a",x"221409",x"1f1208",x"1c1108",x"2c180a",x"301b0b",x"211409",x"311c0c",x"25160a",x"25150a",x"1d1108",x"2e1a0b",x"301a0b",x"381f0e",x"3a200e",x"3c210f",x"371f0d",x"3b210f",x"391f0e",x"361d0d",x"381f0d",x"341c0c",x"2a170a",x"2f190b",x"311a0b",x"3a210f",x"150e07",x"150e07",x"000000",x"000000",x"22170f",x"22170f",x"281a0f",x"342012",x"331d0f",x"331e10",x"351e0f",x"351e0f",x"211409",x"3d220f",x"46372c",x"492c17",x"452a16",x"482b17",x"412512",x"3c2210",x"3f2412",x"432812",x"452813",x"412411",x"412411",x"432611",x"412511",x"3e2310",x"452813",x"422712",x"412612",x"432712",x"412511",x"452813",x"3f2511",x"432713",x"452813",x"422611",x"422712",x"462913",x"492c15",x"442813",x"3a200e",x"432612",x"412611",x"412511",x"3f2410",x"412511",x"3f2410",x"412410",x"3c210f",x"3c210f",x"3c210e",x"402410",x"402511",x"3b200e",x"361e0d",x"321c0c",x"40230f",x"341c0c",x"351d0d",x"371f0d",x"331c0c",x"3b210e",x"3c210e",x"331b0b",x"331c0b",x"381f0d",x"371e0d",x"391f0e",x"3b200e",x"351c0b",x"331b0b",x"351c0c",x"341c0b",x"361c0c",x"321c0c",x"3a200e",x"351d0c",x"3b200d",x"311b0b",x"371e0c",x"361e0d",x"3a200e",x"402410",x"3f230f",x"3e2310",x"3e220f",x"3b210e",x"3b210f",x"3c220f",x"39200e",x"3e220f",x"3e220f",x"3c210e",x"3e220e",x"3c210e",x"3d210e",x"3b200e",x"381e0c",x"3a1f0d",x"3e210f",x"472913",x"482914",x"492a14",x"482a14",x"452712",x"462812",x"492b14",x"492b15",x"442712",x"442813",x"492a14",x"462812",x"452813",x"472914",x"452813",x"472914",x"442813",x"412612",x"432611",x"412410",x"462712",x"432611",x"452813",x"432712",x"432611",x"422511",x"432712",x"412511",x"422612",x"452813",x"462913",x"432612",x"462813",x"432712",x"442712",x"402411",x"422612",x"402410",x"3d2311",x"422612",x"472a14",x"462914",x"351d0d",x"3e2411",x"402511",x"39210f",x"442712",x"432712",x"432711",x"422511",x"402310",x"3e220f",x"3e220f",x"402310",x"432712",x"412511",x"3f220f",x"3c210e",x"3c210f",x"3c210e",x"3a1f0d",x"3a200e",x"3a200e",x"402310",x"412510",x"3a200f",x"371e0e",x"3a200d",x"3b200e",x"3d210e",x"3d210f",x"3a200d",x"361d0c",x"381e0c",x"381e0c",x"371c0c",x"381e0d",x"3e210f",x"3a200e",x"3c210e",x"3a1f0d",x"3b200d",x"3e220e",x"3d210f",x"422510",x"402410",x"3e230f",x"432611",x"40230f",x"422510",x"4a2912",x"4a2912",x"000000",x"000000",x"000000",x"000000",x"381e0d",x"381e0d",x"492c18",x"2b1d14",x"433b32",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"23160b",x"332c24",x"332c24",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"525252",x"525252",x"383838",x"343434",x"484848",x"414141",x"4f4f4f",x"606060",x"656565",x"5e5e5e",x"3d3d3d",x"313131",x"333333",x"303030",x"3c3c3c",x"3f3f3f",x"424242",x"424242",x"464646",x"4a4a4a",x"474747",x"484848",x"434343",x"454545",x"4b4b4b",x"323232",x"313131",x"303030",x"323232",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"333333",x"323232",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"322f2e",x"333333",x"323232",x"323232",x"333333",x"313131",x"2f2f2f",x"2f2f2f",x"323232",x"323232",x"333333",x"323232",x"343434",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"363636",x"363636",x"323232",x"323232",x"333333",x"313131",x"333333",x"424242",x"404040",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"2f2f2f",x"292929",x"313131",x"303030",x"323232",x"2c2a28",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3f2b1d",x"3f2b1d",x"452813",x"422611",x"231409",x"3e2310",x"3f2410",x"3c210f",x"3a220f",x"180f07",x"351d0d",x"432611",x"29160a",x"241509",x"241509",x"4d4c4b",x"333333",x"313131",x"323232",x"333333",x"333333",x"333333",x"333333",x"333333",x"323232",x"2f2f30",x"333333",x"575452",x"333333",x"323232",x"333333",x"333333",x"333333",x"333333",x"323232",x"323232",x"333333",x"323232",x"333333",x"333333",x"333333",x"333333",x"343434",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"333333",x"323232",x"323232",x"303030",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"695547",x"695547",x"462712",x"2e1b0d",x"26160a",x"422713",x"2b180b",x"3d2310",x"3b2210",x"3b210f",x"412612",x"150e07",x"341d0d",x"3c220f",x"432510",x"381f0e",x"3b220f",x"422511",x"412511",x"3f2310",x"3f2310",x"422511",x"3f2410",x"432712",x"462813",x"3f2310",x"432611",x"3a210f",x"3d220f",x"3d220f",x"331c0c",x"3d220f",x"3d220f",x"3c210f",x"3d220f",x"3b210f",x"3c210f",x"3d230f",x"38200e",x"2d1a0b",x"38200e",x"3f2410",x"341d0d",x"3d230f",x"351d0d",x"381f0d",x"331d0c",x"2a170a",x"381f0e",x"381f0d",x"371e0d",x"381f0e",x"381f0e",x"351e0d",x"311b0b",x"311b0b",x"2a180a",x"2b180a",x"361e0d",x"2c190b",x"2f1a0b",x"2c180a",x"301b0b",x"2b180a",x"2b170a",x"301a0b",x"321c0c",x"3c220f",x"321c0c",x"3e220f",x"3a200e",x"3d230f",x"39200e",x"3a200e",x"3b210f",x"412511",x"3d2310",x"3d2310",x"39200f",x"361e0e",x"3d2410",x"3c2310",x"38210f",x"3c2210",x"150e07",x"150e07",x"000000",x"000000",x"20170f",x"20170f",x"27190f",x"2f1c10",x"352011",x"392313",x"361e0f",x"2f1b0d",x"221409",x"402410",x"47362a",x"452714",x"402613",x"432713",x"412613",x"3c2110",x"25150a",x"432511",x"432511",x"452712",x"402410",x"3d220f",x"391f0e",x"3d220f",x"3b200e",x"3a200e",x"3d220f",x"40230f",x"402410",x"412410",x"412410",x"452711",x"422511",x"462813",x"442712",x"432712",x"442712",x"432712",x"472913",x"432611",x"412410",x"442611",x"442611",x"412510",x"442611",x"482912",x"422511",x"4b2b14",x"472813",x"452812",x"442712",x"422511",x"3d220f",x"3f230f",x"442611",x"432511",x"3c220f",x"3f2310",x"442711",x"3c210f",x"3d220f",x"391f0d",x"3e220f",x"3d210e",x"3c200e",x"41240f",x"3d210e",x"3f230f",x"3f230f",x"432510",x"40230f",x"412510",x"40220e",x"40220f",x"40230f",x"472711",x"42240f",x"42240f",x"422510",x"452610",x"43240f",x"40220e",x"3f210e",x"42240f",x"472812",x"442511",x"472814",x"482914",x"412512",x"381e0d",x"3a210e",x"3c210f",x"3e2310",x"3b210f",x"402410",x"3e230f",x"361d0c",x"3b210e",x"402410",x"422612",x"41230f",x"41240f",x"41240f",x"3a200d",x"3f2310",x"3d220f",x"3e230f",x"422510",x"40230f",x"3e220f",x"3e220f",x"3d210f",x"3c200e",x"391e0d",x"3d210e",x"40230f",x"40230f",x"3d210e",x"3f230f",x"3d210f",x"3c220f",x"422510",x"412511",x"422611",x"412510",x"412510",x"412410",x"3e220f",x"3c210f",x"39200e",x"3a200e",x"3c210e",x"402310",x"402410",x"3e230f",x"3f2310",x"412410",x"40230f",x"41240f",x"432510",x"40230f",x"391f0d",x"442611",x"422511",x"3e230f",x"402411",x"442611",x"3a200f",x"371e0d",x"3e230f",x"432511",x"442712",x"452712",x"432611",x"412410",x"442611",x"432611",x"452711",x"472913",x"492a14",x"482915",x"472a15",x"4f2e18",x"482b17",x"482b17",x"3c2110",x"321b0b",x"321b0b",x"341c0c",x"3a210f",x"371f0e",x"3f2411",x"3c220f",x"412612",x"3a200e",x"3a200e",x"40230f",x"3f230f",x"40240f",x"422510",x"40230f",x"432611",x"3e220f",x"432611",x"412511",x"3e220f",x"432611",x"3e220f",x"472813",x"472813",x"000000",x"000000",x"000000",x"000000",x"341c0c",x"341c0c",x"4b2d19",x"271c12",x"3a3229",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"160e07",x"150e07",x"150e07",x"150e07",x"27160a",x"29190d",x"2f2821",x"2f2821",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595959",x"595959",x"595959",x"4a4a4a",x"343434",x"434343",x"4d4d4d",x"505050",x"5f5f5f",x"595959",x"333333",x"343434",x"323232",x"2c2c2c",x"313131",x"323232",x"323232",x"3a3a3a",x"3f3f3f",x"414141",x"3c3c3c",x"363636",x"3c3c3c",x"434343",x"434343",x"444444",x"313131",x"323232",x"333333",x"323232",x"313131",x"323232",x"555555",x"4e4e4e",x"515151",x"4b4b4b",x"393939",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"34302e",x"34302e",x"464646",x"626262",x"505050",x"464646",x"3c3c3c",x"3a3a3a",x"424242",x"3c3c3c",x"424242",x"414141",x"444444",x"444444",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e5e5e",x"5e5e5e",x"5b5b5b",x"535353",x"424242",x"414141",x"434343",x"4c4c4c",x"323232",x"313131",x"323232",x"2b2b2b",x"2d2d2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"323232",x"313131",x"313131",x"323232",x"2e2e2e",x"303030",x"292929",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"352519",x"352519",x"3f2410",x"412612",x"3a210f",x"412410",x"3d2310",x"422612",x"150e07",x"2e1a0b",x"3b210f",x"432611",x"27160a",x"29170a",x"29170a",x"4d4c4b",x"323232",x"323232",x"333333",x"323232",x"323232",x"313131",x"323232",x"333333",x"333333",x"323232",x"5e5d5c",x"61605f",x"504f4f",x"313131",x"323232",x"333333",x"333333",x"333333",x"323232",x"323232",x"333333",x"323232",x"333333",x"333333",x"333333",x"333333",x"343434",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"333333",x"323232",x"323232",x"303030",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"634d3e",x"634d3e",x"492b14",x"2d1a0c",x"221409",x"422713",x"341d0d",x"23150a",x"361e0d",x"3f2411",x"150e07",x"311c0d",x"38200f",x"3f2410",x"472812",x"3c220f",x"3e220f",x"432712",x"452813",x"412611",x"402511",x"402411",x"432611",x"3f230f",x"371e0e",x"3b200e",x"3a200e",x"371e0d",x"381f0d",x"371e0d",x"361d0c",x"331b0b",x"2b1508",x"321a0b",x"331c0b",x"361d0c",x"3a200e",x"371f0d",x"361e0d",x"351d0d",x"3b210f",x"3a200e",x"2d190b",x"321c0c",x"341d0d",x"381f0e",x"3a200e",x"3f2310",x"412510",x"412511",x"3d210f",x"412511",x"432611",x"412511",x"422611",x"351e0d",x"381f0d",x"371e0d",x"301b0c",x"351d0d",x"341c0c",x"351d0c",x"331c0c",x"311a0b",x"30190b",x"2f190b",x"321b0b",x"361d0c",x"361e0d",x"361d0c",x"381f0d",x"3a200e",x"3a200e",x"3a200e",x"391f0d",x"371f0e",x"3f2310",x"412511",x"3a210f",x"37200e",x"39200e",x"39200e",x"412410",x"3a210f",x"150e07",x"150e07",x"000000",x"000000",x"20160f",x"20160f",x"27190e",x"301d0f",x"351f11",x"392110",x"361e0f",x"341e0e",x"231509",x"402410",x"513e2f",x"472915",x"412612",x"402513",x"3f2412",x"392010",x"25150a",x"654630",x"6f4f37",x"75543b",x"77553a",x"735038",x"664731",x"6e4d35",x"77563d",x"74523a",x"7a563c",x"79553b",x"7d593d",x"805c41",x"815c41",x"7d593e",x"7c5a40",x"6d4c34",x"77553b",x"845f44",x"79573c",x"805d42",x"7a583e",x"6e4d35",x"75543b",x"6b4b33",x"6a4a32",x"765338",x"714e36",x"6c4a32",x"6e4c33",x"684730",x"715138",x"6f4c33",x"755138",x"74533a",x"7a563d",x"6d4c34",x"75543a",x"6d4c34",x"674831",x"593d29",x"493222",x"3d2a1c",x"3d220f",x"391f0d",x"3e220f",x"3d210e",x"3c200e",x"41240f",x"3d210e",x"3f230f",x"3f230f",x"432510",x"40230f",x"412510",x"40220e",x"40220f",x"40230f",x"472711",x"42240f",x"42240f",x"422510",x"452610",x"43240f",x"40220e",x"3f210e",x"42240f",x"472812",x"442511",x"472814",x"482914",x"482915",x"482915",x"3f2310",x"422611",x"442711",x"3e2310",x"422511",x"3f2310",x"3d220f",x"3c220f",x"3d230f",x"452812",x"1d1108",x"593c2b",x"6c4b34",x"725036",x"7a573b",x"704d35",x"77533a",x"6d4b35",x"77543a",x"6e4b33",x"62422d",x"684933",x"715138",x"7a573d",x"745139",x"7c593e",x"7d583f",x"7c593f",x"7e5a40",x"77543b",x"75533a",x"725138",x"7f5b40",x"79543b",x"7c593f",x"684831",x"77543b",x"735239",x"745239",x"715038",x"684831",x"7d5c41",x"6b4b35",x"684932",x"654832",x"644530",x"634530",x"573c28",x"362517",x"382618",x"40230f",x"391f0d",x"442611",x"422511",x"3e230f",x"402411",x"442611",x"3a200f",x"371e0d",x"3e230f",x"432511",x"442712",x"452712",x"432611",x"412410",x"442611",x"432611",x"452711",x"472913",x"492a14",x"482915",x"472a15",x"4f2e18",x"482b17",x"563d2d",x"412411",x"341c0d",x"321b0c",x"381e0d",x"381f0e",x"351d0d",x"3f2410",x"412511",x"402511",x"381f0e",x"3f230f",x"29170a",x"3f230f",x"40240f",x"422510",x"40230f",x"432611",x"3e220f",x"432611",x"412511",x"3e220f",x"432611",x"3e220f",x"472813",x"472813",x"000000",x"000000",x"000000",x"000000",x"341c0c",x"341c0c",x"4c2d17",x"2c1d14",x"3f372e",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"21140c",x"2d261e",x"2d261e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c4c4c",x"4c4c4c",x"4e4e4e",x"444444",x"353535",x"3f3f3f",x"404040",x"4c4c4c",x"5b5b5b",x"5b5b5b",x"333333",x"323232",x"323232",x"323232",x"343434",x"333333",x"323232",x"383838",x"373737",x"3d3d3d",x"3f3f3f",x"393939",x"373737",x"404040",x"404040",x"424242",x"464646",x"3f3f3f",x"333333",x"333333",x"323232",x"434343",x"3c3c3c",x"454545",x"4a4a4a",x"505050",x"434343",x"353535",x"323232",x"323232",x"333333",x"323232",x"000000",x"000000",x"4c4c4c",x"4c4c4c",x"505050",x"4b4b4a",x"4f4f4f",x"4c4c4c",x"535353",x"525252",x"4f4f4f",x"515151",x"505050",x"505050",x"5a5a5a",x"515151",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c2c2c",x"2a2a2a",x"333333",x"323232",x"444444",x"4c4c4c",x"4c4c4c",x"4b4b4b",x"505050",x"555555",x"616161",x"3e3e3e",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"323232",x"515151",x"333333",x"393939",x"313131",x"333333",x"292929",x"292929",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"271e16",x"271e16",x"422611",x"402511",x"38200e",x"2d1a0b",x"3f2511",x"442712",x"27160a",x"39200f",x"2f190a",x"3d220d",x"2c180a",x"29180b",x"29180b",x"474747",x"313131",x"414141",x"333333",x"313131",x"333333",x"333333",x"323232",x"313131",x"323232",x"313131",x"313131",x"323232",x"323232",x"323232",x"333333",x"323232",x"313131",x"323232",x"2e2e2e",x"333333",x"333333",x"313131",x"333333",x"323232",x"2f3030",x"313131",x"323232",x"323131",x"313131",x"343434",x"323232",x"313131",x"313131",x"303030",x"323232",x"343434",x"323232",x"323232",x"323232",x"313131",x"2e2e2e",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584133",x"584133",x"492b15",x"2a190c",x"2c1a0b",x"442813",x"371f0e",x"341f0e",x"39200e",x"3c220f",x"150e07",x"3a210f",x"38200f",x"402410",x"543117",x"452812",x"3f2410",x"3d230f",x"452812",x"432712",x"412511",x"402410",x"3f2410",x"3e230f",x"4b2a13",x"160f07",x"321c0c",x"2e1a0b",x"2f1a0b",x"2f190b",x"301a0b",x"2f1a0b",x"311b0b",x"2b1609",x"211106",x"2a1609",x"301b0b",x"321b0b",x"2e180a",x"311b0b",x"321b0c",x"2f190b",x"321b0b",x"2e190b",x"331c0c",x"351d0d",x"371f0d",x"371e0d",x"371f0d",x"331d0c",x"39200e",x"39200f",x"38200e",x"321c0c",x"331c0c",x"2f1a0b",x"331c0c",x"341d0d",x"341c0c",x"321b0b",x"341d0c",x"351d0d",x"311c0c",x"351e0d",x"371f0d",x"341c0c",x"321c0b",x"311b0b",x"3a200e",x"3b2210",x"38200f",x"3b210f",x"412411",x"3b200e",x"381f0d",x"391f0d",x"281509",x"241207",x"201006",x"200f06",x"2e180a",x"351c0c",x"361e0d",x"371f0d",x"150e07",x"150e07",x"000000",x"000000",x"1e140d",x"1e140d",x"26190e",x"2d1b0e",x"341f10",x"382010",x"341d0e",x"331c0c",x"24150a",x"432712",x"503c2f",x"472915",x"422714",x"3d2411",x"3f2412",x"3c220f",x"2f1a0b",x"77543b",x"805c41",x"886245",x"835d41",x"7e5940",x"78543a",x"7e5a40",x"866145",x"7f5b41",x"825b40",x"875f43",x"845d41",x"8e674a",x"896245",x"855e41",x"896347",x"735038",x"845d41",x"8b6446",x"866144",x"8d6648",x"835f42",x"795439",x"815b40",x"7f5a3f",x"7b563c",x"795438",x"7d5639",x"734f34",x"7d573c",x"785338",x"835c40",x"835c3f",x"7e593e",x"875e43",x"866043",x"7e593d",x"856043",x"7e583d",x"78543a",x"6c4a33",x"5a3f2b",x"453120",x"453120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b200e",x"150e07",x"150e07",x"150e07",x"564b41",x"564b41",x"584e44",x"3f2819",x"3f2819",x"150e07",x"150e07",x"150e07",x"492913",x"492913",x"3f2310",x"412511",x"412511",x"402410",x"3f230f",x"3c210e",x"402410",x"3d210e",x"3f2310",x"402410",x"201309",x"7c573d",x"896043",x"865d40",x"896145",x"865e42",x"8b6446",x"815a3f",x"8c6345",x"7d563b",x"7d573d",x"8c6447",x"64442f",x"7a583f",x"845d41",x"8c6547",x"876145",x"896448",x"8a6447",x"7e583d",x"7c583e",x"845d41",x"90684b",x"886043",x"886246",x"745036",x"865f44",x"845e42",x"775339",x"856043",x"795338",x"8b6549",x"845f42",x"755238",x"7b583e",x"755239",x"644530",x"63442d",x"3b2718",x"3c2819",x"3c2819",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412713",x"412713",x"442810",x"402610",x"402610",x"402610",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594233",x"594233",x"412511",x"361d0e",x"39200d",x"381e0d",x"3b200e",x"3b200e",x"3e2310",x"422612",x"412611",x"3b210f",x"432510",x"251509",x"251509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"000000",x"381f0d",x"381f0d",x"4f2d1a",x"2d1d13",x"3f362e",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"1f140a",x"2f261e",x"2f261e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"464646",x"464646",x"404040",x"3a3a3a",x"313131",x"363636",x"3d3d3d",x"444444",x"5b5b5b",x"636362",x"313131",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"353535",x"343434",x"3f3f3f",x"272728",x"535353",x"4c4c4c",x"404040",x"3c3c3c",x"414141",x"414141",x"434343",x"494949",x"4a4a4a",x"383838",x"373737",x"3f3f3f",x"3a3a3a",x"3c3c3c",x"3f3f3f",x"4b4b4b",x"4f4f4f",x"383838",x"313131",x"333333",x"343434",x"303030",x"313131",x"323333",x"505050",x"444444",x"43413f",x"403d3a",x"343333",x"333333",x"454545",x"434343",x"4b4b4b",x"505050",x"595959",x"434343",x"323232",x"323232",x"303030",x"333333",x"313131",x"333333",x"303030",x"323232",x"313131",x"303030",x"323232",x"2f2f2f",x"323232",x"313131",x"323232",x"303030",x"2d2d2d",x"2f2f2f",x"323232",x"323232",x"2a2a2a",x"2b2b2b",x"3b3b3b",x"545454",x"494949",x"525252",x"5b5b5b",x"636363",x"585858",x"464646",x"595958",x"484848",x"484848",x"303030",x"2e2e2e",x"353535",x"313131",x"313131",x"313131",x"323232",x"313131",x"292929",x"333333",x"424242",x"333333",x"4a4a4a",x"444444",x"4d4d4d",x"313131",x"313131",x"000000",x"323232",x"333333",x"333333",x"323232",x"323232",x"333333",x"333333",x"333333",x"323232",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"261d16",x"261d16",x"402511",x"3e2310",x"2a180b",x"2d1a0b",x"3a2210",x"3f2310",x"24150a",x"1f1208",x"2e1a0a",x"361d0b",x"29170a",x"27160a",x"27160a",x"323232",x"323232",x"2f2f2f",x"333333",x"313131",x"323232",x"313131",x"313131",x"333333",x"333333",x"323232",x"343434",x"323232",x"333333",x"303030",x"313131",x"313131",x"323232",x"333333",x"313131",x"323232",x"323232",x"313131",x"333333",x"343434",x"343434",x"313131",x"323232",x"323232",x"313131",x"333333",x"323232",x"343434",x"323232",x"353535",x"313131",x"313131",x"313131",x"323232",x"313131",x"2d2d2d",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543e31",x"543e31",x"4c2a14",x"24150a",x"2b190c",x"3f2512",x"2f1b0c",x"2f1c0d",x"3c2311",x"3f2411",x"150e07",x"2c190b",x"331d0e",x"3e220f",x"4f2f16",x"4a2b15",x"412511",x"3d2310",x"3f2411",x"422713",x"462814",x"432713",x"452813",x"4a2912",x"150e07",x"150e07",x"201309",x"2e1a0b",x"2f1a0b",x"2f190b",x"301a0b",x"2f1a0b",x"311b0b",x"2b1609",x"211106",x"2a1609",x"301b0b",x"321b0b",x"2e180a",x"311b0b",x"321b0c",x"2f190b",x"321b0b",x"2e190b",x"331c0c",x"351d0d",x"371f0d",x"371e0d",x"371f0d",x"331d0c",x"39200e",x"39200f",x"38200e",x"321c0c",x"331c0c",x"2f1a0b",x"331c0c",x"341d0d",x"341c0c",x"321b0b",x"341d0c",x"351d0d",x"311c0c",x"351e0d",x"371f0d",x"341c0c",x"321c0b",x"311b0b",x"3a200e",x"3b2210",x"38200f",x"341d0c",x"402510",x"221409",x"665343",x"1e1208",x"351d0d",x"3c220f",x"351e0d",x"3c2310",x"381f0d",x"3f2310",x"311a0b",x"3c210e",x"170f07",x"170f07",x"000000",x"000000",x"1e150d",x"1e150d",x"26180d",x"2f1c0f",x"321d0e",x"341d0e",x"371f0f",x"311b0c",x"26170b",x"412612",x"4f3b2d",x"492b15",x"412614",x"3e2310",x"3e2310",x"3f2310",x"25150a",x"805b3f",x"835e42",x"8c6649",x"875f43",x"855e42",x"8a6346",x"856044",x"825c41",x"8a6145",x"876043",x"876144",x"825a3e",x"866145",x"866044",x"8b6245",x"8b6344",x"896044",x"7d573a",x"906a4b",x"815a3e",x"896547",x"876043",x"8a6144",x"8d6649",x"845d41",x"815b3f",x"7c573d",x"7b5439",x"7e573b",x"7d573c",x"845e41",x"875f43",x"896042",x"805a3e",x"886043",x"896244",x"896143",x"845c41",x"7f5b3f",x"7a563c",x"79563c",x"563c29",x"442f20",x"442f20",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"241509",x"241509",x"150e07",x"150e07",x"150e07",x"564b41",x"564b41",x"584e44",x"3f2819",x"3f2819",x"150e07",x"150e07",x"150e07",x"150e07",x"422411",x"3c210e",x"402410",x"422611",x"402411",x"412510",x"3c210e",x"432611",x"3a200e",x"412410",x"412410",x"1c1108",x"815c41",x"8b6245",x"8d6345",x"855e42",x"896143",x"936a4b",x"865d40",x"8d6446",x"865e41",x"815b40",x"866044",x"8f6849",x"926a4b",x"8c6447",x"8c6547",x"8b6245",x"936a4d",x"8a6346",x"835c40",x"8b6446",x"896043",x"8f6748",x"8b6447",x"8c6547",x"845c40",x"845e43",x"7f5a3e",x"795338",x"986e4f",x"876144",x"90684c",x"91694b",x"7f593e",x"815c42",x"78543a",x"6f4c34",x"694831",x"402b1c",x"3f2b1c",x"3f2b1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422712",x"422712",x"4b2c12",x"422610",x"4d3b2d",x"4d3b2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"593c29",x"593c29",x"442713",x"361e0d",x"381e0d",x"381f0d",x"381f0e",x"381f0d",x"3a200e",x"412511",x"422612",x"3c220f",x"452611",x"28160a",x"28160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"39200e",x"39200e",x"462b18",x"2a1c11",x"3c332b",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"20130b",x"2d241c",x"2d241c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383838",x"383838",x"363636",x"343434",x"2d2d2d",x"343434",x"333333",x"313131",x"2e2e2e",x"545454",x"4f4f4f",x"424242",x"313131",x"343434",x"343434",x"333333",x"353535",x"323232",x"393939",x"3a3a3a",x"303030",x"3b3b3b",x"484848",x"414141",x"3c3c3c",x"3c3c3c",x"3c3c3c",x"3e3e3e",x"424242",x"444444",x"404040",x"3d3d3d",x"3f3f3f",x"3c3c3c",x"383838",x"3a3a3a",x"3f3f3f",x"404040",x"4b4b4b",x"4d4d4d",x"474747",x"333333",x"333333",x"313131",x"323333",x"333333",x"323232",x"343434",x"323232",x"323232",x"3a3a3a",x"363636",x"393939",x"434343",x"443d39",x"323232",x"323232",x"323232",x"313131",x"303030",x"333333",x"313131",x"333333",x"303030",x"323232",x"313131",x"303030",x"323232",x"2f2f2f",x"323232",x"313131",x"323232",x"303030",x"2d2d2d",x"323232",x"2f2f2f",x"323232",x"333333",x"4b4b4b",x"535353",x"3e3e3e",x"434343",x"3e3e3e",x"333333",x"3b3937",x"43403d",x"333333",x"303030",x"272828",x"292929",x"303030",x"2e2e2e",x"353535",x"313131",x"313131",x"2e2e2e",x"323232",x"333333",x"464646",x"4e4e4e",x"514e4c",x"545454",x"4b4b4b",x"535353",x"525252",x"303030",x"313131",x"333333",x"313131",x"323232",x"333333",x"333333",x"323232",x"333333",x"323232",x"323232",x"323232",x"303030",x"313131",x"313131",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2e2218",x"2e2218",x"3e230f",x"3b210f",x"3f2310",x"1a1008",x"38200e",x"351e0d",x"150e07",x"2b180a",x"1c1108",x"351d0c",x"261609",x"29170a",x"29170a",x"494949",x"3f3f3f",x"323232",x"2a2a2a",x"313131",x"313131",x"2f2f2f",x"333333",x"323232",x"383838",x"383838",x"3b3b3b",x"3e3e3e",x"333333",x"3a3a3a",x"383838",x"333333",x"313131",x"303030",x"2e2e2e",x"303030",x"313131",x"333333",x"323232",x"313131",x"333333",x"323232",x"303030",x"333333",x"333333",x"323232",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"383838",x"3b3b3b",x"363636",x"343434",x"353535",x"3e3b38",x"423e3a",x"252525",x"272727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543e30",x"543e30",x"4f2b14",x"2c190b",x"2d1a0c",x"402511",x"3f2411",x"150e07",x"3a2210",x"3e2411",x"150e07",x"38200f",x"24150a",x"3b200f",x"4f2f17",x"432713",x"402410",x"3c220f",x"361f0f",x"422713",x"402612",x"412612",x"402310",x"422511",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a210f",x"5c493b",x"5c493b",x"26160a",x"351d0d",x"381f0e",x"39200e",x"3a200f",x"371f0e",x"3b220f",x"2e190b",x"3a200d",x"180f08",x"180f08",x"000000",x"000000",x"1e140d",x"1e140d",x"25180d",x"2f1c0d",x"331d0e",x"382010",x"331d0e",x"2e1a0b",x"26160a",x"422713",x"483528",x"4a2b15",x"452813",x"462913",x"442712",x"3f230f",x"301b0c",x"846043",x"8d6548",x"956d4e",x"8d6345",x"956b4c",x"936b4d",x"956c4d",x"8c6547",x"92694b",x"875f43",x"8b6245",x"80593d",x"8f674b",x"886143",x"865e41",x"845c40",x"956b4b",x"876144",x"90684a",x"926a4c",x"936e4e",x"8d6446",x"8b6346",x"8e6447",x"875f43",x"7c563c",x"7d573b",x"8c6343",x"775237",x"875f43",x"875f42",x"896244",x"896043",x"845b3e",x"815a3d",x"8e6648",x"845c3f",x"906749",x"876143",x"7e583d",x"79583f",x"593f2b",x"442f20",x"442f20",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"371f0e",x"371f0e",x"150e07",x"150e07",x"150e07",x"574d43",x"574d43",x"544a3f",x"4d3221",x"4d3221",x"150e07",x"150e07",x"150e07",x"150e07",x"482812",x"3c210e",x"3c210f",x"3f2410",x"3b210f",x"402410",x"402410",x"3f240f",x"3b200e",x"412410",x"422510",x"211409",x"8c6649",x"855e41",x"8b6345",x"90694b",x"805b3f",x"78553c",x"8a5f43",x"936949",x"906647",x"926749",x"845c40",x"936a4b",x"936b4c",x"946a4b",x"91684a",x"956b4d",x"8c6347",x"875f43",x"865d41",x"92694a",x"8d6445",x"896044",x"966b4d",x"91684a",x"875f42",x"886043",x"855e40",x"906647",x"916849",x"91684a",x"956c4e",x"8f6749",x"815a3f",x"815c40",x"79543b",x"704e35",x"6b4a33",x"432e1e",x"442f1e",x"442f1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"36200f",x"36200f",x"37210c",x"271909",x"281909",x"281909",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583a26",x"583a26",x"422410",x"341c0c",x"371e0d",x"381f0d",x"3b210e",x"3a200e",x"3f2310",x"3d220f",x"492a14",x"412511",x"422510",x"211308",x"211308",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"2c190b",x"2c190b",x"3e230f",x"3e230f",x"4c2e1a",x"2a1b10",x"3b332b",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"2a170a",x"24170b",x"2d241a",x"2d241a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"333333",x"2e2e2e",x"323232",x"333333",x"2e2e2e",x"323232",x"323232",x"323232",x"313131",x"323232",x"333333",x"323232",x"333333",x"343434",x"333333",x"383838",x"383838",x"414141",x"393939",x"373737",x"383838",x"3b3b3b",x"3c3c3c",x"3d3d3d",x"3b3b3b",x"3e3e3e",x"3f3f3f",x"3d3d3d",x"404040",x"3c3c3c",x"3e3e3e",x"3b3b3b",x"3b3b3b",x"3f3f3f",x"404040",x"3f3f3f",x"464646",x"414141",x"505050",x"545454",x"404040",x"323232",x"323232",x"313131",x"4f4f4f",x"585858",x"525252",x"454545",x"404040",x"3a3a3a",x"3a3a3a",x"4a4543",x"4e4e4e",x"424242",x"3a3a3a",x"2d2e2e",x"2a2a2a",x"2e2e2e",x"2f2f2f",x"323232",x"2f2f2f",x"434343",x"4b4b4b",x"4f4f4f",x"505050",x"524e4b",x"5e5e5e",x"535353",x"2f2f2f",x"333333",x"333333",x"323232",x"3b3b3b",x"474747",x"3d3d3d",x"434343",x"3f3f3f",x"353535",x"3c3c3c",x"3b3b3b",x"474747",x"4f4f4f",x"4f4f4f",x"444444",x"414141",x"333333",x"333333",x"2f2f2f",x"323232",x"373737",x"303030",x"333333",x"3f3f3f",x"4d4d4d",x"505050",x"4a4a4a",x"454545",x"404040",x"3d3d3d",x"373737",x"3a3a3a",x"333333",x"333333",x"323232",x"333333",x"333333",x"383838",x"383838",x"313131",x"3e2d23",x"3a3a3a",x"363636",x"313131",x"343434",x"2f2f2f",x"313131",x"303030",x"313131",x"2c2c2c",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2e251d",x"2e251d",x"3b200e",x"3d220f",x"3d230f",x"150e07",x"3a200e",x"3a210f",x"150e07",x"381f0d",x"150e07",x"3a1f0d",x"271609",x"29170a",x"29170a",x"474747",x"505050",x"313131",x"343434",x"313131",x"2f2f2f",x"323232",x"333333",x"343434",x"313131",x"323232",x"2f2f2f",x"323232",x"303030",x"303030",x"323232",x"323232",x"333333",x"313131",x"313131",x"333333",x"333333",x"303030",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"3c3c3c",x"323232",x"323232",x"323232",x"343434",x"333333",x"343434",x"323232",x"323232",x"333333",x"2a2a2a",x"1e1e1e",x"2f2c2a",x"3e3b38",x"423e3a",x"252525",x"272727",x"272727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3729",x"4d3729",x"4a2913",x"2d1a0c",x"321d0e",x"3b2210",x"412511",x"150e07",x"3c2311",x"37200f",x"150e07",x"39200f",x"150e07",x"381f0e",x"513017",x"412612",x"3b210f",x"3c210f",x"432713",x"432814",x"3c2311",x"3e2411",x"3e2310",x"371f0e",x"150e07",x"150e07",x"4b4b4a",x"575757",x"515151",x"444444",x"4a4a4a",x"555555",x"4b4b4b",x"494949",x"444444",x"585858",x"404040",x"484745",x"4a4948",x"515050",x"4e4e4e",x"606060",x"545454",x"515151",x"515151",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"534033",x"534033",x"1f1208",x"3b200e",x"321c0c",x"3c210f",x"3a210f",x"3b200e",x"3f2410",x"341c0b",x"361e0d",x"150e07",x"150e07",x"000000",x"000000",x"1e140b",x"1e140b",x"24160b",x"2e1b0d",x"331d0e",x"381f10",x"331c0c",x"2f1a0b",x"25160a",x"442813",x"533b2b",x"4b2b15",x"472914",x"462913",x"442712",x"412410",x"29170a",x"8c6447",x"8c6648",x"956a4a",x"956b4c",x"987051",x"956d4e",x"946c4e",x"946a4c",x"8a6143",x"966d4d",x"95694a",x"7f5a3f",x"977050",x"916648",x"7a553b",x"91684a",x"916748",x"926748",x"967051",x"8c6649",x"936b4d",x"825b3b",x"835c3c",x"8a6042",x"8d6446",x"80593d",x"8b6244",x"8b6143",x"916648",x"8b6245",x"8b6244",x"906649",x"865d41",x"845c40",x"7e583c",x"896144",x"7c563b",x"865e41",x"886144",x"846043",x"79563d",x"5d422d",x"3c281a",x"3c281a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2410",x"3f2410",x"150e07",x"150e07",x"150e07",x"594f45",x"594f45",x"584e43",x"543c2d",x"543c2d",x"150e07",x"150e07",x"150e07",x"150e07",x"482912",x"432510",x"3f230f",x"3b200e",x"3f2310",x"3f2310",x"3c210f",x"412411",x"3a200d",x"40240f",x"3d220f",x"1c1108",x"8e6749",x"886145",x"92694a",x"966d4d",x"7d583c",x"926b4c",x"8d6344",x"9b6f4e",x"906647",x"946a4c",x"906546",x"906749",x"936a4b",x"936a4b",x"946b4d",x"91684a",x"875f43",x"90684a",x"8f6749",x"8f6647",x"8f6648",x"956949",x"9d7253",x"92694b",x"835c41",x"906648",x"8b6143",x"966c4d",x"a17957",x"845b3e",x"93694a",x"8b6140",x"8b6040",x"835c41",x"7b573d",x"735036",x"6c4b33",x"46301f",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38210e",x"38210e",x"2d1c09",x"271809",x"261809",x"261809",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543623",x"543623",x"3c210e",x"341c0c",x"3a200e",x"3d220f",x"3c220f",x"391f0e",x"3d220f",x"3e220f",x"492b14",x"412511",x"42240f",x"221409",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"170f07",x"170f07",x"432611",x"432611",x"391f0d",x"391f0d",x"502f1b",x"311e12",x"342d25",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"27180b",x"2b2117",x"2b2117",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b3b3b",x"373737",x"303030",x"2f2f2f",x"333333",x"333333",x"2e2e2e",x"323232",x"323232",x"323232",x"333333",x"333333",x"333333",x"313131",x"313131",x"323232",x"323232",x"363636",x"393939",x"3a3a3a",x"3a3a3a",x"3c3c3c",x"3b3b3b",x"393939",x"3a3a3a",x"3b3b3b",x"3d3d3d",x"3c3c3c",x"3c3c3c",x"3f3f3f",x"383838",x"3f3f3f",x"3a3a3a",x"393939",x"3c3c3c",x"3b3b3b",x"3e3e3e",x"3e3e3e",x"404040",x"404040",x"414141",x"434343",x"3c3735",x"464646",x"474747",x"4b4b4b",x"484848",x"434343",x"383838",x"3f3f3f",x"3f3f3f",x"3f3f3f",x"3e3e3e",x"3b3b3b",x"464646",x"424242",x"464646",x"464646",x"3f3f3f",x"333333",x"414141",x"454545",x"444444",x"3e3937",x"444444",x"494949",x"434343",x"484949",x"444444",x"484848",x"494949",x"494949",x"4e4e4e",x"4d4d4d",x"3e3e3e",x"404040",x"313131",x"313131",x"323232",x"474747",x"3d3d3d",x"3d3d3d",x"434343",x"434343",x"434343",x"3e3e3e",x"434343",x"474747",x"474747",x"4a4a4a",x"3e3e3e",x"424242",x"464646",x"474848",x"3b3b3b",x"464646",x"414141",x"3c3c3c",x"383838",x"3f3f3f",x"333333",x"3d3d3d",x"383838",x"3f3f3f",x"434343",x"4f4f4f",x"444444",x"414141",x"373737",x"313131",x"383838",x"3f3f3f",x"454545",x"353535",x"353535",x"323232",x"323232",x"333333",x"3f3f3f",x"464646",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2c2016",x"2c2016",x"361d0c",x"3c210f",x"3e2310",x"432612",x"3b2210",x"37200f",x"361e0d",x"3a200d",x"150e07",x"3c210d",x"261609",x"2a180b",x"2a180b",x"525252",x"555555",x"323232",x"313131",x"323232",x"323232",x"323232",x"313131",x"323232",x"313131",x"303030",x"303030",x"303030",x"2e2e2e",x"313131",x"313131",x"333333",x"313131",x"333333",x"343434",x"323232",x"333333",x"333331",x"333333",x"333333",x"323232",x"333333",x"333232",x"333333",x"3d3d3d",x"323232",x"323232",x"303030",x"323232",x"323232",x"343434",x"343434",x"292116",x"323232",x"2c2c2c",x"3b3b3a",x"3c3937",x"342f29",x"3b3632",x"303030",x"2f2f2f",x"2f2f2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3426",x"4a3426",x"4d2c13",x"301c0d",x"2b1a0c",x"37200f",x"422612",x"432713",x"3d2311",x"3b210f",x"3a220f",x"3a210f",x"150e07",x"381f0e",x"492b13",x"3f2411",x"3b210e",x"381f0d",x"39200f",x"432814",x"3d2411",x"3b2310",x"3c2210",x"3a210f",x"150e07",x"4b4b4a",x"4b4b4a",x"595959",x"515151",x"383838",x"4a4a4a",x"636363",x"4b4b4b",x"494949",x"444444",x"585858",x"404040",x"484745",x"4a4948",x"515050",x"4e4e4e",x"606060",x"545454",x"515151",x"515151",x"515151",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"553f30",x"553f30",x"28170a",x"3c210f",x"381f0e",x"39200e",x"3b210f",x"3a210f",x"341d0d",x"2f1a0b",x"371e0d",x"150e07",x"150e07",x"000000",x"000000",x"1d130b",x"1d130b",x"25160c",x"2d1a0d",x"331d0e",x"341d0d",x"341d0c",x"311b0c",x"26160a",x"3f2410",x"4c3628",x"492a13",x"432712",x"432712",x"402410",x"412511",x"27160a",x"8a6346",x"8b6346",x"956c4c",x"92694b",x"936c4e",x"90684a",x"956a4c",x"906748",x"8a6145",x"93694a",x"92694a",x"835b3e",x"966e4e",x"926748",x"835a3e",x"91684a",x"896144",x"a07352",x"997353",x"8c6647",x"865f42",x"875d3e",x"885e40",x"845c3c",x"8f6647",x"91694a",x"956949",x"906647",x"93694a",x"8a6042",x"8d6445",x"91674a",x"8a6042",x"8c6344",x"865e40",x"93684a",x"845d40",x"845e41",x"79553b",x"896247",x"79573d",x"5a3f2d",x"483323",x"483323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"544a40",x"544a40",x"5d5248",x"4e3221",x"4e3221",x"150e07",x"150e07",x"150e07",x"150e07",x"4d2b14",x"3e220f",x"422510",x"3d210e",x"3c220f",x"3d230f",x"3d220f",x"3d220f",x"371e0d",x"381e0d",x"3c210e",x"201309",x"855d41",x"835c41",x"956b4e",x"986e4f",x"93684a",x"906848",x"895f40",x"8f6545",x"976d4d",x"93694b",x"946a4a",x"946a4c",x"866043",x"9b7151",x"997051",x"956c4d",x"90674a",x"946e4f",x"875f43",x"936a4a",x"8d6446",x"8d6346",x"976d4e",x"93684b",x"90674a",x"926849",x"916648",x"996d4d",x"9f7c59",x"996e4f",x"926647",x"89603f",x"8a5f41",x"8a6141",x"865e42",x"79553b",x"735137",x"473120",x"46311f",x"46311f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a220f",x"3a220f",x"2f1e0a",x"291a09",x"291a09",x"291a09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563c2b",x"563c2b",x"3b200e",x"321b0b",x"351d0d",x"3d2310",x"3e2310",x"381e0d",x"432712",x"3b200e",x"462913",x"402511",x"41240f",x"28160a",x"28160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"19110a",x"19110a",x"311c0c",x"311c0c",x"341c0b",x"341c0b",x"52321c",x"2c1c11",x"372f28",x"150e07",x"150e07",x"150e07",x"150e07",x"201308",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"301e0c",x"251c13",x"251c13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"373737",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"333333",x"333333",x"555555",x"323232",x"383838",x"363636",x"383838",x"363636",x"3a3a3a",x"373737",x"383838",x"3b3b3b",x"343434",x"3b3b3b",x"3e3e3e",x"3d3d3d",x"3b3b3b",x"3b3b3b",x"363636",x"393939",x"3b3b3b",x"3e3e3e",x"373737",x"3c3c3c",x"3c3c3c",x"404040",x"3f3f3f",x"404040",x"434343",x"464646",x"454443",x"414141",x"454545",x"454545",x"414141",x"414141",x"414141",x"3b3b3b",x"3e3e3e",x"3d3d3d",x"434343",x"454545",x"434343",x"434343",x"434343",x"3a3b3b",x"323232",x"3b3b3b",x"313131",x"3f3f3f",x"404040",x"434343",x"434343",x"404040",x"383838",x"444444",x"424242",x"454545",x"3e3e3e",x"414141",x"3d3d3d",x"3e3e3e",x"404040",x"313131",x"323232",x"323232",x"434343",x"3d3d3d",x"3c3c3c",x"3d3d3d",x"3c3d3d",x"383838",x"404040",x"414141",x"414141",x"434343",x"383838",x"3d3d3d",x"404040",x"3b3b3b",x"414242",x"404040",x"424242",x"404040",x"373737",x"414141",x"323232",x"3f3f3f",x"323232",x"3d3d3d",x"3f3f3f",x"464646",x"444444",x"3d3d3d",x"3d3d3d",x"3e3e3e",x"444444",x"4a4a4a",x"4d4d4d",x"4d4d4d",x"494949",x"4c4c4c",x"444444",x"4b4b4b",x"454545",x"424242",x"494949",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"241c15",x"241c15",x"351d0c",x"3b210f",x"3b200e",x"3d2310",x"37200f",x"38200f",x"321b0b",x"381f0d",x"150e07",x"381f0d",x"221408",x"2a180b",x"2a180b",x"666666",x"626262",x"5e5e5e",x"4b4b4b",x"4c4c4c",x"323232",x"303030",x"323232",x"313131",x"313131",x"313131",x"303030",x"2d2d2d",x"333333",x"2d2d2d",x"333333",x"313131",x"313131",x"343434",x"323232",x"323232",x"323232",x"353535",x"313131",x"313131",x"292929",x"313131",x"333333",x"333333",x"323232",x"343434",x"313131",x"343434",x"333333",x"323232",x"363636",x"343434",x"333333",x"313131",x"303030",x"303030",x"37322d",x"3e3a37",x"3d3a37",x"292929",x"2a2a2a",x"2a2a2a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3426",x"4a3426",x"472812",x"2a190b",x"23150a",x"3d2411",x"442813",x"3e2511",x"361f0e",x"351d0d",x"26160a",x"39210f",x"150e07",x"371e0d",x"4b2b14",x"412511",x"3b210e",x"351d0c",x"3f2410",x"462914",x"432713",x"3e2311",x"3f2411",x"39210f",x"150e07",x"323232",x"323232",x"333333",x"323232",x"333333",x"313030",x"5f5a57",x"534d47",x"353535",x"333333",x"323232",x"333333",x"343332",x"343332",x"313131",x"343434",x"323232",x"313131",x"48433e",x"4b4742",x"565656",x"333333",x"353535",x"323232",x"313131",x"333333",x"333333",x"313131",x"313131",x"313131",x"343434",x"333333",x"333333",x"343434",x"323232",x"434343",x"323232",x"333333",x"333333",x"333333",x"343434",x"343434",x"323130",x"323232",x"343333",x"343333",x"000000",x"000000",x"533e31",x"533e31",x"27170a",x"3d220f",x"3a200e",x"381f0e",x"3b210e",x"3a210f",x"341c0c",x"361e0d",x"391f0e",x"150e07",x"150e07",x"000000",x"000000",x"1d130a",x"1d130a",x"25170b",x"2d1b0d",x"331d0e",x"311b0c",x"341d0c",x"321c0c",x"26160a",x"3d210e",x"473326",x"492914",x"432814",x"432712",x"412511",x"3d220f",x"321c0d",x"875f42",x"906647",x"926748",x"946a4c",x"997051",x"916749",x"976d4d",x"936949",x"8f6547",x"8d6446",x"8d6548",x"896044",x"986e4f",x"916748",x"8c6243",x"956b4c",x"865d41",x"966e4e",x"927050",x"976b4d",x"8f6749",x"8d6547",x"8b6242",x"8b6141",x"8f6343",x"8c6244",x"966b4d",x"8e6546",x"8f6447",x"885f41",x"926647",x"91684a",x"896042",x"92694a",x"8c6243",x"926849",x"906648",x"8b6345",x"865f43",x"856146",x"7b593d",x"5e4330",x"4b3525",x"4b3525",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"594e44",x"594e44",x"594d43",x"4a2d1a",x"4a2d1a",x"150e07",x"150e07",x"150e07",x"150e07",x"512e15",x"3f2310",x"3f2310",x"3c210e",x"3b200e",x"3e230f",x"402410",x"472913",x"351d0c",x"371e0d",x"3b200d",x"1f1208",x"886144",x"8d6446",x"956d4d",x"8d6547",x"906748",x"936e50",x"8a6142",x"8b6345",x"95694a",x"926849",x"936648",x"9c7250",x"936a4b",x"996f51",x"997151",x"966c4d",x"956a4a",x"90674a",x"8a6143",x"956a4b",x"896143",x"8e6547",x"966c4e",x"926748",x"976c4e",x"9a6e4f",x"956a4a",x"a37656",x"956c4c",x"9b7454",x"966b4d",x"976b4b",x"8f6443",x"885f40",x"7f593a",x"785338",x"74543a",x"473120",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a2210",x"3a2210",x"2d1d0a",x"291a09",x"291a09",x"291a09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"573d2c",x"573d2c",x"3d220f",x"361e0d",x"371e0d",x"432712",x"3e2310",x"3a200e",x"3f2410",x"3d2310",x"492b14",x"3f2410",x"40230f",x"241509",x"241509",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"351d0c",x"351d0c",x"51321e",x"2c1c10",x"393129",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"21150b",x"261d15",x"261d15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d2d2d",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"313131",x"303030",x"323232",x"323232",x"313131",x"333333",x"333333",x"333333",x"323232",x"373737",x"383838",x"363636",x"363636",x"383838",x"373737",x"383838",x"383838",x"3a3a3a",x"3d3d3d",x"393a3a",x"3d3d3d",x"3c3c3c",x"373737",x"373737",x"3d3d3d",x"383838",x"3c3c3c",x"383838",x"3d3d3d",x"3e3e3e",x"414141",x"444444",x"424242",x"484848",x"474747",x"4a4a4a",x"474747",x"4d4d4d",x"464646",x"434343",x"434343",x"3e3e3e",x"3a3a3a",x"3e3e3e",x"3e3e3e",x"3d3d3d",x"404040",x"404040",x"414141",x"444444",x"3d3d3d",x"3f3f3f",x"3d3d3d",x"404040",x"464646",x"414141",x"434343",x"454545",x"444240",x"424242",x"434343",x"474747",x"4a4a4a",x"484848",x"4e4e4e",x"474747",x"424242",x"444444",x"303030",x"343434",x"313131",x"4b4b4b",x"3b3b3b",x"3f3f3f",x"373737",x"414141",x"404040",x"454545",x"434343",x"484848",x"474747",x"414141",x"414141",x"404040",x"474747",x"474747",x"4e4e4e",x"454545",x"3c3c3c",x"3d3d3d",x"3d3d3d",x"3d3e3e",x"4e4e4e",x"313131",x"393939",x"3e3e3e",x"494949",x"535353",x"505151",x"494949",x"474747",x"484847",x"4d4d4d",x"565656",x"4d4d4d",x"4f4f4f",x"505050",x"4e4e4e",x"454545",x"4b4b4b",x"4f4f4f",x"515151",x"4c4c4c",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"322217",x"322217",x"3b200e",x"321c0d",x"3b210e",x"150e07",x"38200f",x"3a200f",x"241509",x"301a0b",x"251509",x"3b200d",x"29180b",x"26160a",x"26160a",x"5d5d5c",x"666666",x"645b53",x"5e5e5e",x"5d5d5d",x"323232",x"323232",x"313232",x"333333",x"303030",x"313131",x"2e2e2e",x"2e2e2e",x"323232",x"2e2e2e",x"2e2e2e",x"323232",x"343434",x"323232",x"313131",x"303030",x"313131",x"333333",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"4a4a4a",x"323232",x"333333",x"333333",x"333333",x"333333",x"333333",x"333333",x"323232",x"323232",x"323232",x"545454",x"3b3b3b",x"414140",x"404040",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c372b",x"4c372b",x"4d2c15",x"2f1c0d",x"2b1a0c",x"3b2210",x"442813",x"150e07",x"36200f",x"3b220f",x"150e07",x"39210f",x"1d1108",x"39200e",x"4b2a14",x"402411",x"3c210f",x"321b0c",x"412511",x"3f2310",x"3c2310",x"3a210f",x"402411",x"3c2311",x"150e07",x"343231",x"343231",x"323232",x"343434",x"333232",x"343333",x"5c5753",x"3b3937",x"323232",x"323232",x"333333",x"333333",x"353433",x"343331",x"353434",x"333232",x"323232",x"323131",x"49453f",x"323232",x"565656",x"333333",x"353535",x"323232",x"313131",x"333333",x"333333",x"313131",x"313131",x"313131",x"343434",x"333333",x"333333",x"343434",x"323232",x"434343",x"323232",x"333333",x"333333",x"333333",x"343434",x"343434",x"323130",x"323232",x"343333",x"343333",x"000000",x"000000",x"4f3828",x"4f3828",x"2b190b",x"3f2310",x"351d0d",x"351d0d",x"3b200e",x"3e2310",x"381f0e",x"371f0e",x"3b210f",x"150e07",x"150e07",x"000000",x"000000",x"1d130b",x"1d130b",x"24170c",x"2e1c0d",x"321c0c",x"321c0c",x"331c0b",x"341d0d",x"25150a",x"3e2410",x"4b3425",x"462813",x"492b16",x"412612",x"422613",x"3c210f",x"27160a",x"80593f",x"8f6547",x"8d6648",x"91684b",x"a07655",x"9b7151",x"9b7050",x"9c7050",x"90674a",x"91684a",x"906647",x"875f42",x"986f50",x"8b6447",x"845d41",x"876044",x"8a6143",x"966c4d",x"957050",x"986f4f",x"90674a",x"8d6447",x"946a4c",x"906543",x"8d6343",x"8a6143",x"966c4c",x"94694a",x"8c6143",x"875d3f",x"936749",x"8e6447",x"8b6143",x"986d4c",x"8b6143",x"8c6245",x"845d40",x"8b6346",x"91694b",x"8d6649",x"73533a",x"59402e",x"4d3727",x"4d3727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"574d43",x"574d43",x"554a41",x"4f3320",x"4f3320",x"3a200e",x"150e07",x"150e07",x"150e07",x"4b2913",x"432711",x"3e220f",x"3c210e",x"331b0b",x"432611",x"3e220f",x"432712",x"3a1f0d",x"341c0c",x"3d210e",x"1b1008",x"825b40",x"936a4b",x"986d4e",x"866043",x"956b4b",x"8e6649",x"875d40",x"8f6446",x"825a3d",x"966a4b",x"8d6344",x"876144",x"966b4c",x"78543c",x"986f50",x"956d4e",x"946b4c",x"7a553d",x"8d6446",x"906546",x"815b40",x"886044",x"8f6649",x"8a6144",x"91684a",x"9a6f4e",x"986c4c",x"a27654",x"956b4b",x"a07655",x"9d7151",x"8f6545",x"93694b",x"8a5f3f",x"865d3f",x"775137",x"714f37",x"463120",x"463120",x"463120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"36200e",x"36200e",x"271909",x"271909",x"281909",x"281909",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543623",x"543623",x"422410",x"371e0d",x"371e0d",x"3e2310",x"3b210f",x"3b210f",x"432611",x"432712",x"412612",x"412510",x"42240f",x"2f1b0c",x"2f1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"1d1209",x"1d1108",x"351c0c",x"351c0c",x"503624",x"2c1b10",x"383028",x"150e07",x"150e07",x"150e07",x"150e07",x"26150a",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"25160b",x"2b1f16",x"2b1f16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d2d2d",x"2d2d2d",x"323232",x"313131",x"323232",x"333333",x"333333",x"323232",x"323232",x"313131",x"303030",x"303030",x"313131",x"333333",x"323232",x"343434",x"383838",x"343434",x"373737",x"353535",x"353535",x"323232",x"3d3d3d",x"3b3b3b",x"383838",x"393939",x"3e3e3e",x"3f3f3f",x"404040",x"3f3f3f",x"3c3c3c",x"3a3a3a",x"3c3c3c",x"3d3d3d",x"353535",x"3b3b3b",x"3b3b3b",x"3c3c3c",x"3f3f3f",x"414141",x"4c4c4c",x"535353",x"5f5f5f",x"606060",x"5f5f5f",x"5c5854",x"67625e",x"5c5956",x"585858",x"4d4d4d",x"414141",x"393939",x"373737",x"373737",x"424242",x"454545",x"494949",x"555555",x"4c4c4c",x"535353",x"5c5c5c",x"4e4e4e",x"545454",x"565656",x"5b5b5b",x"5b5b5b",x"585858",x"5d5d5d",x"5f5f5f",x"5f5f5f",x"595959",x"575757",x"605b57",x"615c57",x"5f5a54",x"484848",x"4f4f4f",x"484848",x"464646",x"4f4f4f",x"3b3b3b",x"3a3a3a",x"3b3b3b",x"4b4b4b",x"515151",x"474747",x"535353",x"575757",x"64605c",x"67615c",x"64605b",x"66615d",x"64605b",x"625d59",x"645e5a",x"5e5a56",x"5a5a5a",x"4b4b4b",x"3c3c3c",x"383838",x"383838",x"383838",x"353535",x"323232",x"333333",x"3e3e3e",x"635d57",x"5b5550",x"51504e",x"494949",x"4b4b4b",x"4a4a4a",x"4c4c4c",x"454545",x"4d4d4d",x"4c4c4c",x"454545",x"4e4e4e",x"525251",x"504f4f",x"4e4e4e",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"342419",x"342419",x"381e0d",x"3d2210",x"301b0c",x"301c0d",x"3b210f",x"3d2411",x"201308",x"261609",x"2f1a0b",x"3b200d",x"2c190c",x"29180b",x"29180b",x"535352",x"7a756f",x"746e67",x"76706b",x"4b4b4b",x"454545",x"323232",x"313232",x"333333",x"303030",x"313131",x"2e2e2e",x"2e2e2e",x"323232",x"2e2e2e",x"2e2e2e",x"323232",x"343434",x"323232",x"313131",x"303030",x"313131",x"333333",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"4a4a4a",x"323232",x"333333",x"333333",x"333333",x"333333",x"333333",x"333333",x"323232",x"323232",x"323232",x"545454",x"3b3b3b",x"414140",x"404040",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3528",x"4a3528",x"4b2c15",x"2c1a0c",x"27170b",x"3d2411",x"3c2311",x"341f0e",x"3c2311",x"3a210f",x"180f07",x"26160a",x"321c0d",x"3c220f",x"4d2b13",x"3e2310",x"3a210f",x"351d0c",x"3f2411",x"3c2210",x"3c230f",x"3d2210",x"432713",x"452914",x"150e07",x"555555",x"5b5b5b",x"616161",x"333333",x"333232",x"373736",x"595653",x"3b3937",x"323232",x"323232",x"333333",x"333333",x"353433",x"5a5a5a",x"4b4b4b",x"4a4a4a",x"313131",x"343434",x"454545",x"454545",x"313131",x"333333",x"313131",x"2a2b2b",x"323232",x"313131",x"333333",x"313131",x"313131",x"343434",x"2f2f2f",x"313131",x"323232",x"343434",x"323232",x"434343",x"323232",x"313131",x"323232",x"313131",x"323232",x"303030",x"333333",x"313131",x"333333",x"333333",x"000000",x"000000",x"4a3425",x"4a3425",x"1e1208",x"341d0d",x"341d0d",x"311b0c",x"311b0b",x"38200e",x"3c2210",x"3b210e",x"361e0d",x"150e07",x"150e07",x"000000",x"000000",x"1c120a",x"1c120a",x"231509",x"2e1a0b",x"311c0c",x"311b0b",x"311b0b",x"331c0c",x"25150a",x"3d220f",x"4a3527",x"472913",x"422714",x"432813",x"432712",x"3e2311",x"311c0d",x"7e583b",x"8c6547",x"8d6548",x"9b714f",x"a07553",x"9e7352",x"9a7051",x"966e4e",x"956b4c",x"946e4e",x"956a4a",x"8e6445",x"a07654",x"946b4c",x"8e6547",x"7b563d",x"8e6547",x"9b7152",x"9a7150",x"9b7150",x"8a6143",x"8c6345",x"8f6445",x"865d42",x"8d6547",x"845b3e",x"986e4e",x"8c6243",x"8e6446",x"8c6143",x"946849",x"8c6244",x"986d4b",x"956b4b",x"8d6344",x"8d6345",x"815b40",x"8c6244",x"876145",x"7c5a3f",x"77543b",x"5c432f",x"4e3928",x"4e3928",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"554b41",x"554b41",x"473c32",x"523624",x"523624",x"39200e",x"150e07",x"150e07",x"150e07",x"432510",x"412511",x"3d220f",x"3e220f",x"361c0c",x"3d2210",x"3d220f",x"3f2411",x"39200d",x"3b200e",x"3d220f",x"201309",x"6f4c35",x"93694a",x"966c4b",x"926748",x"8d6546",x"866247",x"855c3f",x"865e42",x"865c40",x"976c4d",x"956a4b",x"9f7554",x"9a6f4f",x"986e4e",x"866045",x"936a4c",x"8a6447",x"825c42",x"815c41",x"7c573e",x"865e41",x"835d41",x"93694b",x"926949",x"94694a",x"9f7252",x"9c7050",x"9b6f4f",x"976d4e",x"a27655",x"976c4c",x"8a6144",x"896043",x"885f43",x"865f42",x"79543a",x"715139",x"45301f",x"463120",x"463120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200e",x"38200e",x"2f1e0a",x"2a1b09",x"221608",x"221608",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563723",x"563723",x"3f230f",x"39200e",x"371d0c",x"3e2310",x"3c220f",x"381f0d",x"422612",x"402411",x"412612",x"412511",x"40220e",x"28170a",x"28170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"201309",x"381e0d",x"381e0d",x"5c402e",x"261910",x"3a322a",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"150e07",x"150e07",x"150e07",x"191008",x"2d1a0b",x"2a190c",x"271d16",x"271d16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"313131",x"313131",x"323232",x"323232",x"313131",x"303030",x"313131",x"2f2f2f",x"333333",x"313131",x"323232",x"333333",x"323232",x"333333",x"353535",x"393939",x"393939",x"393939",x"343434",x"484848",x"3a3a3a",x"474747",x"3c3c3c",x"3d3d3d",x"3f3f3f",x"444444",x"424242",x"424242",x"3f3f3f",x"3e3e3e",x"3b3b3b",x"383838",x"3a3a3a",x"393939",x"393939",x"3e3e3e",x"404040",x"535353",x"616161",x"464645",x"403f3e",x"454341",x"53504c",x"5c5854",x"6a645e",x"67615b",x"514f4c",x"434343",x"313131",x"3b3b3b",x"313131",x"333333",x"333333",x"323232",x"323232",x"313131",x"615b54",x"655f59",x"665f57",x"645d57",x"66605a",x"655f59",x"655f5a",x"6c645e",x"66615c",x"66605c",x"69645f",x"645e59",x"605a55",x"635d57",x"615b55",x"655f59",x"545351",x"525252",x"4c4c4c",x"454545",x"4b4b4b",x"313131",x"373737",x"333333",x"303030",x"323232",x"323232",x"333333",x"353535",x"333333",x"665e57",x"67615c",x"64605b",x"66615d",x"64605b",x"625d59",x"645e5a",x"555250",x"494949",x"464646",x"5e5e5e",x"484949",x"393939",x"383838",x"3e3e3e",x"3e3e3e",x"3c3c3c",x"333333",x"333333",x"5b5550",x"464545",x"3b3b3b",x"3d3c3c",x"454545",x"565656",x"5a5a5a",x"545454",x"363636",x"383735",x"575350",x"5c5854",x"54524f",x"4d4d4d",x"4e4e4e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2d231b",x"2d231b",x"371d0c",x"3b210f",x"391f0e",x"37200f",x"361e0d",x"3e2310",x"2c1a0c",x"361e0c",x"3a200e",x"402410",x"28180b",x"25150a",x"666666",x"60605f",x"6e6761",x"716b65",x"5b534b",x"454545",x"5b5b5b",x"676665",x"676766",x"6b6966",x"676665",x"666564",x"636261",x"696766",x"696867",x"646463",x"696969",x"616161",x"5e5e5e",x"605f5f",x"5b5a5a",x"585757",x"4a4a4a",x"525252",x"5d5d5d",x"6a6a68",x"686867",x"5b5b5b",x"4a4a4a",x"4f4f4f",x"5b5b5b",x"5d5d5d",x"5d5d5d",x"545454",x"5e5e5e",x"575656",x"585756",x"5e5c5b",x"585654",x"535252",x"454545",x"363636",x"303030",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463225",x"463225",x"4d2d15",x"221409",x"25160a",x"402612",x"412712",x"341d0d",x"3d2311",x"3d230f",x"1e1208",x"2f1b0c",x"351d0d",x"432711",x"573116",x"3f2411",x"3c210f",x"281307",x"3f2411",x"3b2210",x"3a200f",x"3b210f",x"3f2511",x"502f17",x"323232",x"414040",x"4f4f4f",x"5c5c5c",x"666565",x"323232",x"2d2d2d",x"313131",x"535353",x"3b3b3b",x"383838",x"5a5a5a",x"474747",x"383838",x"5a5a5a",x"4b4b4b",x"4a4a4a",x"343434",x"313131",x"323232",x"323232",x"363636",x"2e2e2e",x"313131",x"303030",x"343434",x"323232",x"2f2f2f",x"313131",x"303030",x"333333",x"313131",x"313131",x"313131",x"313131",x"323232",x"333231",x"303030",x"333333",x"333333",x"313131",x"333333",x"333333",x"323232",x"323232",x"323232",x"323232",x"000000",x"000000",x"513a2a",x"513a2a",x"211309",x"3b210e",x"39200f",x"3a200e",x"371f0e",x"341d0d",x"37200f",x"38200e",x"3a200e",x"150e07",x"150e07",x"000000",x"000000",x"1a1008",x"1a1008",x"231409",x"2d1a0b",x"311c0c",x"341c0c",x"321b0b",x"331c0c",x"25150a",x"391f0d",x"4b3426",x"432512",x"412712",x"432714",x"3e2311",x"3c2210",x"29170b",x"6d4932",x"91694a",x"966c4e",x"966d4f",x"9d7454",x"9b7151",x"92694a",x"9b7151",x"95694a",x"986e4e",x"936849",x"906647",x"986f50",x"855f44",x"835c40",x"755139",x"704c35",x"966d4d",x"9e7453",x"9e7453",x"8c6345",x"895f42",x"8a6041",x"8c6346",x"7d553a",x"8b6143",x"8f6648",x"8d6345",x"8c6343",x"8a6041",x"916748",x"926849",x"926647",x"916647",x"8d6346",x"906747",x"885f42",x"936747",x"7e593f",x"8a6548",x"73533b",x"5d432f",x"4e3929",x"4e3929",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"51483e",x"51483e",x"43382e",x"4d2f1a",x"4d2f1a",x"2f1a0b",x"150e07",x"150e07",x"150e07",x"442611",x"3f2411",x"3f230f",x"39200e",x"391f0e",x"3a200e",x"3c230f",x"412612",x"3b200e",x"3b210e",x"3d220f",x"1a1008",x"785339",x"926749",x"986c4d",x"986d4c",x"906648",x"6f4c37",x"865d40",x"906548",x"8f6446",x"8e6446",x"865c41",x"926a4b",x"8f6649",x"9c7353",x"976f4f",x"996f50",x"8c6547",x"7d583e",x"7b563c",x"886144",x"7e583c",x"956c4d",x"966c4d",x"8b6245",x"916749",x"8d6446",x"90674a",x"9e7351",x"966b4c",x"987150",x"9b6f4e",x"885f43",x"734f36",x"79543a",x"7b533a",x"7c573c",x"74523a",x"483322",x"483322",x"483322",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"37210e",x"37210e",x"281909",x"211508",x"201408",x"201408",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503321",x"503321",x"3a1f0d",x"3b200e",x"371d0c",x"3f2410",x"3b210f",x"381f0d",x"3c2310",x"3d2310",x"402512",x"3e2310",x"40230f",x"27160a",x"27160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"2a180b",x"2c190b",x"371e0d",x"573c2b",x"29190e",x"3a322a",x"150e07",x"150e07",x"150e07",x"150e07",x"24150a",x"150e07",x"150e07",x"150e07",x"1a1008",x"2e1a0b",x"24160a",x"312419",x"312419",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"303030",x"333333",x"313131",x"323232",x"363636",x"434343",x"4d4d4d",x"565656",x"616161",x"3b3b3b",x"333333",x"323232",x"313131",x"333333",x"343434",x"363636",x"3a3a3a",x"3b3b3b",x"444444",x"333333",x"505050",x"454545",x"424242",x"3f3f3f",x"414141",x"424242",x"474747",x"434343",x"4f4f4f",x"4d4d4d",x"474747",x"3e3e3e",x"3d3d3d",x"3c3c3c",x"363636",x"474747",x"474747",x"5a5a5a",x"3c3c3c",x"3e3e3e",x"373737",x"434343",x"454341",x"53504c",x"333333",x"333333",x"323232",x"313131",x"323232",x"2f2f2f",x"2f2f2f",x"3c3c3c",x"3b3b3b",x"3f3f3f",x"323232",x"333333",x"313131",x"313131",x"333333",x"665f57",x"645d57",x"66605a",x"655f59",x"655f5a",x"6c645e",x"66615c",x"66605c",x"69645f",x"645e59",x"605a55",x"635d57",x"000000",x"000000",x"000000",x"4f4f4f",x"4e4e4e",x"484747",x"434343",x"505050",x"3a3a3a",x"343434",x"383838",x"3d3d3d",x"393939",x"333333",x"323232",x"323232",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4949",x"3f3f3f",x"3b3b3b",x"323232",x"313231",x"4f4f4f",x"3a3a3a",x"444444",x"5f5f5f",x"565656",x"353535",x"353535",x"000000",x"414140",x"3e3e3d",x"40403f",x"474747",x"5a5755",x"65615b",x"474645",x"363636",x"313131",x"57524e",x"5c5854",x"5d5955",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3c291c",x"3c291c",x"371d0c",x"3d220f",x"361f0e",x"36200f",x"381f0d",x"3d2310",x"231509",x"382210",x"3b210f",x"452812",x"29180b",x"27160a",x"666463",x"666463",x"5d5045",x"6a635c",x"5c544c",x"676059",x"6a645d",x"756f69",x"756f6a",x"746f69",x"706b65",x"78726c",x"75706b",x"726d68",x"706c67",x"736f6b",x"595959",x"525252",x"535353",x"515150",x"605b56",x"504d4a",x"323232",x"585858",x"6b6a6a",x"6b6764",x"605c58",x"444444",x"303030",x"313131",x"363636",x"424242",x"424242",x"494949",x"494848",x"44413e",x"504a45",x"615a54",x"6c655f",x"5d5853",x"454342",x"2e2e2e",x"2b2b2b",x"2d2d2d",x"2d2d2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c372b",x"4c372b",x"512f16",x"28180b",x"26170b",x"412713",x"3d2411",x"381f0e",x"3b2210",x"3d2411",x"150e07",x"331d0d",x"351e0d",x"3a2110",x"4d2c15",x"432611",x"3e2310",x"281408",x"452813",x"150e07",x"331d0e",x"361f0e",x"402511",x"4c2d16",x"150e07",x"323232",x"323232",x"313131",x"333333",x"333333",x"323232",x"343434",x"333333",x"303030",x"323130",x"323232",x"323131",x"323232",x"323232",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"383838",x"3a3a3a",x"373737",x"323232",x"2f2f2f",x"303030",x"323232",x"2a2a2a",x"323232",x"2f2f2f",x"303030",x"2a2a2a",x"292929",x"1c1c1c",x"353535",x"343434",x"333333",x"323232",x"2f2f2f",x"333333",x"313131",x"313131",x"333333",x"444444",x"343434",x"343434",x"000000",x"000000",x"4d3627",x"4d3627",x"26160a",x"3e220f",x"351d0d",x"341d0c",x"3e2310",x"150e07",x"301c0d",x"361e0d",x"381f0d",x"150e07",x"150e07",x"000000",x"000000",x"1b1008",x"1b1008",x"221409",x"2e1a0c",x"321c0c",x"341d0d",x"311b0b",x"321c0c",x"251509",x"39200d",x"422d20",x"472914",x"412714",x"402513",x"3b2110",x"381f0f",x"27170b",x"6e4932",x"916949",x"93694a",x"90674a",x"9e7554",x"9c7252",x"976c4d",x"9a6f4f",x"8f6649",x"977050",x"986b4b",x"93694a",x"a17655",x"986e4e",x"976c4c",x"926849",x"8d6346",x"996f4f",x"956c4c",x"9d7352",x"976b4c",x"875e41",x"885f43",x"845c3f",x"795238",x"916748",x"956949",x"936849",x"976c4d",x"845c3e",x"9b6f4e",x"896245",x"966b4a",x"93694a",x"946949",x"875f43",x"684531",x"825c41",x"8f6647",x"8b6548",x"654632",x"563d2c",x"4f3a29",x"4f3a29",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4e443a",x"4e443a",x"453a30",x"502d19",x"502d19",x"2e1a0b",x"150e07",x"150e07",x"150e07",x"4a2a13",x"432712",x"412510",x"3c210f",x"351d0d",x"3c210e",x"412611",x"3d2310",x"3c210e",x"3b200e",x"341c0c",x"1f1309",x"805a3f",x"7d593d",x"986e4f",x"95694a",x"966b4c",x"966d4d",x"8b6142",x"865d41",x"8b6143",x"906748",x"734e36",x"684630",x"865d41",x"9d7251",x"9b7354",x"996f4f",x"92694b",x"91684a",x"7d573e",x"846044",x"7d563b",x"936b4d",x"8a6144",x"845d40",x"8c6346",x"946a4a",x"896042",x"9c7150",x"956b4a",x"9c6f4e",x"966d4f",x"8b6143",x"906548",x"896043",x"775036",x"815b40",x"6c4b34",x"463121",x"483222",x"483222",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c230f",x"3c230f",x"2f1e0a",x"291a09",x"251709",x"251709",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503422",x"503422",x"41240f",x"391f0d",x"381f0e",x"3f2411",x"381f0e",x"361e0d",x"422612",x"3d2310",x"3e2310",x"3b210f",x"492913",x"28170a",x"28170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"241509",x"2c190b",x"321b0c",x"523828",x"2d1c10",x"39322a",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"150e07",x"150e07",x"351e0f",x"26170b",x"30251c",x"30251c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b3b3b",x"3b3b3b",x"3e3e3e",x"3c3c3c",x"393939",x"424242",x"515151",x"525252",x"606060",x"626262",x"383838",x"323232",x"333333",x"343434",x"333333",x"383838",x"363636",x"3a3a3a",x"3f3f3f",x"444444",x"3f3f3f",x"323232",x"434343",x"444444",x"444444",x"484848",x"505050",x"5a5a5a",x"575757",x"585654",x"58534f",x"4b4b4b",x"4d4d4d",x"4c4c4c",x"4d4d4d",x"4d4d4d",x"4d4d4d",x"525252",x"393939",x"3a3a3a",x"414141",x"383838",x"000000",x"000000",x"393939",x"393939",x"343434",x"333333",x"313131",x"2f2f2f",x"545454",x"4d4d4d",x"4f4f4f",x"4f4f4f",x"4b4b4b",x"525252",x"4b4b4b",x"383838",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434343",x"333333",x"333333",x"373737",x"363636",x"313131",x"333333",x"404040",x"4f4f4f",x"4d4d4d",x"4d4d4d",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"383838",x"4e4e4e",x"515151",x"5a5a5a",x"5f5f5f",x"3c3c3c",x"323232",x"333333",x"000000",x"000000",x"000000",x"444444",x"474747",x"645f5a",x"69625c",x"474645",x"434342",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"322318",x"322318",x"371e0d",x"3d220f",x"3b210f",x"3a2210",x"351e0d",x"371e0d",x"201309",x"38200e",x"3c230f",x"432611",x"251509",x"26160a",x"51504e",x"51504e",x"726b65",x"6a625b",x"7a756f",x"69635c",x"685f59",x"635b53",x"6e6760",x"6e6862",x"716c66",x"6d6761",x"5b534b",x"595149",x"574f48",x"625c58",x"595959",x"484848",x"444444",x"3d3b39",x"5d554e",x"2f2c28",x"323232",x"5d5d5d",x"4a4847",x"66615c",x"5a5855",x"585858",x"3a3a3a",x"3d3d3c",x"4e4e4e",x"494848",x"313131",x"343333",x"3f3d3b",x"4d4945",x"565049",x"5c544c",x"5c544d",x"4c4641",x"3a3937",x"343434",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513d31",x"513d31",x"533116",x"1c1108",x"2a190b",x"412612",x"3e2511",x"361f0e",x"432713",x"3f2511",x"150e07",x"341d0d",x"331d0d",x"402512",x"543118",x"3e2310",x"381f0e",x"29170a",x"422612",x"201309",x"2d1a0c",x"341d0d",x"3a210f",x"4a2c15",x"383736",x"606060",x"3e3e3e",x"343434",x"313131",x"323232",x"333333",x"323232",x"323232",x"333333",x"323232",x"424242",x"434343",x"363636",x"323232",x"323232",x"333333",x"323232",x"313131",x"444444",x"353535",x"353535",x"313131",x"313131",x"323232",x"2f2f2f",x"303030",x"323232",x"2a2a2a",x"323232",x"2f2f2f",x"303030",x"2a2a2a",x"292929",x"1c1c1c",x"353535",x"343434",x"333333",x"323232",x"2f2f2f",x"333333",x"313131",x"313131",x"333333",x"444444",x"343434",x"343434",x"000000",x"000000",x"4e3829",x"4e3829",x"28170b",x"3f2310",x"331d0d",x"2f1b0c",x"3c220f",x"341c0c",x"27170b",x"38200e",x"371f0e",x"150e07",x"150e07",x"000000",x"000000",x"1a1008",x"1a1008",x"211409",x"2e1a0c",x"321c0c",x"361e0d",x"311a0b",x"2f1a0b",x"25160a",x"361e0d",x"483426",x"482b16",x"422815",x"3f2413",x"3c2412",x"3c2211",x"321d0e",x"5c361c",x"855f43",x"886043",x"956c4c",x"a27856",x"9c7050",x"9c704f",x"996e4e",x"9b7050",x"946e4f",x"8f6546",x"936a4c",x"9a6f4e",x"9b7050",x"976d4c",x"926949",x"936949",x"9a6f4f",x"9b7151",x"906748",x"976b4b",x"865d40",x"8e6345",x"845b3f",x"754f36",x"956b4c",x"916648",x"996d4c",x"966a4b",x"865d3f",x"966c4c",x"8e6445",x"9c704f",x"916748",x"906546",x"8a6043",x"845b3f",x"825b3f",x"8b6043",x"866144",x"715138",x"5b412d",x"4f3a29",x"4f3a29",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4f463c",x"4f463c",x"42372e",x"4b2d19",x"4b2d19",x"381e0c",x"150e07",x"150e07",x"150e07",x"462812",x"3c220f",x"3e2310",x"3e230f",x"30190b",x"3b200e",x"3f2410",x"3e2310",x"3c210f",x"3b200e",x"3b200e",x"1d1108",x"8a6446",x"815b3f",x"96694b",x"916546",x"7b573d",x"8b6345",x"885e41",x"8f6445",x"996d4c",x"996d4d",x"794f34",x"714e37",x"896145",x"845c40",x"a07454",x"996e4e",x"8a6245",x"855d42",x"8a6144",x"7a5a3f",x"81593e",x"90694a",x"8d6648",x"8f6446",x"8b6245",x"91684a",x"885f41",x"94694a",x"9b7050",x"9d7050",x"926748",x"8b6244",x"896043",x"8b6345",x"6f4c32",x"7b583d",x"664630",x"452f20",x"463020",x"463020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b220f",x"3b220f",x"311f0a",x"2b1b09",x"271909",x"271909",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503422",x"503422",x"432511",x"371e0d",x"3e2310",x"3f2310",x"361e0d",x"3b210f",x"38200f",x"412511",x"412511",x"39200e",x"472812",x"2b180b",x"2b180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"201309",x"2d190b",x"381e0d",x"593f2e",x"2a1a0f",x"3a322a",x"150e07",x"150e07",x"150e07",x"150e07",x"191008",x"150e07",x"150e07",x"150e07",x"1d1108",x"351f0f",x"28170c",x"32271d",x"32271d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5b5b5b",x"515151",x"4e4e4e",x"4a4a4a",x"3c3c3c",x"4b4b4b",x"575757",x"595959",x"5d5d5d",x"646464",x"414141",x"323232",x"323232",x"333333",x"333333",x"3c3c3c",x"444444",x"434343",x"464646",x"494949",x"484848",x"494a4a",x"4d4d4d",x"484848",x"4d4d4d",x"656565",x"4d4d4d",x"454545",x"454545",x"585654",x"353535",x"343434",x"4d4d4d",x"595959",x"525252",x"4f4f4f",x"5d5d5d",x"343434",x"363636",x"393939",x"000000",x"000000",x"000000",x"000000",x"555555",x"555555",x"636363",x"6c6c6c",x"5f5f5f",x"575757",x"545454",x"545454",x"535353",x"565656",x"515151",x"545454",x"515151",x"5d5d5d",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"414141",x"414141",x"343434",x"4d4d4d",x"4a4a4a",x"3e3e3e",x"313131",x"4e4e4e",x"484848",x"303030",x"323232",x"383838",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595858",x"595858",x"717171",x"525252",x"5f5a55",x"454545",x"575452",x"373635",x"373635",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"352419",x"352419",x"3a200e",x"3a200e",x"3b210f",x"351f0e",x"371e0d",x"39200e",x"201308",x"351d0d",x"3a210f",x"442711",x"211409",x"25150a",x"595756",x"595756",x"605850",x"736d66",x"726c66",x"5c544b",x"5d544b",x"5a5148",x"5f574f",x"5d564d",x"5e564f",x"5a5148",x"574f47",x"4e463d",x"4f473e",x"534c45",x"2b2a29",x"313131",x"343333",x"423f3c",x"5c544c",x"272421",x"313131",x"313131",x"433f3c",x"5a544c",x"383634",x"333333",x"313131",x"2e2e2d",x"383838",x"303030",x"2c2c2c",x"383736",x"3b3631",x"48423b",x"59514a",x"5f574e",x"59524b",x"494540",x"333231",x"313131",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d382b",x"4d382b",x"482913",x"28170b",x"29180b",x"39200f",x"3b2210",x"341d0d",x"3d2311",x"3f2512",x"150e07",x"321d0d",x"2d190b",x"412612",x"492a14",x"341d0d",x"331c0c",x"361d0c",x"442713",x"402612",x"2b190b",x"351d0d",x"39200e",x"4b2c15",x"333333",x"313131",x"323232",x"323232",x"555555",x"454545",x"5c5c5c",x"595959",x"323232",x"333333",x"323232",x"434343",x"454545",x"5e5e5e",x"606060",x"5b5b5b",x"525252",x"505050",x"4b4b4b",x"383838",x"323232",x"343434",x"323232",x"323232",x"323232",x"515151",x"323232",x"333333",x"323232",x"333333",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"333333",x"323232",x"323232",x"313131",x"333231",x"282828",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c372a",x"4c372a",x"27160a",x"3c210f",x"361e0d",x"321c0c",x"341d0d",x"371f0d",x"150e07",x"351d0d",x"3f230f",x"150e07",x"150e07",x"000000",x"000000",x"1a1008",x"1a1008",x"211309",x"2d190b",x"301a0b",x"371f0d",x"301a0b",x"361e0d",x"251509",x"3b200e",x"4e3627",x"482a16",x"432814",x"3e2413",x"3f2513",x"371f10",x"27170b",x"69442f",x"7c5940",x"825b3f",x"8c6346",x"986f4e",x"926849",x"986d4e",x"936749",x"966b4c",x"9b7453",x"956949",x"966d4f",x"9d7253",x"986e4e",x"956b4b",x"976b4c",x"966b4b",x"8e684a",x"9b7050",x"9d704d",x"845e43",x"825a3e",x"926747",x"8c6243",x"83593d",x"956b4c",x"916748",x"906747",x"916646",x"734b31",x"976c4c",x"8f6647",x"9a6f4f",x"906648",x"875d40",x"885e42",x"8a6143",x"8c6243",x"855e40",x"866043",x"78563c",x"5d432e",x"4e3928",x"4e3928",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1c1108",x"1c1108",x"150e07",x"150e07",x"150e07",x"50473d",x"50473d",x"3d332a",x"4a2e1c",x"4a2e1c",x"381f0d",x"150e07",x"150e07",x"150e07",x"432611",x"412410",x"3f2410",x"381f0e",x"3a200e",x"3c220f",x"361f0e",x"3b210f",x"3c220f",x"381f0d",x"3a1f0d",x"201308",x"7e573c",x"815a3f",x"956a49",x"8f6545",x"94694a",x"926748",x"845c3f",x"885f43",x"896042",x"92684a",x"845b3d",x"8b6245",x"7d593f",x"9b7051",x"9f7454",x"8f6547",x"936a4c",x"845c40",x"805b40",x"8b6346",x"80593f",x"8e6546",x"9e7454",x"8d6346",x"916749",x"966d4d",x"996e4e",x"9d7050",x"9f7352",x"9d7150",x"946a4a",x"815a3d",x"906647",x"845d41",x"6f4a31",x"6e4d35",x"6b4a34",x"432e1e",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"35200d",x"35200d",x"301e0a",x"281909",x"231608",x"231608",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"553827",x"553827",x"432511",x"331c0c",x"3f230f",x"3d2310",x"3a200e",x"3a200e",x"3f2411",x"402511",x"422712",x"351e0d",x"432611",x"311c0d",x"311c0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"341d0d",x"381d0d",x"523828",x"2a1a0d",x"3c342c",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"150e07",x"150e07",x"150e07",x"150e07",x"2f1c0e",x"26170c",x"2d221a",x"2d221a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"59524b",x"59524b",x"686868",x"656565",x"565656",x"636363",x"636262",x"636363",x"626261",x"666666",x"535353",x"3c3c3c",x"333333",x"373737",x"555555",x"575757",x"575757",x"636363",x"5f5f5f",x"5c5c5c",x"5c5c5c",x"595959",x"585858",x"686461",x"676360",x"565655",x"434343",x"464646",x"454545",x"000000",x"383838",x"434343",x"494949",x"5b5b5b",x"646464",x"5c5c5c",x"353535",x"363636",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"555555",x"585858",x"484848",x"424242",x"3a3938",x"555555",x"626262",x"5f5f5f",x"676767",x"5a5a5a",x"575757",x"555555",x"4d4c4a",x"464646",x"333232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"474747",x"474747",x"4b4b4b",x"4d4d4d",x"4a4a4a",x"4d4d4d",x"636363",x"505050",x"515151",x"333434",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595858",x"5f5e5e",x"696765",x"56524e",x"6d6761",x"6e6862",x"66625d",x"414141",x"373635",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2c2018",x"2c2018",x"3f230f",x"3a200e",x"3b210e",x"3d2410",x"3a200e",x"371e0d",x"251509",x"361f0e",x"39200f",x"432712",x"1c1108",x"25150a",x"25150a",x"5a5856",x"414141",x"504e4d",x"545251",x"5d5a58",x"585551",x"5a5754",x"595652",x"5b5957",x"535353",x"515151",x"575654",x"555352",x"5a5958",x"575656",x"4f4e4d",x"555453",x"5b5957",x"575655",x"4d4c4c",x"515151",x"4f4f4f",x"494949",x"3f3f3f",x"353535",x"333333",x"494949",x"525252",x"545352",x"484746",x"484746",x"585452",x"585858",x"393939",x"353535",x"474747",x"4b4b4b",x"333333",x"303030",x"2f2f2f",x"333333",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3528",x"4a3528",x"522f17",x"23150a",x"1d1208",x"3b2210",x"3b2210",x"37200f",x"3c2310",x"3b2210",x"150e07",x"351e0e",x"2d190b",x"3e2411",x"533017",x"3d220f",x"341d0d",x"321c0c",x"452814",x"452914",x"28170a",x"371f0e",x"3f2311",x"442712",x"150e07",x"333333",x"333333",x"313131",x"343434",x"383838",x"3c3b39",x"494949",x"494949",x"4b4b4b",x"414141",x"3f3f3f",x"515151",x"525252",x"3f3e3d",x"333333",x"313131",x"303030",x"323232",x"3c3c3c",x"333232",x"323130",x"323232",x"3b3a38",x"423f3d",x"515151",x"323232",x"333333",x"323232",x"333333",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"333333",x"323232",x"323232",x"313131",x"333231",x"282828",x"2a2a2a",x"2a2a2a",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3a2d",x"4e3a2d",x"231409",x"39200e",x"381f0e",x"39200e",x"371e0d",x"381f0e",x"150e07",x"331d0d",x"38200e",x"180f07",x"180f07",x"000000",x"000000",x"1a1008",x"1a1008",x"201309",x"2e1a0c",x"321c0c",x"39200e",x"2e190b",x"311b0b",x"25150a",x"351d0d",x"4b3628",x"452815",x"422816",x"412714",x"3d2512",x"3e2513",x"331e0f",x"5c3a27",x"7e593f",x"81593e",x"976d4d",x"986e4f",x"996c4c",x"9b6f4e",x"8d6548",x"93684a",x"a37856",x"936849",x"9b7150",x"9b7151",x"966d4e",x"9b6f4f",x"9c7050",x"986c4c",x"976b4a",x"9e7351",x"a37756",x"946949",x"8b6144",x"906648",x"916547",x"81583c",x"9b6f4e",x"936849",x"8f6747",x"916748",x"70472d",x"926748",x"8b6042",x"956b4c",x"8f6445",x"8d6345",x"8e6344",x"8a6144",x"865d41",x"845d3f",x"845e42",x"75533b",x"604530",x"513a29",x"513a29",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341e0e",x"341e0e",x"150e07",x"150e07",x"150e07",x"51473d",x"51473d",x"3c3229",x"4e2d17",x"4e2d17",x"311c0d",x"150e07",x"150e07",x"150e07",x"3f220f",x"412511",x"3d220f",x"3f230f",x"3c220f",x"39200f",x"351e0d",x"3e2310",x"3e230f",x"371d0c",x"3b200d",x"201308",x"865f41",x"855e41",x"9f7152",x"936849",x"8f6447",x"8b6446",x"815b3e",x"865d40",x"8e6344",x"8a6346",x"8e6445",x"8d6548",x"966c4d",x"996e4e",x"9c7150",x"8e6545",x"956c4c",x"865c3f",x"8e6547",x"906748",x"855e42",x"886146",x"9a7150",x"986d4e",x"976d4d",x"825b3f",x"926749",x"9b704f",x"956c4c",x"9e7351",x"926849",x"80593e",x"93694a",x"855d41",x"744f36",x"755138",x"6f4d35",x"442f1f",x"442f1f",x"442f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200e",x"38200e",x"2e1d0a",x"281909",x"281909",x"281909",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513524",x"513524",x"422510",x"341c0c",x"39200e",x"3c210f",x"381f0d",x"381f0e",x"3a2210",x"39200f",x"3f2511",x"361d0d",x"432611",x"29170b",x"29170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"311c0d",x"371d0c",x"4f3424",x"27170c",x"423a31",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"150e07",x"2b1a0d",x"29180c",x"271d15",x"271d15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"59524b",x"59524b",x"5e564f",x"655e58",x"6f6a64",x"716c67",x"69625c",x"6b655f",x"6e6762",x"6b655f",x"74706b",x"6d6762",x"716b65",x"65625e",x"666360",x"6a6663",x"6e6b68",x"716e6a",x"75706c",x"6b6765",x"736f6a",x"6e6a67",x"706b66",x"716c67",x"676360",x"5f5d5c",x"504f4f",x"000000",x"000000",x"000000",x"000000",x"444444",x"505050",x"5d5a58",x"5f5b56",x"58524c",x"373736",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434242",x"40403f",x"444341",x"514d4a",x"57524f",x"605953",x"625b54",x"5f5954",x"5b554f",x"534e49",x"4c4947",x"585858",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b4b4b",x"4d4d4d",x"605f5d",x"5f5b58",x"5d5956",x"595654",x"3d3d3d",x"585755",x"444444",x"444444",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"696765",x"56524e",x"000000",x"6e6862",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2a2019",x"2a2019",x"3d230f",x"371e0d",x"381f0e",x"351f0e",x"361e0d",x"321b0b",x"28170a",x"361f0e",x"361f0e",x"412410",x"28170a",x"241509",x"241509",x"313131",x"313131",x"5a524a",x"5d554d",x"5d564e",x"5c544d",x"5b534b",x"625952",x"635b54",x"625b53",x"655e57",x"635c55",x"625b55",x"68615a",x"59534d",x"59524c",x"58514b",x"57493d",x"565049",x"454341",x"434343",x"3b3b3a",x"3b3b3a",x"333333",x"333333",x"333333",x"484848",x"525252",x"575350",x"494540",x"4e4b49",x"625c55",x"525150",x"333333",x"313131",x"35312e",x"393939",x"323232",x"323232",x"323232",x"2f2f2f",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"493326",x"493326",x"4f2d15",x"29180b",x"1d1108",x"422713",x"361f0e",x"2e1b0d",x"341e0e",x"392110",x"1d1209",x"331e0e",x"361f0e",x"452914",x"543017",x"3d220f",x"3b210f",x"26160a",x"3a2110",x"150e07",x"27160a",x"331d0d",x"39210f",x"422511",x"150e07",x"4f4f4f",x"323232",x"333333",x"525252",x"616161",x"505050",x"353535",x"333333",x"333333",x"313131",x"323232",x"323232",x"323232",x"353535",x"313131",x"323232",x"323232",x"343434",x"363636",x"303030",x"343434",x"323232",x"3b3a38",x"3e3b39",x"4e4e4e",x"323232",x"333333",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"303030",x"333333",x"282828",x"2a2a2a",x"2a2a2a",x"000000",x"000000",x"000000",x"000000",x"000000",x"483121",x"483121",x"26160a",x"3c210f",x"3a210f",x"2d190b",x"3a200e",x"371e0d",x"27170a",x"321d0d",x"38200e",x"180f07",x"180f07",x"000000",x"000000",x"191008",x"191008",x"211309",x"2c190b",x"2d190b",x"361d0d",x"301a0b",x"351d0d",x"25150a",x"38200f",x"443327",x"472b16",x"412615",x"3f2614",x"3f2614",x"422714",x"2d1a0d",x"64412d",x"9d7050",x"8b6143",x"8e6546",x"8e6446",x"956a4b",x"9b7050",x"a17453",x"976b4c",x"a07453",x"986d4c",x"966b4b",x"9a6e4c",x"9b7252",x"956a4b",x"936949",x"9b6e4d",x"9d704f",x"9c7151",x"a27655",x"966b4a",x"8c6143",x"865d41",x"8f6446",x"7f563a",x"986c4d",x"9a6d4c",x"966d4d",x"906547",x"835b3d",x"906647",x"916747",x"996e4e",x"8d6244",x"906648",x"8e6344",x"885f42",x"875e41",x"8b6244",x"8e6649",x"7b573d",x"654733",x"4f3928",x"4f3928",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402511",x"402511",x"150e07",x"150e07",x"150e07",x"52483e",x"52483e",x"3d342b",x"482a15",x"482a15",x"2f1c0d",x"150e07",x"150e07",x"150e07",x"482712",x"3c210f",x"39200e",x"3c210f",x"371e0d",x"39200e",x"3c210f",x"3c210e",x"3c220f",x"371e0d",x"3a200d",x"1c1108",x"8b6145",x"8b6244",x"9e7252",x"946849",x"926749",x"916646",x"8e6445",x"7f583b",x"946849",x"946b4b",x"8e6545",x"9b7050",x"91684a",x"92684a",x"996f4d",x"8a6144",x"956c4c",x"8b6143",x"9a6d4d",x"986e4f",x"8f6647",x"936b4d",x"875f43",x"8f6648",x"956c4d",x"865e41",x"7e573d",x"966b4c",x"966d4d",x"986f4e",x"976b4c",x"845c3f",x"8e6546",x"865e41",x"7a543a",x"724f36",x"684932",x"4a3323",x"4a3323",x"4a3323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a220f",x"3a220f",x"32200a",x"2d1d0a",x"2c1c09",x"2c1c09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"493021",x"493021",x"432611",x"361d0d",x"361d0d",x"381f0e",x"3a200e",x"351d0c",x"442813",x"38200f",x"442813",x"341d0d",x"3d230f",x"2f1b0c",x"2f1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"3f2411",x"361c0c",x"4f3321",x"21140b",x"4a4239",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"150e07",x"150e07",x"150e07",x"170f07",x"28190d",x"23160b",x"2c1f16",x"2c1f16",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e4e4e",x"4e4e4e",x"353535",x"323232",x"3d3d3d",x"323232",x"333333",x"363636",x"383838",x"404040",x"313131",x"323232",x"313131",x"2e2e2e",x"323232",x"2b2b2b",x"313131",x"323232",x"2f2f2f",x"323232",x"313232",x"323232",x"3a3a3a",x"393939",x"404040",x"383838",x"323232",x"323232",x"000000",x"000000",x"323232",x"323232",x"323232",x"303030",x"343434",x"313131",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"333333",x"323232",x"343434",x"303030",x"2f2f2f",x"333333",x"323232",x"323232",x"313131",x"323232",x"2f2f2f",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"373737",x"313131",x"313131",x"323232",x"313131",x"323232",x"323232",x"313131",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"313131",x"333333",x"313131",x"323232",x"333232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2c221b",x"2c221b",x"402410",x"361e0d",x"341d0d",x"2d1a0c",x"331c0c",x"29160a",x"191008",x"2f1b0c",x"331e0e",x"412410",x"201309",x"241609",x"241609",x"363636",x"323232",x"615951",x"605850",x"5f5850",x"655e57",x"5f574f",x"615951",x"665f58",x"69625a",x"6a635c",x"59524a",x"5b544d",x"6f6963",x"5a534d",x"5b544e",x"5c5650",x"5e5852",x"5d564e",x"383635",x"3e3e3d",x"414140",x"343434",x"323232",x"313131",x"313131",x"666666",x"474747",x"514b46",x"413e3a",x"504d4a",x"5f5850",x"373636",x"333333",x"323232",x"333333",x"363636",x"323232",x"323233",x"313131",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3729",x"4d3729",x"4e2d15",x"2a190b",x"24150a",x"402612",x"341e0e",x"341e0e",x"3b2211",x"2f1c0d",x"150e07",x"351f0f",x"311c0d",x"452914",x"543219",x"3c220f",x"381f0e",x"150e07",x"37200f",x"150e07",x"1a1008",x"331d0d",x"3a210f",x"412511",x"323232",x"3e3e3e",x"555555",x"4f4f4f",x"616161",x"545454",x"5d5d5d",x"5f5e5e",x"323232",x"515151",x"323232",x"333232",x"323232",x"525252",x"5f5f5f",x"5b5b5b",x"585857",x"434343",x"323232",x"323232",x"2a2a2a",x"303030",x"323232",x"3f3d3a",x"3e3c3a",x"4c4c4c",x"313131",x"2f2f2f",x"323232",x"333333",x"333333",x"343434",x"323232",x"2f2f2f",x"343434",x"323232",x"323232",x"323232",x"313131",x"333333",x"353535",x"323232",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"473123",x"473123",x"2b180b",x"3a200f",x"3a210f",x"150e07",x"2f1a0b",x"150e07",x"150e07",x"2f1b0c",x"3a220f",x"180f07",x"180f07",x"000000",x"000000",x"1a1008",x"1a1008",x"221409",x"2c190b",x"311b0c",x"321c0c",x"2f190b",x"341d0d",x"25150a",x"38200e",x"3e2f24",x"472915",x"412716",x"432816",x"3d2514",x"3e2514",x"2a180b",x"7e563b",x"9a6e4f",x"875f43",x"895f43",x"976b4b",x"996c4c",x"9d7051",x"986d4c",x"8e6448",x"9d7453",x"9b6f4f",x"94694a",x"966949",x"996e4f",x"996d4d",x"93684a",x"996d4c",x"9e7251",x"a27655",x"a27755",x"956949",x"8f6547",x"946849",x"8b6144",x"7e553a",x"906648",x"8f6647",x"9b7150",x"956b4a",x"855c3f",x"8a6143",x"946848",x"966a4a",x"8d6546",x"936749",x"80593c",x"8b6244",x"8a6042",x"8b6244",x"8b6447",x"7a563b",x"5c422d",x"4e3827",x"4e3827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2310",x"3d2310",x"150e07",x"150e07",x"150e07",x"52483f",x"52483f",x"41372e",x"4e2f1b",x"4e2f1b",x"371f0e",x"150e07",x"150e07",x"150e07",x"422511",x"3a200e",x"3b200f",x"3b220f",x"341d0c",x"371f0e",x"39200e",x"39200e",x"402410",x"381e0d",x"3b210e",x"201309",x"8c6446",x"8b6143",x"946b4d",x"8b6143",x"906648",x"815940",x"885e41",x"865d3f",x"8e6345",x"8f6546",x"8e6445",x"986e50",x"956c4c",x"95694a",x"9b6f4f",x"855d3f",x"896245",x"8e6447",x"966a4b",x"976d4e",x"93694a",x"946b4c",x"896144",x"7e583d",x"896144",x"906647",x"7b553b",x"966c4c",x"8e684a",x"9a7151",x"8f6547",x"885f41",x"8f6547",x"855d3f",x"754f36",x"755238",x"644630",x"47301f",x"473020",x"473020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"39210d",x"39210d",x"311f0a",x"2d1d0a",x"2a1b09",x"2a1b09",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f3423",x"4f3423",x"442812",x"361d0c",x"391f0e",x"3b210f",x"3c210f",x"351d0d",x"442813",x"3a210f",x"412612",x"331c0c",x"452711",x"2d1a0b",x"2d1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"452913",x"331b0a",x"543724",x"28190e",x"443b33",x"150e07",x"150e07",x"150e07",x"150e07",x"28170b",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1b0d",x"23150b",x"261e17",x"261e17",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595959",x"595959",x"5d5d5d",x"545454",x"434343",x"4d4d4d",x"535353",x"5b5b5b",x"656565",x"575757",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"383838",x"373737",x"3c3c3c",x"3c3c3c",x"393939",x"3d3d3d",x"404040",x"464646",x"464646",x"3d3d3d",x"323232",x"333333",x"323232",x"333333",x"323232",x"333333",x"383838",x"323232",x"333333",x"393939",x"343434",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"313131",x"3b3b3b",x"464646",x"424242",x"383838",x"343434",x"323232",x"313131",x"343434",x"323232",x"343434",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d3d3d",x"3d3d3d",x"4f4f4f",x"494949",x"3d3d3d",x"323232",x"363636",x"4b4b4b",x"343434",x"323232",x"333333",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"313131",x"323232",x"313131",x"323232",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"35251a",x"35251a",x"3f2410",x"311b0c",x"221409",x"361f0e",x"150e07",x"211308",x"150e07",x"170f07",x"2b180b",x"3b220f",x"241509",x"26160a",x"26160a",x"4e4d4d",x"454543",x"615951",x"5e564e",x"625b53",x"655e57",x"5e564e",x"615a53",x"645c55",x"655e57",x"665e57",x"5d574f",x"69635c",x"6f6962",x"514b44",x"564f48",x"5c564f",x"605952",x"5b534c",x"373636",x"3e3d3d",x"3b3b3a",x"313131",x"343434",x"333333",x"323232",x"606060",x"3c3c3b",x"504b45",x"3e3a37",x"605c58",x"6f6964",x"303030",x"323232",x"303030",x"313131",x"333333",x"333333",x"333333",x"313131",x"313131",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3729",x"4d3729",x"512f16",x"28180b",x"1c1108",x"402512",x"29180b",x"37200f",x"150e07",x"1a1008",x"150e07",x"150e07",x"28170a",x"3b210f",x"4f2f17",x"321c0d",x"3a210f",x"381f0e",x"2c190b",x"301c0d",x"351f0e",x"2c190b",x"3b210f",x"472913",x"323232",x"323232",x"323232",x"313131",x"343434",x"343434",x"343434",x"313131",x"323232",x"323232",x"303030",x"333333",x"323232",x"313131",x"323232",x"313131",x"313131",x"333333",x"323232",x"333130",x"333130",x"323232",x"333333",x"403e3a",x"312f2e",x"454545",x"323232",x"303030",x"333333",x"343434",x"333333",x"313131",x"323232",x"2f2f2f",x"323232",x"323232",x"2d2d2d",x"313131",x"323232",x"313131",x"313131",x"313131",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3626",x"4e3626",x"28170a",x"3d2310",x"301b0b",x"311b0b",x"341d0d",x"251509",x"301a0b",x"201309",x"3a210f",x"150e07",x"150e07",x"000000",x"000000",x"1a1008",x"1a1008",x"211409",x"2b180b",x"311b0c",x"311b0c",x"2c180a",x"351e0d",x"26160a",x"3e230f",x"3d2f24",x"482a17",x"472c18",x"442915",x"412815",x"3d2414",x"362010",x"724d36",x"a07553",x"9c7050",x"865c3f",x"a27654",x"926647",x"976b4b",x"9a7050",x"8c6245",x"876044",x"9b6f4f",x"95694a",x"976c4c",x"996e4f",x"8f6547",x"906445",x"9c7050",x"a17453",x"966c4d",x"9a704f",x"976b4b",x"946748",x"966a4b",x"8d6344",x"81583d",x"906648",x"926849",x"986f50",x"936a4a",x"825a3d",x"865e41",x"885f42",x"906647",x"976d4d",x"8f6344",x"8a5f41",x"8c6244",x"8f6647",x"865e41",x"896246",x"755138",x"5e422e",x"4e3727",x"4e3727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1a0c",x"2f1a0c",x"150e07",x"150e07",x"150e07",x"51483d",x"51483d",x"42382f",x"4c2f1b",x"4c2f1b",x"2e1b0d",x"150e07",x"150e07",x"150e07",x"452711",x"381f0e",x"3d220f",x"351d0d",x"351d0c",x"38200e",x"311c0b",x"3d230f",x"3f2411",x"361d0c",x"3b200e",x"1a1008",x"79563c",x"906447",x"986d4d",x"795338",x"986e4e",x"896042",x"8a6043",x"8e6445",x"8e6445",x"976c4c",x"936849",x"92694b",x"91694c",x"946a4a",x"966c4d",x"886143",x"8d6548",x"976e4e",x"966a4b",x"936a4b",x"95694a",x"9b7150",x"926749",x"916849",x"8c6345",x"936848",x"926848",x"835d42",x"8a6145",x"966e4e",x"8b6144",x"80583d",x"926749",x"875f41",x"735036",x"745037",x"714f38",x"432e1e",x"422d1d",x"422d1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2310",x"3d2310",x"3c250d",x"8e7355",x"7e664c",x"7e664c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f3321",x"4f3321",x"482913",x"351c0c",x"3c220f",x"381f0e",x"3a200e",x"361e0d",x"422713",x"38200f",x"402511",x"381f0d",x"442611",x"2b190b",x"2b190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"38200f",x"371d0c",x"4d311f",x"2a1a0e",x"423a32",x"150e07",x"150e07",x"150e07",x"150e07",x"29180a",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1a0d",x"27170b",x"29211a",x"29211a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"565656",x"4e4e4e",x"4a4a4a",x"444444",x"3b3b3b",x"444444",x"4d4d4d",x"505050",x"616161",x"5c5c5c",x"2f2f2f",x"343434",x"313131",x"333333",x"333333",x"323232",x"303030",x"313131",x"383838",x"373737",x"383838",x"363636",x"373737",x"3b3b3b",x"393939",x"4a4a4a",x"424242",x"333333",x"323232",x"333333",x"313131",x"313131",x"414141",x"474747",x"414141",x"474747",x"303030",x"313131",x"323232",x"323232",x"313131",x"000000",x"000000",x"000000",x"4a4a4a",x"4a4a4a",x"666666",x"5c5c5c",x"505050",x"4c4c4c",x"505050",x"454545",x"454545",x"474747",x"414141",x"484848",x"4d4d4d",x"575757",x"454545",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"515151",x"515151",x"353535",x"414141",x"3f3f3f",x"4d4d4d",x"4d4d4d",x"454545",x"4d4d4d",x"404040",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383838",x"383838",x"555555",x"424242",x"313131",x"323232",x"303030",x"333333",x"2e2e2e",x"323232",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"2e2720",x"2e2720",x"3b210f",x"321c0c",x"381f0e",x"3b210f",x"341d0d",x"281609",x"341d0c",x"38200e",x"150e07",x"3f2410",x"26160a",x"27170a",x"27170a",x"4b4b4a",x"333333",x"333333",x"333333",x"323232",x"333333",x"323232",x"333333",x"323232",x"2f2f2f",x"333333",x"323232",x"2e2d2d",x"313131",x"313131",x"323232",x"313131",x"333333",x"333333",x"333333",x"313131",x"323232",x"333333",x"333333",x"333333",x"332c29",x"373737",x"333232",x"323232",x"323232",x"303030",x"323232",x"323232",x"2f2f2f",x"323232",x"323232",x"343434",x"6d6c6c",x"484645",x"3f3b37",x"33302d",x"2f2f2f",x"2f2f2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523b2c",x"523b2c",x"523017",x"29190b",x"2b1a0c",x"3b2311",x"39210f",x"402512",x"3c2310",x"22140a",x"3b2210",x"3a210f",x"150e07",x"402511",x"563219",x"3a2210",x"3d2310",x"3b210f",x"150e07",x"311e0e",x"38200f",x"311c0d",x"39200f",x"482a14",x"150e07",x"363636",x"323232",x"323232",x"323232",x"323232",x"464646",x"434141",x"333232",x"323131",x"323232",x"323232",x"333333",x"333333",x"333333",x"343434",x"3a3a3a",x"373737",x"333333",x"333333",x"323232",x"373737",x"323232",x"363636",x"515151",x"646464",x"323232",x"323232",x"313131",x"333333",x"333333",x"313131",x"333333",x"323232",x"323232",x"323232",x"313131",x"4a4a4a",x"3d3d3d",x"363636",x"3f3f3f",x"393939",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"463123",x"463123",x"241509",x"3c210f",x"2d190b",x"321c0c",x"311c0d",x"231409",x"341d0c",x"25160a",x"351d0d",x"150e07",x"150e07",x"000000",x"000000",x"1a1008",x"1a1008",x"231409",x"2d1a0b",x"2f1a0b",x"321b0c",x"2d180a",x"361f0d",x"26160a",x"402511",x"3d2e24",x"472b17",x"3e2515",x"422816",x"432816",x"3a2313",x"2a190c",x"805b3f",x"956b4d",x"9b7151",x"996d4c",x"9d7050",x"9a6d4d",x"9a6e4d",x"9d7151",x"986c4c",x"a27655",x"8d6548",x"946a4c",x"986d4e",x"986e4f",x"916748",x"956b4b",x"916749",x"9a6f50",x"956b4b",x"9d7353",x"93694a",x"906648",x"936949",x"906648",x"82593e",x"946849",x"936a4b",x"99704f",x"936849",x"7f573b",x"956949",x"936748",x"926748",x"9c7050",x"936849",x"875f41",x"825b3f",x"946a4a",x"8a6143",x"7d573f",x"77543a",x"614531",x"4d3726",x"4d3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351f0e",x"351f0e",x"150e07",x"150e07",x"150e07",x"4f453c",x"4f453c",x"382d24",x"4e2e19",x"4e2e19",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"472711",x"371e0d",x"371f0d",x"38200e",x"321b0c",x"351e0d",x"371e0d",x"38200e",x"3c230f",x"351d0c",x"3a200e",x"1f1208",x"896345",x"8d6445",x"95694a",x"8e6445",x"976d4d",x"8f6545",x"845c3f",x"8a6143",x"8e6447",x"8e6345",x"956a4c",x"9c7454",x"8b6347",x"906547",x"90684a",x"8c6546",x"956c4d",x"9b6f50",x"946a4b",x"996f4f",x"93694a",x"966f4f",x"966c4e",x"996e4e",x"976c4c",x"916748",x"966c4d",x"8a6347",x"876044",x"926b4d",x"855d3f",x"825b3f",x"8d6244",x"815a3e",x"734f36",x"805a3e",x"6c4c34",x"402c1d",x"442f1e",x"442f1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2310",x"3d2310",x"3c250d",x"8e7355",x"7e664c",x"7e664c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b3222",x"4b3222",x"442712",x"341c0c",x"3d220f",x"381f0d",x"3b210f",x"381f0e",x"442813",x"412511",x"412612",x"351d0c",x"442611",x"331d0d",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"3f2511",x"391f0e",x"4f3323",x"29190e",x"3b332b",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"150e07",x"150e07",x"150e07",x"170f07",x"2e1b0d",x"27170b",x"30241c",x"30241c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4a4a",x"404040",x"3c3c3c",x"424242",x"373737",x"3c3c3c",x"464646",x"4f4f4f",x"626262",x"606060",x"333333",x"313131",x"323232",x"313131",x"333333",x"343434",x"303030",x"323232",x"363636",x"383838",x"2f2f2f",x"343434",x"323232",x"414141",x"3c3c3c",x"414141",x"414141",x"3f4040",x"4a4a4a",x"4b4b4b",x"444444",x"3e3e3e",x"3f3f3f",x"3c3c3c",x"404040",x"4d4d4d",x"4f4f4f",x"393939",x"303030",x"333333",x"323232",x"2c2c2c",x"2b2b2b",x"000000",x"4a4a4a",x"5a5a5a",x"484848",x"3f3d3b",x"3f3f3f",x"3a3a3a",x"4b4b4b",x"474747",x"4c4c4c",x"4c4c4c",x"4c4c4c",x"545454",x"4f4f4f",x"474747",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"323232",x"323232",x"333333",x"454545",x"3f3f3f",x"4b4b4b",x"4e4e4e",x"4b4b4b",x"525252",x"5b5b5b",x"5d5d5d",x"4b4b4b",x"4b4b4b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"313131",x"323232",x"545454",x"303030",x"4f4f4f",x"444444",x"323232",x"323232",x"323232",x"000000",x"000000",x"323232",x"333333",x"333333",x"323232",x"323232",x"343434",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"362e26",x"362e26",x"3d220f",x"3a200e",x"3a200e",x"3f2411",x"38200e",x"341d0c",x"2d190b",x"3c2210",x"150e07",x"3f2411",x"28170a",x"24150a",x"24150a",x"333333",x"333333",x"343434",x"333333",x"323232",x"333333",x"333333",x"303030",x"2d2d2d",x"2f2f2f",x"343434",x"323232",x"313131",x"303030",x"313131",x"333333",x"323232",x"313131",x"333333",x"323232",x"303030",x"303030",x"313131",x"323232",x"323232",x"313131",x"322f2d",x"313131",x"323232",x"323232",x"333333",x"313131",x"2c2c2c",x"303030",x"323232",x"303030",x"333333",x"686867",x"4f4d4a",x"45413d",x"3a3836",x"2e2e2e",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543d2e",x"543d2e",x"4c2c15",x"2a190b",x"301c0d",x"341d0d",x"3b210f",x"422612",x"38200f",x"38200f",x"341f0f",x"3e2411",x"150e07",x"311d0d",x"56361b",x"3d2310",x"2f1b0c",x"371f0e",x"39200f",x"3a2310",x"1d1208",x"361f0f",x"402511",x"432713",x"150e07",x"525252",x"525252",x"333333",x"323232",x"333333",x"303030",x"3e3e3e",x"323232",x"313131",x"313131",x"323232",x"313131",x"303030",x"2a2a2a",x"2f2f2f",x"313131",x"333333",x"333333",x"333333",x"323232",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"343434",x"323232",x"323232",x"323232",x"323232",x"343434",x"323232",x"333333",x"292929",x"2f2f2f",x"323232",x"333333",x"313131",x"323232",x"333333",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3628",x"4d3628",x"2a180b",x"381e0d",x"341d0d",x"1c1108",x"2d190b",x"2d190b",x"150e07",x"2f1b0c",x"381f0d",x"150e07",x"150e07",x"000000",x"000000",x"191008",x"191008",x"211409",x"2f1b0d",x"2d190b",x"331c0c",x"301a0b",x"351d0d",x"26160a",x"3d220f",x"3f3025",x"472c18",x"3c2314",x"3f2716",x"422816",x"3f2514",x"331e0e",x"946b4c",x"a37856",x"9b6f4f",x"986c4b",x"9a6d4c",x"9a6f4f",x"91684a",x"825c41",x"7e583f",x"a37756",x"8d6648",x"a37757",x"966b4c",x"95694a",x"926849",x"8f6546",x"95694a",x"946b4c",x"956c4c",x"92694a",x"906446",x"906647",x"8a6243",x"895f43",x"875c3f",x"805b3f",x"866043",x"936a4b",x"986d4d",x"845b3f",x"986c4b",x"8c6244",x"946849",x"8c6244",x"926647",x"81593d",x"885e40",x"926747",x"8b6143",x"835c40",x"7a573d",x"644732",x"4e3827",x"4e3827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200f",x"38200f",x"150e07",x"150e07",x"150e07",x"4e453d",x"4e453d",x"3b3026",x"4e2e18",x"4e2e18",x"2b190b",x"150e07",x"150e07",x"150e07",x"371e0d",x"391f0d",x"361e0d",x"331c0c",x"311b0b",x"351f0d",x"321c0c",x"3e230f",x"3f2410",x"3b210e",x"3e220f",x"1d1208",x"90694a",x"8b6244",x"8c6242",x"936747",x"986e4e",x"906545",x"8b6142",x"8f6546",x"936849",x"8c6244",x"966c4c",x"946b4d",x"8f6547",x"845d40",x"996f4f",x"855f44",x"966e4e",x"92684b",x"94694c",x"91694b",x"8c6244",x"9b7353",x"93694a",x"93694b",x"8f6648",x"855f42",x"986d4c",x"946a4b",x"8d6547",x"976d4d",x"8d6445",x"8c6345",x"8a6345",x"825b3f",x"7d573c",x"7b553a",x"66462f",x"422e1e",x"453020",x"453020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"483020",x"483020",x"442611",x"351c0c",x"3f2410",x"381f0d",x"381f0e",x"3c220f",x"432712",x"442812",x"3e220f",x"3c210f",x"4a2812",x"2f1b0c",x"2f1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"311d0d",x"331a0b",x"513524",x"2f1c0f",x"362e26",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"28180c",x"32271e",x"32271e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d3d3d",x"3b3b3b",x"3d3d3d",x"383838",x"333333",x"343434",x"393939",x"434343",x"595959",x"696969",x"474747",x"333333",x"323232",x"323232",x"323232",x"323130",x"333333",x"343434",x"373737",x"3b3b3b",x"323232",x"333333",x"343434",x"444444",x"3a3a3a",x"3f3f3f",x"3b3b3b",x"3d3d3d",x"404040",x"414141",x"3d3d3d",x"373737",x"3b3b3b",x"3b3b3b",x"3a3a3a",x"353535",x"3f3f3f",x"464646",x"3e3e3e",x"454545",x"323232",x"272727",x"2b2b2b",x"1f1f1f",x"2f2f2f",x"323232",x"323232",x"44423f",x"3c3a39",x"343433",x"362f2d",x"414141",x"414141",x"404040",x"454545",x"3f3f3f",x"333333",x"333333",x"323232",x"313131",x"313131",x"2e2e2e",x"333333",x"313131",x"313131",x"323232",x"323232",x"323232",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"333333",x"333333",x"313131",x"313131",x"333333",x"4b4b4b",x"484848",x"484848",x"4c4c4c",x"4a4a4a",x"434343",x"423f3c",x"433f3c",x"585756",x"575757",x"333333",x"313131",x"323232",x"333434",x"2f3030",x"2e2e2e",x"323232",x"323232",x"333333",x"202020",x"2f2f2f",x"444444",x"545454",x"313131",x"434343",x"525252",x"323232",x"323232",x"313131",x"313131",x"313131",x"343434",x"2d2d2d",x"323232",x"323232",x"333333",x"313131",x"323232",x"323232",x"313131",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"403126",x"403126",x"3b210f",x"3d220f",x"3a200e",x"150e07",x"321c0d",x"2e190b",x"1d1108",x"341e0d",x"150e07",x"3d220f",x"231509",x"26160a",x"26160a",x"323232",x"333333",x"313131",x"323232",x"323232",x"323232",x"333333",x"333333",x"2f2f2f",x"313131",x"303030",x"2f2f2f",x"2f2f2f",x"303030",x"323232",x"333333",x"323232",x"323232",x"323232",x"333333",x"313131",x"313131",x"323232",x"313131",x"323232",x"323232",x"333333",x"313131",x"313131",x"343434",x"303030",x"373838",x"2f2f2f",x"343434",x"32302f",x"313131",x"333333",x"444342",x"45413e",x"45413e",x"343230",x"302f2e",x"302f2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513d30",x"513d30",x"4a2b13",x"29180b",x"23150a",x"3c2311",x"391f0e",x"150e07",x"2d1b0d",x"37200f",x"180f08",x"3b2311",x"38210f",x"3c2210",x"563319",x"38200f",x"39200f",x"311b0c",x"3c2310",x"150e07",x"2f1b0c",x"3a210f",x"412611",x"4f2e16",x"150e07",x"525252",x"525252",x"454545",x"313131",x"323232",x"323232",x"323232",x"343434",x"343434",x"2f2f2f",x"353535",x"323232",x"2d2d2d",x"2d2d2d",x"2e2e2e",x"313131",x"323232",x"2e2e2e",x"313131",x"303030",x"313131",x"313131",x"303030",x"323232",x"313131",x"323232",x"323232",x"323232",x"333232",x"313131",x"323232",x"303030",x"353535",x"2f2f2f",x"303030",x"2a2a2a",x"333333",x"333333",x"313131",x"303030",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3628",x"4a3628",x"1e1208",x"3b210e",x"361e0d",x"311c0d",x"321c0c",x"311b0b",x"26160a",x"341e0d",x"371f0d",x"150e07",x"150e07",x"000000",x"000000",x"191008",x"191008",x"201309",x"2b180b",x"2d190b",x"311b0c",x"2e190b",x"341d0d",x"25150a",x"3f2411",x"443226",x"4a2c18",x"422816",x"3e2615",x"422715",x"3e2514",x"28180c",x"916748",x"966d4f",x"956a49",x"966a4b",x"9c6f50",x"a07554",x"886146",x"93694c",x"734f37",x"875f44",x"91684a",x"a47957",x"996f4f",x"986d4d",x"835b3f",x"956948",x"976b4b",x"966c4d",x"9a6f4e",x"9d7151",x"976b4c",x"93694a",x"95694b",x"8a6142",x"775239",x"926748",x"8b6244",x"956b4b",x"93694b",x"855b3e",x"8e6444",x"926647",x"946949",x"9a6e4e",x"906546",x"875d3f",x"895f41",x"8c6445",x"8a6042",x"7f593e",x"77553b",x"664a33",x"4e3827",x"4e3827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a2110",x"3a2110",x"150e07",x"150e07",x"150e07",x"4c4239",x"4c4239",x"3e342c",x"4f331f",x"4f331f",x"371f0e",x"150e07",x"150e07",x"150e07",x"41240f",x"3b200e",x"371e0d",x"3b210f",x"371e0d",x"3a210f",x"351e0d",x"351d0c",x"3f2410",x"3c210f",x"3b200e",x"1f1209",x"93694a",x"805a3f",x"885e43",x"8c6243",x"9a6d4d",x"865d41",x"8a5f41",x"8a6143",x"7e583c",x"835d40",x"866042",x"956c4e",x"855d40",x"946b4b",x"91694b",x"946c4c",x"986e4e",x"916749",x"936a4b",x"a07453",x"896043",x"a07757",x"94694a",x"93684a",x"976c4c",x"845d40",x"835d41",x"956c4c",x"875f43",x"946a4c",x"896144",x"8b6244",x"886144",x"7b563b",x"7c583c",x"7b563b",x"694931",x"493323",x"4a3423",x"4a3423",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452b1c",x"452b1c",x"442510",x"351d0c",x"3f2410",x"381f0e",x"38200e",x"3d220f",x"412612",x"3a210f",x"3f2310",x"3c210f",x"4c2c14",x"331d0d",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"311d0d",x"361d0d",x"533624",x"2f1d11",x"352d25",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"150e07",x"311d0d",x"29180c",x"2e261f",x"2e261f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"3b3b3b",x"3c3c3c",x"323232",x"323232",x"343434",x"323232",x"333333",x"313131",x"2f2f2f",x"2f2f2f",x"323232",x"313131",x"333333",x"323232",x"333333",x"333333",x"343434",x"313131",x"393939",x"3b3b3b",x"323232",x"333333",x"454545",x"3e3e3e",x"3e3f3f",x"3b3b3b",x"3f3f3f",x"3c3c3c",x"3c3d3d",x"3b3b3b",x"3c3c3c",x"3e3e3e",x"383838",x"3c3c3c",x"3b3b3b",x"363636",x"434343",x"454545",x"414141",x"4f4f4f",x"3d3d3d",x"323232",x"2d2d2d",x"2f2f2f",x"323232",x"333333",x"323232",x"323232",x"3e3e3e",x"484848",x"3b3b3b",x"373737",x"404040",x"313131",x"323232",x"353535",x"323232",x"323232",x"313131",x"313131",x"2e2e2e",x"333333",x"313131",x"313131",x"313131",x"313131",x"373737",x"393939",x"333333",x"323232",x"313131",x"333333",x"323232",x"333333",x"323232",x"333333",x"4a4a4a",x"4a4a4a",x"3f3f3f",x"373737",x"383838",x"363636",x"343434",x"323232",x"313131",x"303030",x"2a2a2a",x"2c2c2c",x"333333",x"313131",x"323232",x"333434",x"2f3030",x"2e2e2e",x"333333",x"313131",x"414141",x"414141",x"464646",x"434343",x"393939",x"4b4b4b",x"484848",x"474747",x"313131",x"313131",x"333333",x"323232",x"313131",x"343434",x"323232",x"323232",x"323232",x"333333",x"2f2f2f",x"2e2e2e",x"2d2d2d",x"313131",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3b3129",x"3b3129",x"381f0d",x"351e0d",x"361e0d",x"150e07",x"381f0e",x"341d0d",x"201308",x"150e07",x"2e1a0b",x"3f2310",x"27160a",x"26160a",x"26160a",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"323232",x"313131",x"333333",x"333333",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"303030",x"313131",x"313131",x"323232",x"353535",x"323232",x"323232",x"323232",x"343434",x"313131",x"323232",x"2d2d2d",x"303030",x"333333",x"333333",x"333333",x"323131",x"313131",x"323232",x"3f3f3f",x"555554",x"504d4a",x"413e3b",x"31302f",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d382b",x"4d382b",x"4e2c14",x"29170a",x"28170a",x"3b2210",x"231409",x"150e07",x"39210f",x"3a2210",x"150e07",x"150e07",x"2a180b",x"39200f",x"4d2c14",x"412511",x"38200f",x"311b0c",x"402612",x"150e07",x"2a180b",x"3a2210",x"3f2411",x"512f17",x"150e07",x"333333",x"333333",x"323232",x"303030",x"333333",x"323232",x"313131",x"333333",x"313131",x"313131",x"333333",x"2d2d2d",x"323232",x"303030",x"313131",x"323232",x"323232",x"323232",x"323232",x"333333",x"313131",x"323232",x"323232",x"333333",x"343434",x"323232",x"323232",x"323232",x"313131",x"333333",x"343434",x"303030",x"2d2d2d",x"282828",x"1f1f1f",x"2f2f2f",x"313131",x"333333",x"323232",x"303030",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513929",x"513929",x"26160a",x"3b210f",x"2f1a0b",x"2f1a0c",x"331c0c",x"341d0c",x"26170a",x"301b0c",x"39200e",x"150e07",x"150e07",x"000000",x"000000",x"191008",x"191008",x"201309",x"2b180b",x"2b180a",x"301a0b",x"2f1a0b",x"331c0c",x"231409",x"412511",x"402f24",x"482b18",x"402615",x"3b2414",x"3e2514",x"402614",x"311c0e",x"8e6549",x"9e7453",x"9a6f4f",x"94684a",x"976e4d",x"9d7253",x"956b4c",x"996e4e",x"946949",x"8f684b",x"94694a",x"a37857",x"946a4a",x"996d4e",x"926748",x"8a6143",x"956b4a",x"926748",x"906748",x"986c4c",x"956846",x"916545",x"906748",x"8c6244",x"825b3d",x"966a4a",x"966b4b",x"9d7050",x"906949",x"8a5f42",x"916645",x"926749",x"8c623f",x"916646",x"895e41",x"8a6142",x"8c6344",x"8c6244",x"8b6143",x"805a3f",x"755237",x"5f442e",x"4c3624",x"4c3624",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2311",x"3e2311",x"150e07",x"150e07",x"150e07",x"4c433a",x"4c433a",x"433930",x"52311c",x"52311c",x"2b180b",x"150e07",x"150e07",x"150e07",x"3e220e",x"3b210f",x"391f0d",x"3f2410",x"361d0d",x"371e0d",x"3c230f",x"331c0c",x"3b200e",x"3c210f",x"3c200e",x"211409",x"724e36",x"8d6345",x"855d40",x"875d41",x"9a6f4e",x"855c41",x"8a6041",x"845c3f",x"865d3f",x"8e6445",x"8f6447",x"966d4f",x"8d6345",x"926a4c",x"916548",x"956d4d",x"996f4e",x"996f4f",x"996d4c",x"976f4e",x"8a6144",x"987051",x"956d4d",x"956b4b",x"8f6547",x"8d6446",x"8e6446",x"805b3f",x"93694b",x"865f42",x"7b5639",x"8b6141",x"7e593d",x"7f593d",x"825c3f",x"755138",x"6a4932",x"483221",x"493322",x"493322",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462b1a",x"462b1a",x"462712",x"361d0c",x"39200e",x"381f0e",x"3c220f",x"3e2310",x"3f2410",x"3d220f",x"3e2310",x"3c210f",x"4a2912",x"2e1a0b",x"2e1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381e0d",x"381e0d",x"533623",x"2b1a10",x"373028",x"150e07",x"150e07",x"150e07",x"150e07",x"231509",x"150e07",x"150e07",x"150e07",x"150e07",x"311c0d",x"2b1a0d",x"332921",x"332921",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"404040",x"404040",x"414141",x"333333",x"322f2d",x"333333",x"333333",x"333232",x"2f2f2f",x"303030",x"2f2f2f",x"323232",x"323232",x"313131",x"323232",x"333333",x"303031",x"303131",x"373737",x"3a3a3a",x"3e3e3e",x"454545",x"444444",x"3f3f3f",x"3c3c3c",x"3b3b3b",x"3c3c3c",x"3c3c3c",x"3b3b3b",x"373737",x"393939",x"373737",x"3b3b3b",x"3c3c3c",x"3a3a3a",x"3a3a3a",x"3a3a3a",x"3c3c3c",x"3f3f3f",x"404040",x"444444",x"444444",x"424242",x"454545",x"505050",x"4c4c4c",x"4e4e4e",x"4e4e4e",x"464646",x"434343",x"414141",x"3b3b3b",x"363636",x"3b3b3b",x"414141",x"4e4e4e",x"4a4a4a",x"545454",x"4e4e4e",x"505050",x"535353",x"505050",x"545454",x"4c4c4c",x"4e4e4e",x"494949",x"444444",x"4c4c4c",x"424242",x"444444",x"4a4a4a",x"4c4c4c",x"505050",x"4f4f4f",x"404040",x"454545",x"3b3b3b",x"3a3a3a",x"343434",x"333333",x"383838",x"393939",x"3d3d3d",x"414141",x"484848",x"4a4a4a",x"4b4b4b",x"505050",x"4f4f4f",x"494949",x"525252",x"535353",x"505050",x"4f4f4f",x"505050",x"4a4a4a",x"424242",x"3e3e3e",x"353535",x"333333",x"323232",x"2f2f2f",x"333333",x"333333",x"333333",x"3d3d3d",x"383838",x"3c3c3c",x"3c3c3c",x"313131",x"343434",x"343434",x"343434",x"313131",x"313131",x"323232",x"323232",x"323232",x"373737",x"414141",x"282828",x"262626",x"262626",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"463428",x"463428",x"3a200e",x"321c0d",x"331c0c",x"361e0e",x"3b210f",x"3b200e",x"1a1008",x"29180b",x"351d0d",x"412410",x"251509",x"231509",x"231509",x"323232",x"333333",x"313131",x"313131",x"333333",x"313131",x"323232",x"333333",x"323232",x"313131",x"323232",x"333333",x"313131",x"303030",x"313131",x"343434",x"333333",x"2b221b",x"323232",x"343333",x"4d4742",x"504a44",x"343333",x"353535",x"44413d",x"575049",x"333232",x"363636",x"313131",x"3c3a38",x"4d4843",x"5e564f",x"46423f",x"313131",x"333333",x"2f2f2f",x"484848",x"575757",x"4a4a4a",x"434342",x"3d3d3c",x"2f2f2f",x"2f2f2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50392b",x"50392b",x"4d2c15",x"2a180b",x"29180b",x"3d2310",x"331d0c",x"351f0e",x"442713",x"402612",x"1c1108",x"331e0e",x"37200f",x"3d2210",x"4d2c15",x"3a210f",x"331d0d",x"27160a",x"432813",x"150e07",x"1c1108",x"331d0d",x"3a210f",x"4f2f16",x"150e07",x"474646",x"474646",x"313131",x"313131",x"303030",x"313131",x"323232",x"2c2c2c",x"343434",x"313131",x"333333",x"333333",x"3b3b3b",x"3c3c3c",x"3a3b3b",x"383838",x"333333",x"343434",x"323232",x"333434",x"313131",x"323232",x"333333",x"313131",x"333333",x"313131",x"323232",x"333333",x"323232",x"313131",x"313131",x"303030",x"2e2e2e",x"303030",x"313131",x"323232",x"313131",x"333333",x"333333",x"323232",x"343333",x"343333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3729",x"4e3729",x"27160a",x"3b210f",x"2e190b",x"26160a",x"311b0b",x"351d0d",x"25160a",x"231409",x"371e0d",x"150e07",x"150e07",x"000000",x"000000",x"190f08",x"190f08",x"1f1208",x"29180b",x"2a180a",x"301a0b",x"2e190b",x"341d0d",x"211409",x"422511",x"433429",x"4b2c18",x"412815",x"3d2414",x"3d2313",x"3c2414",x"2f1c0e",x"845d41",x"9a7151",x"966b4c",x"996e4f",x"a47958",x"a37756",x"986d4e",x"956c4d",x"9a6f50",x"9a6f4e",x"8d6445",x"a87c59",x"976d4e",x"886145",x"916647",x"845c3f",x"976e4e",x"956849",x"9b6f4f",x"986d4e",x"8d6342",x"8a603f",x"956a4b",x"986c4c",x"8b6143",x"976b4b",x"976c4c",x"986c4c",x"a17453",x"8c6143",x"8d6243",x"956a47",x"8a603f",x"916645",x"875e40",x"885f41",x"81573b",x"8b6244",x"896043",x"815b41",x"6f4e35",x"5f422d",x"4e3726",x"4e3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"361f0e",x"361f0e",x"150e07",x"150e07",x"150e07",x"544a40",x"544a40",x"443a31",x"462a15",x"462a15",x"2c190b",x"150e07",x"150e07",x"150e07",x"391e0c",x"3c220f",x"381f0d",x"3e230f",x"311a0b",x"391f0e",x"412611",x"371f0d",x"3b210e",x"361e0d",x"3c210e",x"1c1108",x"7f573e",x"966a4b",x"885f42",x"896042",x"966a4a",x"936a4a",x"714c35",x"916648",x"8a6042",x"8f6547",x"93694b",x"a27855",x"916748",x"916748",x"8a6144",x"8b6447",x"986e4e",x"926849",x"916749",x"9a704f",x"906446",x"a37856",x"9c7051",x"966b4c",x"8a6142",x"8f6647",x"976d4d",x"8d6546",x"8e6446",x"875e3f",x"795437",x"845c3d",x"815b40",x"805b3f",x"7e593e",x"7d573c",x"684931",x"4b3423",x"4a3423",x"4a3423",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432816",x"432816",x"452711",x"351c0c",x"3b210f",x"391f0e",x"381f0e",x"3f2410",x"442813",x"3b210e",x"422612",x"3a200e",x"482812",x"351f0e",x"351f0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"331a0b",x"331a0b",x"573722",x"27190f",x"352e26",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1209",x"150e07",x"150e07",x"150e07",x"191008",x"2d1a0c",x"25170c",x"312821",x"312821",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383838",x"414141",x"333333",x"322f2d",x"333333",x"333333",x"323232",x"2f2f2f",x"303030",x"000000",x"323232",x"323232",x"343434",x"343434",x"313131",x"505050",x"343434",x"393939",x"353535",x"3b3b3b",x"383838",x"393939",x"3b3b3b",x"3a3a3a",x"424242",x"3e3e3e",x"3d3d3d",x"3b3b3b",x"3a3a3a",x"3d3d3d",x"383838",x"3b3b3b",x"3c3c3c",x"393939",x"3a3a3a",x"393939",x"393939",x"393939",x"424242",x"434343",x"434343",x"474747",x"434444",x"434444",x"434343",x"424242",x"424343",x"424242",x"404040",x"3d3d3d",x"3c3c3c",x"404040",x"353535",x"3c3c3c",x"363636",x"3c3c3c",x"444444",x"404040",x"444444",x"393939",x"2d2d2d",x"484949",x"444444",x"414141",x"393939",x"454545",x"434343",x"434343",x"424242",x"3e3e3e",x"3f3f3f",x"434343",x"3a3a3a",x"414141",x"343434",x"494949",x"323232",x"575757",x"323232",x"444444",x"343434",x"383838",x"3f3f3f",x"414141",x"414141",x"3c3c3c",x"404040",x"414141",x"444444",x"444444",x"414141",x"414141",x"3a3a3a",x"3d3d3d",x"424242",x"383838",x"252525",x"393939",x"3c3c3c",x"333333",x"343434",x"333333",x"353535",x"393939",x"363636",x"3d3d3d",x"393939",x"303030",x"323232",x"343434",x"3a3a3a",x"3a3a3a",x"454545",x"3b3938",x"333333",x"373737",x"3a3735",x"3f3f3f",x"3f3f3f",x"414141",x"272727",x"272727",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"413329",x"413329",x"3e230f",x"402410",x"3c210f",x"3f2511",x"3b210e",x"361e0d",x"1c1108",x"361e0d",x"371f0e",x"462813",x"251509",x"231509",x"231509",x"333333",x"313131",x"343434",x"313131",x"323232",x"343434",x"323232",x"323232",x"323232",x"313131",x"313131",x"313131",x"343434",x"313131",x"343434",x"323231",x"323232",x"3c3c3c",x"3a3a3a",x"4f4d4b",x"66605b",x"504a44",x"343434",x"4d4c4c",x"453e38",x"4c453d",x"4e4d4b",x"565656",x"454444",x"423f3c",x"504841",x"5e564e",x"373635",x"373635",x"333333",x"2f2f2f",x"484848",x"575757",x"4a4a4a",x"434342",x"3d3d3c",x"2f2f2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3728",x"4e3728",x"583218",x"29180a",x"25160a",x"371f0e",x"361e0d",x"3b2210",x"412612",x"3e2411",x"1c1108",x"3c2310",x"371f0e",x"402410",x"4d2c15",x"341d0d",x"39200e",x"150e07",x"371f0e",x"150e07",x"311b0c",x"150e07",x"39200f",x"482914",x"150e07",x"4e4e4e",x"515151",x"323232",x"333333",x"333333",x"323232",x"2f2f2f",x"1b1b1b",x"313131",x"313131",x"2e2e2e",x"393736",x"59514a",x"544e48",x"575049",x"323232",x"323232",x"333333",x"2b2a29",x"383736",x"443f3b",x"5f574f",x"686059",x"625a52",x"595046",x"5a5147",x"5f564f",x"5e564f",x"5e564e",x"5d554d",x"4d4743",x"343434",x"343434",x"303030",x"313131",x"323232",x"313131",x"333333",x"333333",x"323232",x"343333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533f31",x"533f31",x"251509",x"351d0d",x"150e07",x"351d0d",x"2a180a",x"2d190b",x"341e0d",x"150e07",x"341d0d",x"150e07",x"150e07",x"000000",x"000000",x"191008",x"191008",x"1f1208",x"2a180b",x"2d190b",x"2c180a",x"2e190b",x"321c0c",x"201309",x"3f2410",x"44342a",x"4d2e19",x"422816",x"3e2514",x"3b2313",x"3c2413",x"29180b",x"875f43",x"936a4b",x"966b4c",x"986c4c",x"a07555",x"a47957",x"9c6f4e",x"9d7050",x"986b4c",x"9c7050",x"845c3f",x"a47958",x"9b7252",x"936b4b",x"7f593d",x"8c6344",x"956b4b",x"976b4b",x"8e6345",x"986c48",x"966a47",x"946744",x"9c7150",x"a07353",x"8f6445",x"895f42",x"9d7150",x"9d7151",x"9b6f50",x"8e6345",x"956948",x"976a48",x"956947",x"8e6346",x"956848",x"895e40",x"835a3c",x"8e6546",x"865e41",x"805a3f",x"6f4e35",x"5d412c",x"4f3726",x"4f3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"371e0d",x"371e0d",x"150e07",x"150e07",x"150e07",x"574d43",x"574d43",x"40372d",x"482c18",x"482c18",x"2b180b",x"150e07",x"150e07",x"150e07",x"3c200d",x"381f0e",x"361d0c",x"402511",x"361e0d",x"3b210e",x"402511",x"3f2310",x"3d220f",x"422511",x"40230f",x"211309",x"7d573d",x"825b3f",x"845c40",x"8c6344",x"8b6043",x"936748",x"926849",x"8e6547",x"835b3e",x"906647",x"926748",x"9a7151",x"976d4d",x"906747",x"8c6347",x"946a4b",x"976c4d",x"8a6045",x"926749",x"946b4b",x"956a4a",x"9a7152",x"996f4f",x"996e4e",x"956a4a",x"855d40",x"896144",x"91684a",x"7f593f",x"875e3e",x"8c6241",x"825b3b",x"815c40",x"6c4a33",x"855d42",x"785338",x"6a4b34",x"483322",x"4a3423",x"4a3423",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432917",x"432917",x"442711",x"341c0b",x"3d220f",x"402310",x"3b210e",x"3f2411",x"402511",x"3c210f",x"3a200e",x"3b210e",x"4a2a13",x"301c0c",x"301c0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402510",x"402510",x"523420",x"24190f",x"362f27",x"150e07",x"150e07",x"150e07",x"150e07",x"28170b",x"150e07",x"150e07",x"150e07",x"1a1008",x"2f1a0b",x"28180d",x"322921",x"322921",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"333333",x"323232",x"2f2f2f",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"333333",x"323232",x"555555",x"323232",x"373737",x"363636",x"323232",x"373737",x"373737",x"393939",x"393939",x"3c3c3c",x"3c3c3c",x"3c3c3c",x"3a3a3a",x"393939",x"3a3a3a",x"3e3e3e",x"3c3c3c",x"393a3a",x"3c3c3c",x"3c3c3c",x"3c3c3c",x"343434",x"363636",x"383838",x"3a3a3a",x"393939",x"474747",x"424242",x"3a3b3b",x"353535",x"3b3c3c",x"424242",x"393939",x"414141",x"3b3b3b",x"3f3f3f",x"373737",x"343434",x"373737",x"474747",x"3f3f3f",x"3b3b3b",x"494949",x"434343",x"373737",x"444444",x"474747",x"3f3f3f",x"434343",x"3c3c3c",x"3a3a3a",x"424242",x"404040",x"424242",x"414141",x"404040",x"3d3d3d",x"3b3b3b",x"3e3e3e",x"3d3d3d",x"3e3e3e",x"313131",x"555555",x"333333",x"4d4d4d",x"353535",x"3a3a3a",x"404040",x"404040",x"3b3b3b",x"414141",x"444444",x"3d3d3d",x"3a3a3a",x"464646",x"484848",x"3e3e3e",x"404040",x"464646",x"3c3c3c",x"3d3d3d",x"2d2d2d",x"343434",x"424242",x"313131",x"353535",x"323232",x"3c3c3c",x"353535",x"3d3d3d",x"464646",x"444444",x"3a3a3a",x"3f3f3f",x"363636",x"4a4a4a",x"4c4c4c",x"454545",x"4d4d4d",x"535353",x"585351",x"545454",x"4a4a4a",x"4a4a4a",x"4f4f4f",x"3e3e3e",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"473427",x"473427",x"3c220f",x"351e0e",x"361e0d",x"321c0d",x"39200e",x"351d0d",x"1e1208",x"29180b",x"341d0d",x"432712",x"27160a",x"231409",x"231409",x"333333",x"343434",x"333333",x"303030",x"323232",x"323232",x"313131",x"313131",x"333333",x"333333",x"313131",x"313131",x"323232",x"313131",x"333333",x"333333",x"333333",x"313131",x"393939",x"4a4847",x"645f5b",x"4b4742",x"333333",x"3d3d3d",x"65615c",x"625e5c",x"4b4b4b",x"414140",x"353535",x"44403c",x"59534c",x"5e564e",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513828",x"513828",x"4f2e15",x"2a180b",x"24150a",x"3a200e",x"3b210f",x"39200f",x"422611",x"3b210f",x"150e07",x"351f0f",x"341d0c",x"3f2310",x"482912",x"361f0d",x"3e2310",x"150e07",x"2f1b0c",x"150e07",x"351d0d",x"150e07",x"371f0e",x"452813",x"150e07",x"150e07",x"565656",x"333333",x"313131",x"333333",x"2f2f2f",x"292929",x"2d2d2d",x"333333",x"323232",x"444444",x"595756",x"69635b",x"4d4741",x"655d56",x"313131",x"323232",x"2c2d2d",x"4d4d4d",x"4a4a4a",x"55514d",x"655e57",x"6c665f",x"6d665f",x"6f6761",x"6d6660",x"6d6660",x"655e58",x"645c55",x"635b53",x"4c4641",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3c2f",x"4e3c2f",x"27160a",x"351d0d",x"371f0d",x"351d0d",x"301b0c",x"29170a",x"361f0e",x"39210f",x"2e1a0c",x"150e07",x"150e07",x"000000",x"000000",x"1b1008",x"1b1008",x"221409",x"29170a",x"2d1a0b",x"2b170a",x"2d190b",x"351d0d",x"201309",x"3f2411",x"46392e",x"4c2e19",x"3f2715",x"3a2314",x"3a2313",x"3d2313",x"301c0e",x"835c41",x"9f7252",x"966b4b",x"9a6d4d",x"a27654",x"a47958",x"9e7251",x"9c7050",x"986b4c",x"996e4d",x"7b5337",x"a27856",x"9e7454",x"946b4c",x"946849",x"8f6445",x"8d6446",x"8f6546",x"966c4c",x"9a7150",x"8a603f",x"986d4c",x"9b6f4f",x"986c4d",x"916647",x"8f6343",x"986b4c",x"9a6f4f",x"a07452",x"906547",x"7e563b",x"8a5f42",x"926647",x"926748",x"896042",x"855b3d",x"8b6244",x"936848",x"8b6343",x"845c41",x"755137",x"593e2a",x"4d3625",x"4d3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b210e",x"3b210e",x"150e07",x"150e07",x"150e07",x"574e43",x"574e43",x"453a31",x"4f311e",x"4f311e",x"331d0d",x"150e07",x"150e07",x"150e07",x"42240f",x"3c220f",x"321b0b",x"3e2310",x"3a200d",x"3a200e",x"3b220f",x"402511",x"3f2310",x"371f0e",x"3f230f",x"1b1008",x"8d6546",x"674531",x"8b6044",x"845c3f",x"916646",x"865d40",x"946a4a",x"8a6144",x"865b3f",x"966949",x"936849",x"a27655",x"9a7051",x"946a4a",x"9a6f4f",x"8c6447",x"8f6749",x"886043",x"946a4a",x"8e6445",x"926747",x"9c7454",x"996e4e",x"9b7051",x"956949",x"835d3f",x"815c41",x"8e6547",x"714d36",x"90674a",x"765236",x"8a6245",x"815b3f",x"855e41",x"7e593d",x"714e33",x"6b4a32",x"463120",x"453020",x"453020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432817",x"432817",x"432511",x"351c0c",x"3c210f",x"381f0e",x"39200e",x"402410",x"432712",x"371f0d",x"3b200e",x"402310",x"452611",x"301c0c",x"301c0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c200d",x"3c200d",x"563723",x"28190f",x"3b332c",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"191008",x"1b1108",x"2e1c0f",x"362e26",x"362e26",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"333333",x"323232",x"2f2f2f",x"333333",x"333231",x"313131",x"3e3f3f",x"383939",x"333333",x"34302e",x"323232",x"323232",x"333333",x"323232",x"2b2b2b",x"3a3a3a",x"383838",x"353535",x"363636",x"353535",x"3d3d3d",x"3a3a3a",x"3e3e3e",x"3d3d3d",x"3b3b3b",x"3b3b3b",x"3c3c3c",x"393939",x"3b3b3b",x"3a3a3a",x"363636",x"393939",x"3c3c3c",x"3a3a3a",x"3e3e3e",x"3f3f3f",x"3e3e3e",x"3e3e3e",x"3e3e3e",x"484848",x"4f4f4f",x"545454",x"5b5b5b",x"5a5a5a",x"555555",x"515151",x"494949",x"434343",x"424242",x"3d3d3d",x"323232",x"303030",x"434343",x"4f4f4f",x"515151",x"515151",x"585858",x"4f4f4f",x"555555",x"555555",x"545454",x"505050",x"555555",x"4d4d4d",x"444444",x"464646",x"434343",x"4b4b4b",x"505050",x"575757",x"5c5c5c",x"5b5b5b",x"555555",x"4d4d4d",x"4c4c4c",x"353535",x"333333",x"3a3a3a",x"474747",x"3b3b3b",x"383838",x"3f3f3f",x"4b4b4b",x"4f4f4f",x"545454",x"575757",x"5c5c5c",x"5c5c5c",x"595959",x"5c5c5c",x"525252",x"5c5c5c",x"555555",x"525252",x"4a4a4a",x"3a3a3a",x"414141",x"353535",x"3b3b3b",x"2f2f2f",x"373737",x"373737",x"3d3d3d",x"4f4f4f",x"4c4c4c",x"505050",x"4a4a4a",x"474747",x"434343",x"434343",x"494949",x"474747",x"494949",x"4b4b4b",x"494949",x"484848",x"454545",x"5d5d5d",x"474747",x"474747",x"474747",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"392c22",x"392c22",x"3d220f",x"3a210f",x"301b0c",x"1b1108",x"351d0d",x"331d0d",x"150e07",x"29180b",x"331c0d",x"412511",x"28170a",x"211309",x"211309",x"323232",x"333333",x"313131",x"323232",x"323232",x"323232",x"343434",x"323232",x"303030",x"313131",x"333333",x"323232",x"323232",x"323232",x"333333",x"3d3d3d",x"464646",x"575757",x"5b5b5b",x"595959",x"5a5959",x"4e4e4e",x"494949",x"5a5a5a",x"5c5c5b",x"575756",x"515151",x"444444",x"484848",x"565656",x"575757",x"515151",x"373737",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523827",x"523827",x"533116",x"29180b",x"29180b",x"391f0e",x"361e0d",x"27160a",x"3d2411",x"361e0e",x"150e07",x"28170b",x"311b0c",x"402411",x"4c2c15",x"341d0d",x"3f2310",x"3c220f",x"341e0e",x"301d0d",x"331c0c",x"150e07",x"3a210f",x"4f2e17",x"150e07",x"150e07",x"5b5b5b",x"606060",x"575757",x"494949",x"202020",x"202020",x"343434",x"333333",x"323232",x"333333",x"48433f",x"635b52",x"4f4a44",x"66605a",x"303030",x"343434",x"323232",x"333333",x"333333",x"4a4541",x"625a52",x"605850",x"615a51",x"605850",x"615a52",x"5e564e",x"5b534a",x"615952",x"5e564e",x"494541",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503c2f",x"503c2f",x"25150a",x"39200f",x"381f0d",x"391f0e",x"321c0c",x"28170a",x"3a210f",x"3a210f",x"341d0d",x"150e07",x"150e07",x"000000",x"000000",x"1d1208",x"1d1208",x"231509",x"2a180b",x"2d190b",x"2a160a",x"301b0b",x"2c190b",x"1f1309",x"3a200e",x"45362c",x"462a17",x"3d2414",x"382213",x"382211",x"3c2313",x"28170b",x"7b553a",x"956c4c",x"9b6f4f",x"946a4a",x"a07655",x"9a704f",x"a37756",x"986d4c",x"966a4b",x"946a4b",x"8f6345",x"956a4c",x"9c7253",x"896145",x"8a6144",x"885e40",x"906647",x"966a4a",x"9c7150",x"9b6f4f",x"956c4c",x"946949",x"996d4e",x"9e7252",x"956a4b",x"926646",x"986c4c",x"a17555",x"a57958",x"906547",x"936847",x"926848",x"986c4c",x"946849",x"8c6143",x"8b6040",x"906646",x"936748",x"865d40",x"835b40",x"755239",x"5c412b",x"493322",x"493322",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c220f",x"3c220f",x"150e07",x"150e07",x"150e07",x"544b41",x"544b41",x"40352b",x"50301a",x"50301a",x"28170a",x"150e07",x"150e07",x"150e07",x"3e220e",x"402410",x"371e0d",x"3c220f",x"3a200e",x"3e220f",x"381f0e",x"422611",x"3e2310",x"3a210f",x"3d220f",x"1e1208",x"896144",x"875e41",x"77523a",x"8f6647",x"946949",x"885e41",x"956a4b",x"906548",x"80573b",x"906445",x"956949",x"976f4e",x"996f4d",x"936a4b",x"966d4f",x"946b4d",x"996f4f",x"8d6446",x"90674b",x"8d6245",x"9a6f4e",x"997051",x"8f6549",x"966b4c",x"95694a",x"855c3e",x"996d4d",x"845c41",x"835c41",x"996e4e",x"875f42",x"7d563b",x"78533b",x"876145",x"815b3f",x"765238",x"62452e",x"473221",x"483221",x"483221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462a18",x"462a18",x"41230f",x"351d0c",x"3c210f",x"391f0d",x"3c220f",x"3d230f",x"3d2310",x"3c220f",x"3c210e",x"422611",x"41240f",x"361f0e",x"361f0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381f0c",x"381f0c",x"563722",x"24180f",x"3a322a",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"28180c",x"2f1f14",x"433a31",x"433a31",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"313131",x"323232",x"323232",x"303030",x"353330",x"313131",x"3e3f3f",x"383939",x"333333",x"34302e",x"323232",x"343434",x"333333",x"333333",x"2f2f2f",x"333333",x"393939",x"343434",x"333333",x"424242",x"343434",x"424242",x"3b3b3b",x"404040",x"3e3e3e",x"3d3d3d",x"3b3b3b",x"3b3b3b",x"3a3a3a",x"393939",x"393939",x"383838",x"3a3a3a",x"383838",x"373737",x"393939",x"3f3f3f",x"494949",x"535353",x"606060",x"464544",x"4a4947",x"514e4b",x"5d5751",x"6c6660",x"6b6560",x"5f5c5a",x"3f3f3f",x"3d3d3d",x"333333",x"323232",x"2d2d2d",x"2e2e2e",x"59544f",x"57534d",x"5a5550",x"5c5854",x"595550",x"5c5854",x"5b5753",x"655e57",x"615b54",x"67605a",x"655f59",x"5f5a56",x"5c5955",x"595959",x"5d5955",x"58534e",x"5c5752",x"59544e",x"59534e",x"5d5751",x"4d4d4d",x"575757",x"515151",x"474747",x"393939",x"353535",x"323232",x"363636",x"333333",x"514c47",x"5c564f",x"5d564f",x"59534c",x"5e5751",x"615a54",x"615b55",x"645e58",x"645c55",x"605954",x"625c56",x"4a4540",x"383838",x"5b5b5b",x"4e4e4e",x"373737",x"353535",x"383838",x"343434",x"323232",x"313131",x"323232",x"5f5852",x"56514b",x"474645",x"373736",x"3a3a3a",x"4c4c4c",x"4d4d4d",x"4a4a4a",x"4d4d4d",x"3c342d",x"363636",x"57534f",x"5c5855",x"504e4d",x"4f4f4f",x"474747",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"442f21",x"442f21",x"3d220f",x"3a210f",x"2b180b",x"3a220f",x"351d0d",x"2f1b0c",x"29170a",x"2b180b",x"2d1a0b",x"422611",x"28170a",x"28170a",x"28170a",x"333333",x"313131",x"313131",x"343434",x"323232",x"323232",x"333333",x"343434",x"333333",x"303030",x"313131",x"333333",x"333333",x"313131",x"323232",x"343434",x"2f2f2f",x"2e2e2e",x"2a2a2a",x"363533",x"4b453f",x"47423e",x"313131",x"313131",x"4f4a45",x"514b46",x"323131",x"343434",x"343434",x"3f3d3a",x"524c46",x"5d564e",x"45413d",x"45413d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513726",x"513726",x"502e15",x"2a190b",x"29180b",x"3b200e",x"3b210f",x"351d0d",x"3a2210",x"241509",x"3e2411",x"37200f",x"2f1a0b",x"3c210f",x"502d15",x"381f0e",x"2e1b0c",x"3c220f",x"150e07",x"37210f",x"1c1108",x"331d0d",x"3c210f",x"4d2d16",x"150e07",x"150e07",x"606060",x"585858",x"575757",x"515151",x"343434",x"343434",x"323232",x"3f3f3f",x"3e3d3d",x"454545",x"545453",x"565453",x"555555",x"6e6d6d",x"3c3c3c",x"313131",x"494949",x"4d4d4d",x"535353",x"575756",x"5a5957",x"5e5c5b",x"5e5c5b",x"605f5d",x"5e5c5b",x"605e5d",x"585858",x"575757",x"4a4a4a",x"434242",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3a2d",x"4e3a2d",x"211409",x"3d230f",x"321c0d",x"201309",x"150e07",x"221409",x"150e07",x"2b190b",x"39200e",x"191008",x"191008",x"000000",x"000000",x"201309",x"201309",x"27170a",x"2a180a",x"2c180b",x"29170a",x"311b0c",x"321d0d",x"1d1108",x"3b210f",x"493a2f",x"412615",x"432917",x"3b2213",x"392213",x"361f10",x"321d0e",x"8d6446",x"986d4f",x"684732",x"9a6e4d",x"a17453",x"9f7352",x"a17655",x"996f4f",x"92684a",x"996e4e",x"8b6245",x"986f4e",x"9d7251",x"92684b",x"956b4a",x"785037",x"946747",x"916646",x"996f4f",x"875d41",x"9b6f4e",x"855f43",x"946a4b",x"986e4e",x"93684a",x"956849",x"9a6d4c",x"a27654",x"a67957",x"926647",x"966948",x"986b4a",x"986c4b",x"966a49",x"8f6446",x"906444",x"936848",x"936848",x"825b3f",x"835c40",x"6f4c35",x"553b27",x"4b3523",x"4b3523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2411",x"3f2411",x"150e07",x"150e07",x"150e07",x"4f463c",x"4f463c",x"3c322a",x"4f2e17",x"4f2e17",x"2a180b",x"150e07",x"150e07",x"150e07",x"3a1f0d",x"412511",x"3d2210",x"432712",x"3b200e",x"3b200e",x"3e2310",x"422611",x"402410",x"3f2410",x"38200e",x"1d1108",x"8b6144",x"845b3f",x"926749",x"956949",x"8e6445",x"80573e",x"94684a",x"8e6446",x"885f41",x"926747",x"976b4b",x"94694a",x"916647",x"986f4f",x"8e6748",x"997050",x"9a6f51",x"94684a",x"9b7050",x"8c6243",x"896246",x"966d4d",x"90674a",x"91684a",x"916949",x"8b6143",x"845d3f",x"815a3e",x"896144",x"865e40",x"875f42",x"78533a",x"916a4b",x"79553c",x"7a553a",x"755138",x"6b4a32",x"4c3625",x"4b3524",x"4b3524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2e1d",x"4a2e1d",x"41230f",x"361e0d",x"3a200e",x"3a200e",x"3c210f",x"412511",x"3e2310",x"3c220f",x"3f230f",x"3c210f",x"492812",x"341e0e",x"341e0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b200c",x"3b200c",x"583620",x"2c1d11",x"393129",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"150e07",x"150e07",x"150e07",x"170f07",x"2d1a0d",x"312016",x"453c33",x"453c33",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"363636",x"363636",x"333333",x"303030",x"343434",x"313131",x"343434",x"3d3d3d",x"484848",x"565656",x"282828",x"232323",x"333333",x"323232",x"313131",x"303030",x"313131",x"353535",x"353535",x"3c3c3c",x"313131",x"4d4d4d",x"404040",x"414141",x"3b3b3b",x"3e3e3e",x"434343",x"414141",x"454545",x"3c3c3c",x"434343",x"3e3e3e",x"383838",x"313131",x"323232",x"343434",x"323232",x"414141",x"484848",x"5c5c5c",x"424242",x"3c3c3c",x"3f3f3f",x"43413f",x"484440",x"5d5751",x"313131",x"303030",x"323232",x"303030",x"323232",x"303031",x"303030",x"2f3030",x"323232",x"303030",x"323232",x"333333",x"343434",x"595550",x"5c5854",x"5b5753",x"655e57",x"615b54",x"67605a",x"655f59",x"635c57",x"5f5953",x"64605b",x"5d5955",x"58534e",x"5c5752",x"59544e",x"59534e",x"5d5751",x"4e4d4d",x"464545",x"474545",x"484848",x"515151",x"363636",x"333333",x"343434",x"363636",x"313131",x"313131",x"323232",x"323232",x"3b3b3b",x"615a54",x"615b55",x"645e58",x"645c55",x"605954",x"625c56",x"4a4540",x"383838",x"333333",x"3f3f3f",x"565656",x"484848",x"3b3b3b",x"3c3c3c",x"4b4b4b",x"3f3f3f",x"333333",x"2e2e2e",x"56514b",x"424141",x"3e3e3e",x"424141",x"3a3a3a",x"525252",x"555555",x"4d4d4d",x"343434",x"2e2e2e",x"57534f",x"5c5855",x"504e4d",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"453122",x"453122",x"3b210e",x"422712",x"301a0b",x"361f0e",x"150e07",x"2e1a0c",x"301b0c",x"150e07",x"29170a",x"3c210e",x"27160a",x"25150a",x"25150a",x"313030",x"313131",x"313131",x"343434",x"323232",x"323232",x"2f2f2f",x"323232",x"323232",x"323232",x"333333",x"323232",x"333333",x"323232",x"313131",x"2f2f2f",x"2d2d2d",x"242424",x"555555",x"4f4d4b",x"4d463f",x"3b3632",x"323232",x"3a3a3a",x"615b56",x"524f4c",x"3a3939",x"383838",x"343434",x"47433f",x"524c45",x"5b544c",x"353433",x"353433",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503828",x"503828",x"553117",x"27160a",x"2e1b0c",x"371e0d",x"3a200e",x"3c2210",x"331d0e",x"27170b",x"372110",x"3b2311",x"2f1a0c",x"3e220f",x"502d14",x"39200e",x"3f2411",x"321c0d",x"331d0e",x"150e07",x"341d0d",x"3a210f",x"3d220f",x"4c2d16",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"343434",x"343434",x"323232",x"3f3f3f",x"333333",x"343434",x"363636",x"2f2f2f",x"3a3a3a",x"333333",x"323232",x"393939",x"494949",x"4d4d4d",x"535353",x"575756",x"5a5957",x"5e5c5b",x"5e5c5b",x"605f5d",x"5e5c5b",x"605e5d",x"585858",x"575757",x"4a4a4a",x"434242",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"483629",x"483629",x"201309",x"422612",x"351e0e",x"331d0d",x"38200f",x"321c0c",x"251509",x"311c0c",x"371f0e",x"190f08",x"190f08",x"000000",x"000000",x"211409",x"211409",x"26160a",x"2a180a",x"2b180a",x"2c180a",x"2d190b",x"2e1b0c",x"1b1008",x"3a200f",x"4a3a2f",x"452a17",x"3d2413",x"3b2211",x"362012",x"372011",x"2a190c",x"896144",x"936a4b",x"876144",x"7a553d",x"9f7252",x"9f7251",x"a17555",x"966b4d",x"966c4d",x"976d4d",x"8e6245",x"9e7454",x"90694b",x"926849",x"976e4f",x"865c3e",x"8f6444",x"8a6143",x"9e7250",x"916444",x"936849",x"906749",x"946b4c",x"976c4c",x"966a4b",x"966a4b",x"976a4b",x"a67a58",x"9c7050",x"926646",x"956948",x"976a4b",x"966a4b",x"8e6344",x"926646",x"8f6444",x"8f6343",x"966a4a",x"795338",x"8a6245",x"6a4933",x"593e2b",x"4b3524",x"4b3524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"361f0e",x"361f0e",x"150e07",x"150e07",x"150e07",x"4c433a",x"4c433a",x"40362d",x"51311b",x"51311b",x"321c0d",x"150e07",x"150e07",x"150e07",x"3a1f0d",x"432712",x"432612",x"432712",x"381f0d",x"3f2310",x"3d220f",x"3f2411",x"3e2310",x"442611",x"38200e",x"1c1108",x"8b6447",x"8d6244",x"886042",x"926849",x"8f6447",x"8b6143",x"8d6345",x"916648",x"8e6445",x"886041",x"986e4e",x"9b7151",x"916647",x"966d4e",x"8f6547",x"956b4b",x"9c7352",x"92694b",x"9d7453",x"8e6445",x"986e4e",x"8d6649",x"966c4e",x"986d4c",x"8f6647",x"7f563b",x"875f42",x"845c3f",x"855c40",x"865e41",x"886043",x"855e42",x"8f6749",x"8d6447",x"7f5a3f",x"7c573d",x"6c4c34",x"4e3725",x"4b3524",x"4b3524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c3322",x"4c3322",x"442611",x"381f0e",x"331c0c",x"361d0c",x"3b200e",x"3e2310",x"3f2410",x"402410",x"3b200e",x"3b200e",x"4a2a13",x"361f0f",x"361f0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c210e",x"3c210e",x"54351f",x"2c1d11",x"3b332b",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1309",x"150e07",x"150e07",x"150e07",x"1b1008",x"2a180c",x"2c1f16",x"4a4037",x"4a4037",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494949",x"494949",x"474747",x"414141",x"3a3a3a",x"404040",x"494949",x"4d4d4d",x"525252",x"535353",x"282828",x"2e2e2e",x"2e2e2e",x"323232",x"333333",x"353535",x"383838",x"383838",x"3b3b3b",x"434343",x"313131",x"4f4f4f",x"333333",x"434343",x"3e3e3e",x"434343",x"474747",x"4b4b4b",x"535353",x"585858",x"595959",x"4e4e4e",x"464646",x"404040",x"404040",x"434343",x"4b4b4b",x"4e4e4e",x"555555",x"383838",x"3f3f3f",x"3c3c3c",x"3d3c3c",x"000000",x"484848",x"313131",x"323232",x"313131",x"333333",x"323232",x"333333",x"414141",x"424242",x"424242",x"474747",x"464646",x"353535",x"2e2f2f",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"64605b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"464545",x"454444",x"373737",x"333333",x"4a4a4a",x"373737",x"333333",x"323232",x"424242",x"323232",x"606060",x"575757",x"444444",x"444444",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"313131",x"313131",x"333333",x"474747",x"4a4a4a",x"4c4c4c",x"585858",x"484848",x"2e2e2e",x"2d2d2d",x"000000",x"000000",x"403f3f",x"444343",x"464646",x"5c5854",x"67605b",x"4a4948",x"3f3e3e",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"412d20",x"412d20",x"381e0d",x"39200e",x"371e0d",x"39200f",x"2f1a0b",x"2d190b",x"331d0d",x"150e07",x"341d0d",x"3a1f0d",x"25150a",x"25150a",x"25150a",x"323232",x"313131",x"313131",x"313131",x"313131",x"323232",x"313131",x"333333",x"313131",x"303030",x"313131",x"323232",x"333333",x"343434",x"313131",x"2a2a2a",x"1b1b1b",x"282828",x"313131",x"53504d",x"59544e",x"373431",x"303030",x"3d3d3d",x"68625d",x"585654",x"464545",x"363636",x"343333",x"4c4743",x"5b544d",x"565049",x"303030",x"303030",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f3728",x"4f3728",x"532f16",x"27160a",x"2d1a0b",x"341e0d",x"361e0d",x"3a210f",x"3d2310",x"2e1a0c",x"341e0e",x"150e07",x"331d0d",x"381e0d",x"492812",x"3c220f",x"3f2310",x"38200e",x"3f2411",x"150e07",x"2e190b",x"3b220f",x"452813",x"462812",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"313131",x"343434",x"313131",x"323232",x"313131",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a382b",x"4a382b",x"201309",x"3f2411",x"3d2311",x"321c0c",x"381f0e",x"3c220f",x"2c190b",x"341d0d",x"3e2310",x"150e07",x"150e07",x"000000",x"000000",x"211309",x"211309",x"28170b",x"271509",x"251409",x"2a170a",x"271609",x"221309",x"1b1008",x"3a210f",x"4f3b2e",x"4a2c18",x"3f2715",x"422715",x"402514",x"382012",x"2a190c",x"896244",x"9b7051",x"8f6749",x"8b6345",x"a37957",x"936849",x"996f51",x"996d4e",x"90674a",x"9a7050",x"946849",x"9d7453",x"976c4d",x"8c6346",x"946a4a",x"6c432a",x"926647",x"926746",x"976b4b",x"926646",x"926648",x"956b4c",x"92694a",x"95694a",x"936747",x"966949",x"976c4d",x"a47856",x"986d4b",x"956848",x"926748",x"906445",x"926747",x"7f573d",x"8b6243",x"946848",x"785239",x"916646",x"8e6546",x"805a3e",x"7b583d",x"5c402c",x"4c3525",x"4c3525",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2410",x"3e2410",x"150e07",x"150e07",x"150e07",x"4d443b",x"4d443b",x"42382f",x"4f321f",x"4f321f",x"341d0d",x"150e07",x"150e07",x"150e07",x"422510",x"452814",x"412612",x"432712",x"3e230f",x"3d220f",x"3c210f",x"402510",x"412511",x"361e0d",x"412410",x"1d1108",x"815a3e",x"8c6244",x"8b6143",x"946a4a",x"95694a",x"926647",x"916646",x"926749",x"885f41",x"8e6445",x"92684a",x"91694b",x"8c6244",x"92694a",x"966b4c",x"8d6346",x"8f664a",x"966d4e",x"936a4c",x"906648",x"956a4a",x"966d4d",x"a27655",x"9b7150",x"94694a",x"643c14",x"906648",x"885f41",x"8a6144",x"7f593c",x"8d6446",x"8a6244",x"865f44",x"866042",x"815a3f",x"79553a",x"6a4a33",x"4b3525",x"4c3626",x"4c3626",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513727",x"513727",x"402310",x"3b210f",x"321c0c",x"361e0d",x"3b210e",x"3f2410",x"3c210f",x"3f2310",x"3c2310",x"3f230f",x"472812",x"311c0d",x"311c0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422511",x"422511",x"4f311e",x"2e1e14",x"3d352d",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"180f07",x"26170d",x"2c1f16",x"4b4138",x"4b4138",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595959",x"595959",x"444444",x"474747",x"3c3c3c",x"484848",x"4e4e4e",x"525252",x"545454",x"5b5b5b",x"323131",x"313131",x"333333",x"313131",x"343434",x"363636",x"393939",x"3d3d3d",x"3d3d3d",x"3f3f3f",x"474747",x"444444",x"474747",x"434343",x"464646",x"4d4d4d",x"585858",x"505050",x"535252",x"5d5a56",x"494746",x"434343",x"4e4e4e",x"535353",x"4c4c4c",x"494949",x"4c4c4c",x"474747",x"313131",x"333333",x"3a3a3a",x"000000",x"000000",x"000000",x"484848",x"484848",x"595554",x"585858",x"484949",x"555555",x"545454",x"515151",x"505050",x"545454",x"525252",x"535353",x"5d5d5d",x"535353",x"373737",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"303030",x"343434",x"343434",x"3b3b3b",x"484848",x"515151",x"4c4c4c",x"3e3e3e",x"444444",x"404040",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"303030",x"656565",x"585858",x"4a4a4a",x"525252",x"585858",x"343434",x"2d2d2d",x"2e2e2e",x"000000",x"000000",x"000000",x"000000",x"4a4847",x"5c5854",x"67605b",x"575552",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3f2e23",x"3f2e23",x"331c0c",x"311a0b",x"2f1a0b",x"1c1108",x"351d0d",x"331c0c",x"150e07",x"28160a",x"321c0c",x"391e0d",x"27160a",x"251509",x"251509",x"333333",x"343434",x"323232",x"323232",x"333333",x"313131",x"313131",x"302e2c",x"323232",x"323232",x"2f2f2f",x"313131",x"2d2d2d",x"313131",x"323232",x"363636",x"2a2a2a",x"4e4e4e",x"555555",x"545352",x"555251",x"3e3d3c",x"353535",x"4c4c4c",x"545250",x"454545",x"3b3b3b",x"353535",x"353535",x"4d4c4b",x"4f4e4d",x"494949",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"373635",x"373636",x"585653",x"545454",x"363636",x"2f2f2f",x"323232",x"313131",x"343434",x"313131",x"333333",x"323232",x"323232",x"323232",x"323232",x"313131",x"313131",x"2f2f2f",x"383838",x"323232",x"503829",x"462711",x"28160a",x"2b180b",x"3e2310",x"311b0b",x"1c1108",x"331d0d",x"321c0d",x"150e07",x"24150a",x"321c0d",x"381f0d",x"4d2a13",x"3d220f",x"331b0b",x"331d0d",x"402511",x"150e07",x"2b170a",x"3b2310",x"3c210f",x"482813",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"32302f",x"333333",x"323232",x"323232",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"473427",x"473427",x"29180b",x"402410",x"38200e",x"301b0c",x"3b220f",x"3b210f",x"2b190b",x"351d0d",x"361e0d",x"150e07",x"150e07",x"000000",x"000000",x"22150b",x"22150b",x"27180c",x"231309",x"241308",x"281609",x"271609",x"29160a",x"180f08",x"371f0d",x"4f3c2e",x"4c2f19",x"412614",x"402614",x"3c2513",x"392212",x"321d0e",x"8c6345",x"8b6245",x"8e6446",x"986d4d",x"90684a",x"835c40",x"9c7152",x"9c7151",x"90684a",x"8d6649",x"956a4a",x"9c7052",x"936a4b",x"956a4a",x"80583e",x"875f41",x"82583d",x"996d4c",x"976c4d",x"8d6242",x"95694a",x"8f6649",x"8a6345",x"946849",x"95694a",x"916546",x"9d7150",x"9b6f4f",x"9f7351",x"966a4b",x"966a4a",x"946747",x"8d6143",x"916647",x"8d6242",x"906546",x"795239",x"946948",x"926848",x"865d41",x"7b563c",x"5f422d",x"4d3625",x"4d3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2411",x"3e2411",x"150e07",x"150e07",x"150e07",x"4b4238",x"4b4238",x"43372d",x"52321c",x"52321c",x"2a180b",x"150e07",x"150e07",x"150e07",x"40230f",x"452814",x"3e2310",x"3f2411",x"3c220f",x"3e230f",x"3f2410",x"3f2411",x"39200e",x"3d2310",x"412410",x"1b1108",x"886042",x"8e6546",x"8c6343",x"986c4b",x"946949",x"906646",x"976c4c",x"956b4c",x"895e41",x"986c4c",x"8d6344",x"94694a",x"7f573b",x"956b4b",x"9b7050",x"926849",x"9c7051",x"996e4f",x"936849",x"926749",x"996f4f",x"966b4c",x"997050",x"906748",x"986c4c",x"865e40",x"8a6244",x"896043",x"825c40",x"835c3e",x"865e41",x"916647",x"7f5b40",x"855e42",x"855e41",x"76533a",x"6a4a33",x"4a3424",x"493323",x"493323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422d22",x"422d22",x"452711",x"3d2310",x"351e0d",x"371e0d",x"381f0d",x"3c220f",x"3e230f",x"3f2410",x"472914",x"3f2410",x"4b2c14",x"321c0d",x"321c0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432712",x"432712",x"603e27",x"332115",x"3c332b",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1209",x"150e07",x"150e07",x"150e07",x"1e1208",x"21150c",x"312319",x"4c4238",x"4c4238",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"636363",x"636363",x"606060",x"545454",x"434343",x"505050",x"5c5c5c",x"545454",x"5f5f5f",x"616161",x"2a2a29",x"323232",x"303030",x"313131",x"3a3a3a",x"444444",x"4d4d4d",x"4e4e4e",x"555555",x"555555",x"535353",x"555555",x"545454",x"555555",x"585858",x"5a5a5a",x"484848",x"4c4c4c",x"4f4f4f",x"5d5a56",x"393939",x"494949",x"424242",x"5e5e5e",x"565656",x"515151",x"565656",x"313131",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"616161",x"616161",x"535353",x"4c4c4c",x"5c5c5c",x"5e5e5e",x"5d5d5d",x"5a5a5a",x"565656",x"505050",x"4e4e4e",x"4f4f4f",x"595959",x"4a4949",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"484848",x"484848",x"444444",x"636363",x"525252",x"575757",x"4e4e4e",x"575757",x"3c3c3c",x"323232",x"323232",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"606060",x"646361",x"59534d",x"605852",x"615d58",x"474645",x"393735",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a3427",x"4a3427",x"371e0d",x"361e0d",x"321b0b",x"341e0d",x"3d220f",x"351d0d",x"180f07",x"301b0c",x"351d0d",x"452712",x"26160a",x"241509",x"241509",x"343434",x"343434",x"343434",x"313131",x"313131",x"343434",x"333333",x"313131",x"313131",x"303030",x"343434",x"313131",x"353535",x"333333",x"292929",x"2c2c2c",x"242424",x"303030",x"404040",x"413d3a",x"4f4943",x"383633",x"333333",x"40403f",x"625c55",x"504d4a",x"3c3c3b",x"333333",x"313030",x"413d3a",x"544d47",x"5a534d",x"47433f",x"47433f",x"000000",x"000000",x"000000",x"000000",x"000000",x"373635",x"373636",x"585653",x"545454",x"363636",x"2f2f2f",x"323232",x"313131",x"343434",x"313131",x"333333",x"323232",x"323232",x"323232",x"323232",x"313131",x"313131",x"2f2f2f",x"383838",x"323232",x"2f1b0c",x"432511",x"261509",x"29170a",x"3c220f",x"361d0d",x"331c0c",x"381e0d",x"3a200f",x"150e07",x"2f1b0c",x"361f0e",x"391f0d",x"4f2c14",x"371f0d",x"31190b",x"331d0d",x"402511",x"150e07",x"301a0b",x"3d2310",x"3d220f",x"492a13",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"32302f",x"333333",x"323232",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463326",x"463326",x"2a180b",x"472914",x"39210f",x"361f0e",x"38200f",x"371f0e",x"2b190b",x"351d0d",x"361e0d",x"150e07",x"150e07",x"000000",x"000000",x"20140b",x"20140b",x"26170b",x"24150b",x"221208",x"28160a",x"241409",x"251409",x"170f07",x"341d0d",x"4b392c",x"4c2d19",x"422716",x"3f2514",x"3f2514",x"392213",x"29180b",x"63432f",x"875f44",x"885f41",x"986f4e",x"845c40",x"8d6345",x"966d4d",x"99704f",x"886044",x"896144",x"936848",x"9a704f",x"8f674b",x"896346",x"8e6446",x"926749",x"855c3e",x"966b4a",x"976c4b",x"926747",x"926749",x"986d4e",x"906647",x"7f573c",x"875f43",x"8b6145",x"996e4e",x"90694a",x"a17452",x"996e4c",x"95694b",x"976a4b",x"906545",x"8f6445",x"7e573a",x"845c3e",x"8e6345",x"956949",x"896043",x"8f6547",x"7e5a3e",x"60422e",x"4f3726",x"4f3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432712",x"432712",x"150e07",x"150e07",x"150e07",x"4e453c",x"4e453c",x"463b31",x"513017",x"513017",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"422410",x"3e2310",x"3f2310",x"432713",x"3a200e",x"371f0e",x"37200e",x"412510",x"3d220f",x"3f2410",x"432610",x"211409",x"926848",x"8d6344",x"9a6f4e",x"976a4a",x"956a4a",x"936847",x"94694a",x"916647",x"865b3f",x"966a4b",x"916546",x"996c4c",x"8d6242",x"91694a",x"9d7251",x"875f43",x"a17555",x"92684a",x"94694a",x"936849",x"986f50",x"986c4d",x"9c7352",x"8f6849",x"946949",x"896142",x"926849",x"8b6345",x"845c40",x"896043",x"845e41",x"8d6346",x"93694a",x"7c563c",x"7c573d",x"7c573c",x"694932",x"483221",x"493321",x"493321",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412f25",x"412f25",x"432611",x"3a210f",x"3d220f",x"341c0c",x"3b210e",x"341d0d",x"3d220f",x"3f2310",x"432712",x"412511",x"4e2d15",x"2b190b",x"2b190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2c1a0c",x"2e1b0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442712",x"442712",x"49301f",x"302117",x"3f372f",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"150e07",x"150e07",x"150e07",x"150e07",x"23140a",x"2b2017",x"4a4037",x"4a4037",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"625e5a",x"625e5a",x"625c58",x"5a5147",x"6a6561",x"706963",x"6f6a64",x"706a65",x"6e6963",x"6d6965",x"67625e",x"59544f",x"5f5852",x"6c655f",x"68645f",x"6e6964",x"6f6a65",x"6f6a66",x"6f6a65",x"736d68",x"706a63",x"6b6863",x"6e6965",x"6c6863",x"6c6863",x"565655",x"4d4d4d",x"484848",x"000000",x"000000",x"4c4c4c",x"4d4d4d",x"4f4f4f",x"595857",x"5f5953",x"494643",x"363636",x"353535",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"626262",x"4b4b4b",x"444444",x"474544",x"4e4c4a",x"54514f",x"424242",x"565656",x"535353",x"595551",x"58534f",x"504d4c",x"595959",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4a4a",x"4e4e4e",x"565655",x"54514e",x"494949",x"4b4b4b",x"5c5c5c",x"595959",x"414141",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"626161",x"646361",x"59534d",x"605852",x"615d58",x"53504d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"493528",x"493528",x"381f0d",x"3b210f",x"341c0c",x"3b210e",x"3c220f",x"3a200e",x"150e07",x"351f0f",x"3d2310",x"482a13",x"29170a",x"261509",x"261509",x"313131",x"333333",x"333333",x"313131",x"343434",x"333333",x"323232",x"313131",x"2f2f2f",x"353535",x"333333",x"313131",x"333333",x"333333",x"303030",x"2d2d2d",x"2c2926",x"2f2f2f",x"545454",x"5f5c59",x"565049",x"383735",x"383837",x"595858",x"6b655f",x"585554",x"4a4a4a",x"4b4b4b",x"353434",x"4c4843",x"5a534c",x"534d47",x"393837",x"393837",x"000000",x"000000",x"000000",x"000000",x"373635",x"373635",x"373635",x"5d5a58",x"565655",x"302f2e",x"313131",x"323232",x"323232",x"303030",x"343434",x"303030",x"343434",x"323232",x"323232",x"323232",x"333333",x"2f2f2f",x"2e2e2e",x"383838",x"333333",x"252525",x"482811",x"231409",x"29170a",x"391f0e",x"331c0c",x"412511",x"391f0d",x"3c210f",x"3c210f",x"2c1a0b",x"39210f",x"3d220f",x"4c2b14",x"371f0d",x"341c0c",x"2e190a",x"39200e",x"150e07",x"2e190b",x"3c220f",x"3c210f",x"442611",x"150e07",x"150e07",x"4f4f4f",x"3f3f3f",x"111111",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"2f2f2f",x"313131",x"333333",x"313131",x"323232",x"343434",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"303030",x"333333",x"323232",x"323232",x"323232",x"323232",x"2c2c2c",x"313131",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"433024",x"433024",x"29180b",x"3f2410",x"3d2411",x"311c0c",x"371f0e",x"341d0d",x"251509",x"341c0c",x"381f0e",x"150e07",x"150e07",x"000000",x"000000",x"20140b",x"20140b",x"25170b",x"25160b",x"23140a",x"29170a",x"241409",x"27160a",x"160e07",x"311c0d",x"4b3b2f",x"452915",x"442815",x"402514",x"412615",x"3b2313",x"341e0f",x"8d6446",x"845d41",x"8b6141",x"956b4b",x"956b4b",x"976b4b",x"9d7151",x"9d7454",x"906748",x"875f43",x"8d6548",x"896244",x"8d6649",x"90694a",x"9f7251",x"906648",x"845b3f",x"9c7050",x"9b6f4f",x"946848",x"8e6446",x"936a4a",x"8d6445",x"82593e",x"996e4e",x"8f6546",x"966b4b",x"9a6f4f",x"9d7150",x"9c704e",x"986c4b",x"8e6244",x"8d6345",x"8b6143",x"8f6445",x"8d6244",x"8d6345",x"946a49",x"895f41",x"885f44",x"6c4b35",x"634630",x"4f3726",x"4f3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a210f",x"3a210f",x"150e07",x"150e07",x"150e07",x"4b4238",x"4b4238",x"3f342b",x"4f301b",x"4f301b",x"351d0d",x"150e07",x"150e07",x"150e07",x"412410",x"422712",x"412511",x"442813",x"3a200e",x"3a210f",x"39200e",x"3f2411",x"3e2310",x"3f2310",x"412510",x"1c1108",x"8a6042",x"8d6344",x"936a4a",x"926748",x"9b6e4d",x"966a49",x"956a48",x"865b3f",x"885d40",x"9c7050",x"996c4c",x"93684a",x"8e6344",x"996d4d",x"9a6f4f",x"956848",x"946b4d",x"956a4b",x"9b6e4e",x"8c6345",x"956c4d",x"936949",x"926a4c",x"966d4d",x"976d4e",x"886042",x"896244",x"8f6849",x"8e6546",x"8a6243",x"835c3e",x"8b6144",x"8d6446",x"815a3e",x"825b3f",x"7d583c",x"6d4c35",x"483322",x"493322",x"493322",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3224",x"4a3224",x"482913",x"3f2410",x"371f0e",x"2b170a",x"3c220f",x"3b200e",x"3d220f",x"3d220f",x"402411",x"412511",x"502e16",x"301b0c",x"301b0c",x"000000",x"000000",x"000000",x"000000",x"351f0e",x"241409",x"2c1a0c",x"2e1b0c",x"1c1108",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f230f",x"3f230f",x"4d3323",x"2f2017",x"413931",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"150e07",x"150e07",x"150e07",x"1a1008",x"25150b",x"2e2016",x"453b31",x"453b31",x"000000",x"000000",x"5e4e42",x"4d2c15",x"482812",x"482812",x"482812",x"625e5a",x"625c58",x"5a5147",x"6a6561",x"706963",x"6f6a64",x"706a65",x"6e6963",x"6d6965",x"67625e",x"59544f",x"5f5852",x"6c655f",x"68645f",x"6e6964",x"746d67",x"6f6a66",x"6f6a65",x"736d68",x"706a63",x"6b6863",x"6e6965",x"6c6863",x"6c6863",x"4b2b14",x"452712",x"4d2d15",x"513017",x"523117",x"4b2b14",x"533117",x"4f4f4f",x"5c5a57",x"5f5953",x"605951",x"4e2d15",x"4c2c15",x"4f2d15",x"4a2a14",x"4f2e16",x"4c2c15",x"502e15",x"4a2a13",x"4a2a13",x"4a2a14",x"4f2e15",x"4c2d15",x"4b4947",x"53504d",x"54514f",x"5d5651",x"625c56",x"5e5955",x"625b54",x"58534f",x"565350",x"5b3a21",x"5f3c22",x"5f3e24",x"59381f",x"5d3a21",x"54341d",x"54341d",x"4e301a",x"52321c",x"4f2f19",x"53321c",x"4f301a",x"53331c",x"4b2c16",x"4f311c",x"4b2e18",x"4e301b",x"4a2c18",x"4c2f1a",x"4d2f19",x"55351e",x"51321c",x"515151",x"5a5958",x"54514e",x"4f4c49",x"565350",x"6a635d",x"5b5956",x"4c4c4c",x"563822",x"53351f",x"54361f",x"4e301c",x"4f331e",x"4e301b",x"51331d",x"4f311b",x"50321b",x"55341c",x"52331c",x"4e301a",x"50311c",x"50311b",x"51311b",x"512f18",x"52321c",x"56341c",x"5a371f",x"59361d",x"56341d",x"4f301a",x"6a4c33",x"6a4c33",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"403328",x"403328",x"3a200e",x"3c210f",x"341c0c",x"381f0e",x"3a210f",x"371f0d",x"412511",x"321d0d",x"39200e",x"452813",x"29170a",x"241409",x"241409",x"333333",x"343434",x"303030",x"313131",x"333333",x"323232",x"343434",x"313131",x"323232",x"313131",x"333333",x"313131",x"313131",x"313131",x"2e2e2e",x"323232",x"323232",x"3e3e3e",x"444444",x"5c5854",x"625d58",x"333231",x"333333",x"424241",x"67615a",x"4e4d4c",x"434343",x"393939",x"363534",x"4e4943",x"5e564f",x"3f3d3b",x"323232",x"313131",x"303030",x"5a5959",x"4a4846",x"393531",x"31302f",x"383533",x"383533",x"5e5c5b",x"575757",x"323232",x"303030",x"323232",x"323232",x"323232",x"313131",x"323232",x"313131",x"2f2f2f",x"333333",x"303030",x"343434",x"333333",x"454545",x"383837",x"323232",x"312f2d",x"4a2912",x"1c1108",x"29170a",x"3a200e",x"331c0c",x"361e0d",x"3d230f",x"402411",x"3a200e",x"29180b",x"371f0e",x"381f0e",x"472611",x"381e0d",x"381f0d",x"29170a",x"381f0e",x"150e07",x"301a0b",x"341d0e",x"371f0d",x"472812",x"150e07",x"4f4f4f",x"4f4f4f",x"3f3f3f",x"111111",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"2f2f2f",x"313131",x"333333",x"313131",x"323232",x"343434",x"333333",x"323232",x"333333",x"323232",x"323232",x"333333",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"303030",x"333333",x"323232",x"323232",x"323232",x"323232",x"2c2c2c",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422f23",x"422f23",x"2c190b",x"432712",x"38200f",x"331d0d",x"361f0e",x"311c0c",x"28160a",x"2f1a0b",x"351d0d",x"150e07",x"150e07",x"000000",x"000000",x"20140b",x"20140b",x"27180c",x"29190c",x"27180b",x"29180c",x"25170b",x"221309",x"160f07",x"3a2210",x"544032",x"452915",x"3b2314",x"3c2314",x"362012",x"331e10",x"28170b",x"906647",x"926748",x"8c6242",x"8f6749",x"9b704f",x"875e41",x"976e4d",x"9c7152",x"936849",x"896144",x"835b41",x"8c6548",x"896247",x"936a4c",x"9b6f4e",x"906648",x"916648",x"976d4d",x"966b4a",x"976c4b",x"8f6445",x"936849",x"956b4b",x"8b6042",x"8f6345",x"8b6144",x"885f41",x"956a4b",x"976b4a",x"956b4b",x"946a4a",x"8d6344",x"916647",x"896041",x"8a6143",x"865e42",x"8f6647",x"9a704f",x"8f6546",x"805a3f",x"7a573d",x"61452f",x"4e3626",x"4e3626",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a220f",x"3a220f",x"150e07",x"150e07",x"150e07",x"4f453c",x"4f453c",x"473a31",x"4d3120",x"4d3120",x"331d0d",x"150e07",x"150e07",x"150e07",x"442611",x"402511",x"432612",x"432712",x"3b210f",x"3b210f",x"3a210f",x"3f2411",x"3f2410",x"3d220f",x"422511",x"1d1108",x"8f6749",x"8b6243",x"956b4b",x"996c4c",x"896145",x"845b3e",x"95694a",x"845b3e",x"8a6042",x"9b6e4d",x"976a4b",x"976c4b",x"966a49",x"a07351",x"9b6f4e",x"966b4b",x"9d7051",x"9d7151",x"93684a",x"926749",x"956d4d",x"936849",x"976e4e",x"996f50",x"946b4c",x"8d6346",x"976d4c",x"8a6144",x"8c6446",x"8b6243",x"855d41",x"8d6446",x"8d6245",x"815a3d",x"815a3f",x"724f36",x"66472f",x"442f1f",x"453020",x"453020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a3527",x"4a3527",x"4b2a13",x"3b220f",x"3b210f",x"2e180a",x"39200e",x"3b200e",x"371e0d",x"3b210f",x"422611",x"432712",x"462812",x"331d0d",x"331d0d",x"000000",x"000000",x"000000",x"000000",x"3b2210",x"351f0e",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e230f",x"3e230f",x"4f3220",x"2b1e14",x"3f372e",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"150e07",x"150e07",x"150e07",x"170f07",x"29170a",x"2d1e13",x"433930",x"433930",x"000000",x"5e4e42",x"5e4e42",x"4d2c15",x"482812",x"482812",x"482812",x"442611",x"452711",x"452611",x"482811",x"492913",x"4a2a13",x"4a2a14",x"4a2913",x"4a2a13",x"482812",x"432510",x"482813",x"442511",x"4d2d15",x"4b2a13",x"4f2e15",x"4f2d15",x"4c2b14",x"4b2b14",x"4d2d15",x"4d2d15",x"4f2f17",x"513018",x"513017",x"4b2b14",x"452712",x"4d2d15",x"513017",x"523117",x"4b2b14",x"533117",x"4f2d15",x"4b2b13",x"482813",x"4d2c14",x"4e2d15",x"4c2c15",x"4f2d15",x"4a2a14",x"4f2e16",x"4c2c15",x"502e15",x"4a2a13",x"4a2a13",x"4a2a14",x"4f2e15",x"4c2d15",x"4d2c14",x"422410",x"452610",x"472711",x"4c2a13",x"936c4a",x"5c3a21",x"5d3d24",x"5b3a21",x"5b3a21",x"5f3c22",x"5f3e24",x"59381f",x"5d3a21",x"54341d",x"54341d",x"4e301a",x"52321c",x"4f2f19",x"53321c",x"4f301a",x"53331c",x"4b2c16",x"4f311c",x"4b2e18",x"4e301b",x"4a2c18",x"4c2f1a",x"4d2f19",x"55351e",x"51321c",x"5a3921",x"50321d",x"573820",x"58371f",x"523520",x"54361f",x"573720",x"50321d",x"563822",x"53351f",x"54361f",x"4e301c",x"4f331e",x"4e301b",x"51331d",x"4f311b",x"50321b",x"55341c",x"52331c",x"4e301a",x"50311c",x"50311b",x"51311b",x"512f18",x"52321c",x"56341c",x"5a371f",x"59361d",x"56341d",x"4f301a",x"6a4c33",x"6a4c33",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3f332a",x"3f332a",x"391f0e",x"3e2310",x"361e0d",x"3d2310",x"3c230f",x"3d220f",x"150e07",x"331d0d",x"3a220f",x"482914",x"241509",x"221309",x"221309",x"323232",x"333333",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"313131",x"333333",x"323232",x"313131",x"323232",x"202020",x"313131",x"3a3a3a",x"4a4a4a",x"454545",x"424242",x"424242",x"333333",x"3a3a3a",x"444444",x"414141",x"494949",x"404040",x"454545",x"4a4a4a",x"4b4b4b",x"444444",x"343434",x"313131",x"303030",x"5a5959",x"4a4846",x"393531",x"31302f",x"2f2f2f",x"393939",x"444240",x"3c3c3c",x"313131",x"333333",x"2d2e2e",x"303030",x"303030",x"2d2d2d",x"2f2f2f",x"2f2f2f",x"2c2c2c",x"323232",x"2e2e2e",x"333333",x"323232",x"323232",x"343434",x"333333",x"333333",x"4c2b13",x"1f1208",x"2d190b",x"2d190b",x"2d180a",x"1f1208",x"3d2310",x"3d2210",x"150e07",x"2f1a0b",x"3b2210",x"3e210f",x"442611",x"391f0e",x"3c2310",x"1b1008",x"3b2210",x"150e07",x"311b0b",x"28170b",x"39200f",x"432712",x"150e07",x"555555",x"555555",x"484848",x"202020",x"323232",x"333333",x"313131",x"333333",x"313131",x"333333",x"313131",x"313131",x"313131",x"2e2e2e",x"323232",x"313131",x"323232",x"313131",x"333333",x"323232",x"333333",x"323232",x"323232",x"343434",x"343434",x"313131",x"313131",x"303030",x"323232",x"333333",x"323232",x"313131",x"303030",x"323232",x"333333",x"313131",x"313131",x"303030",x"2c2c2c",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f3026",x"3f3026",x"311c0c",x"412511",x"321d0d",x"150e07",x"311c0c",x"2b180b",x"1f1208",x"150e07",x"38200e",x"150e07",x"150e07",x"000000",x"000000",x"24170d",x"24170d",x"2b1a0f",x"2a190c",x"2b190c",x"2b1a0d",x"28180c",x"2a190d",x"160e07",x"3d2310",x"503f33",x"462916",x"432917",x"372012",x"392211",x"371f10",x"27170b",x"855f42",x"986d4e",x"946949",x"885e42",x"946849",x"7e573c",x"9f7252",x"9b6f50",x"916648",x"926849",x"9b6f4d",x"986c4c",x"896044",x"896143",x"926b4c",x"8b6446",x"906547",x"8a6043",x"996d4c",x"916646",x"926748",x"936748",x"906546",x"745036",x"8f6547",x"966b4c",x"8c6142",x"986d4d",x"9e7353",x"95694a",x"976c4b",x"966b4b",x"875d3e",x"81583c",x"8b6244",x"976d4d",x"926849",x"956c4c",x"8c6244",x"855d43",x"805b40",x"5d412d",x"4d3625",x"4d3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412611",x"412611",x"150e07",x"150e07",x"150e07",x"4e453b",x"4e453b",x"46392e",x"4e2f1b",x"4e2f1b",x"2b190b",x"150e07",x"150e07",x"150e07",x"3d220f",x"3b210f",x"432712",x"402612",x"3f2410",x"3d220f",x"402511",x"412511",x"3c220f",x"3b200d",x"432712",x"1e1208",x"8e6748",x"8e6547",x"986c4c",x"9a6e4c",x"976b4b",x"7f583d",x"855d3f",x"653d1b",x"8c6143",x"885f42",x"8c6144",x"956a4b",x"906546",x"986b4a",x"8a6043",x"8c6244",x"916649",x"906649",x"916547",x"8c6244",x"8a6041",x"926949",x"966c4d",x"8d6242",x"986f50",x"8a6143",x"92694b",x"845d3f",x"8d6547",x"8f6647",x"8b6243",x"8a6042",x"906849",x"8a6244",x"8c6446",x"79553a",x"6e4d35",x"473120",x"45301f",x"45301f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3728",x"4e3728",x"472913",x"402410",x"371e0d",x"30190a",x"301b0c",x"3c220f",x"361e0d",x"3d220f",x"331e0e",x"3d2310",x"462812",x"2d1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"3b2210",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"391e0d",x"391e0d",x"50321f",x"2b1d12",x"433b33",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"150e07",x"1c1108",x"2c190b",x"2e1e12",x"42372e",x"42372e",x"000000",x"5b4b3f",x"5b4b3f",x"462a15",x"3f2613",x"3a2311",x"3d2411",x"402612",x"301c0d",x"301c0d",x"351f0e",x"2f1b0c",x"2b190b",x"331d0d",x"351f0f",x"2e1b0d",x"311c0d",x"2e1a0c",x"2d1a0b",x"2d1a0b",x"2f1b0c",x"361f0f",x"37200f",x"29180b",x"2f1b0c",x"2b190b",x"2a180b",x"2f1b0c",x"29180b",x"2a170a",x"2b180b",x"2b170a",x"2c180b",x"2c190b",x"28170a",x"2d190b",x"231409",x"2b180a",x"271609",x"271509",x"281609",x"211308",x"271509",x"241409",x"271509",x"28160a",x"29170a",x"221409",x"2d190b",x"29170a",x"2a170a",x"2c180b",x"251509",x"2f1a0c",x"2c190b",x"2e1a0b",x"2f1a0b",x"2a180b",x"402511",x"150e07",x"896546",x"876343",x"916c4c",x"876546",x"8b6646",x"866243",x"876243",x"876141",x"7e5c3d",x"755336",x"755236",x"835f40",x"846040",x"715136",x"7d5c40",x"816043",x"805e41",x"876445",x"876445",x"896445",x"8b6748",x"856142",x"8e6949",x"8c6849",x"8e694a",x"886546",x"8b6648",x"8b6646",x"916c4b",x"906d4c",x"8c6848",x"8c6748",x"896445",x"8b6646",x"8f6a4b",x"8b6748",x"8b6646",x"8a6646",x"8c6747",x"896342",x"815e3e",x"7e5a3b",x"795538",x"896343",x"8c6544",x"7a583a",x"8a6748",x"906b4b",x"8c6748",x"906a4b",x"8c6848",x"8d6747",x"926d4c",x"8c6646",x"956e4d",x"5c4d42",x"5c4d42",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"493b31",x"493b31",x"3d220f",x"412612",x"361e0d",x"2f1c0c",x"361e0d",x"3b200e",x"191008",x"321c0c",x"3a210f",x"4a2a14",x"26160a",x"231409",x"231409",x"333333",x"2d2520",x"313131",x"343434",x"333333",x"353535",x"313131",x"313131",x"343434",x"333333",x"323232",x"323232",x"313131",x"333333",x"2d2d2d",x"2c2c2c",x"2a2a2a",x"2e2e2e",x"303030",x"303030",x"313131",x"2d2d2d",x"313131",x"2f2f2f",x"4f4f4f",x"2e2e2e",x"313131",x"323232",x"323232",x"313131",x"313131",x"303030",x"323232",x"333333",x"323232",x"5e5e5d",x"504e4b",x"494541",x"302f2e",x"323232",x"343434",x"343434",x"323232",x"323232",x"323232",x"323232",x"353434",x"3d3935",x"4f4841",x"5e564e",x"5a5149",x"5a524a",x"4c463f",x"3b3938",x"343333",x"595959",x"343434",x"313131",x"323232",x"303030",x"492811",x"221308",x"2a180a",x"3a200e",x"331b0b",x"361f0e",x"3d220f",x"3d220f",x"150e07",x"351e0d",x"3b210f",x"3c220f",x"4e2b14",x"38200e",x"3e2310",x"150e07",x"3e2411",x"150e07",x"321c0b",x"150e07",x"39200e",x"432611",x"150e07",x"494949",x"494949",x"292929",x"323232",x"323232",x"313131",x"303030",x"303030",x"323232",x"313131",x"343434",x"333333",x"323232",x"333333",x"323232",x"343434",x"323232",x"323232",x"323232",x"333333",x"333333",x"313131",x"323232",x"323232",x"333333",x"343434",x"333333",x"323232",x"323232",x"313131",x"323232",x"333333",x"333333",x"313131",x"313131",x"313131",x"323232",x"2f2f2f",x"333333",x"343434",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2e25",x"3d2e25",x"2d1a0c",x"412612",x"412611",x"39200e",x"331c0d",x"301b0c",x"311c0c",x"341c0c",x"37200f",x"150e07",x"150e07",x"000000",x"000000",x"27180e",x"27180e",x"2e1c0f",x"2f1c0f",x"2c1b0d",x"2a190c",x"28180c",x"2f1c0d",x"160e07",x"341d0d",x"523d2f",x"452915",x"442916",x"362012",x"372011",x"382010",x"2e1b0d",x"8b6347",x"906748",x"7e573c",x"96694a",x"936847",x"8a6041",x"956b4c",x"9d7150",x"906547",x"865d40",x"7a5439",x"926648",x"976b4c",x"996f4f",x"956e4f",x"8b6245",x"8e6548",x"966a4a",x"986e4e",x"885e41",x"966d4d",x"976b4b",x"8e6445",x"896044",x"95694a",x"8e6346",x"885f41",x"916748",x"9c704f",x"9e7150",x"986b4b",x"9a6e4c",x"8e6444",x"8a6043",x"8a5f42",x"936a4a",x"8d6446",x"91684a",x"885f43",x"644430",x"835c41",x"5e422d",x"4e3625",x"4e3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2411",x"3f2411",x"150e07",x"150e07",x"150e07",x"50473e",x"50473e",x"40342b",x"4d2d15",x"4d2d15",x"28170a",x"150e07",x"150e07",x"150e07",x"3d2210",x"3a200e",x"412612",x"452913",x"3e2310",x"3e230f",x"3a200e",x"432611",x"3e230f",x"3a200e",x"402410",x"1c1108",x"8e6749",x"946a4a",x"8f6647",x"926849",x"926546",x"926647",x"8c6143",x"6f462f",x"855c3e",x"9e7151",x"936849",x"976b4b",x"916647",x"916646",x"875c40",x"865c40",x"936747",x"8c6346",x"876043",x"8d6345",x"855d42",x"8b6144",x"9c6f4f",x"8d6345",x"91684a",x"8a6143",x"815a3f",x"8e6445",x"8e6647",x"966b4a",x"92694a",x"8a6143",x"835c40",x"8b6345",x"8f6547",x"805a3f",x"714f37",x"422d1e",x"463020",x"463020",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3525",x"4e3525",x"482914",x"412511",x"311b0c",x"291509",x"311a0b",x"3d220f",x"3b200e",x"3c210f",x"452712",x"452812",x"482812",x"2a170a",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"150e07",x"150e07",x"150e07",x"170f07",x"29180b",x"29180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b200e",x"3b200e",x"553a28",x"2d1d11",x"463e35",x"150e07",x"150e07",x"150e07",x"150e07",x"26160a",x"150e07",x"150e07",x"150e07",x"1a1008",x"321c0c",x"2d1d13",x"3f352d",x"3f352d",x"000000",x"5b4a3e",x"5b4a3e",x"3c2311",x"2d1b0d",x"311d0e",x"2f1b0c",x"2e1a0c",x"2e1b0c",x"2f1b0d",x"2d1b0d",x"26170b",x"2f1b0c",x"2b190b",x"27170a",x"2c1a0c",x"1e1309",x"22150a",x"2a190c",x"1c1108",x"26160a",x"23150a",x"29190c",x"211409",x"27170b",x"191008",x"24150a",x"28180b",x"26160b",x"29180b",x"26160a",x"2d1b0d",x"2a190c",x"2b190b",x"2b190b",x"29180a",x"25150a",x"221409",x"251509",x"2a180b",x"1c1108",x"1d1108",x"241509",x"221409",x"241509",x"211409",x"29180b",x"24150a",x"28170b",x"25160a",x"26160a",x"2c190b",x"28170a",x"241509",x"1f1309",x"28170a",x"2a190b",x"221409",x"3b220f",x"150e07",x"815d3f",x"7e5c3f",x"805e40",x"805d3e",x"825f41",x"846041",x"7f5b3d",x"7b583a",x"815d3e",x"815e3e",x"755338",x"836141",x"846141",x"886445",x"866445",x"7b593d",x"78583b",x"79593c",x"846142",x"825f41",x"846244",x"856444",x"8d6a4a",x"876344",x"805d41",x"8b6748",x"846142",x"805c3e",x"7f5d3d",x"876243",x"8d6746",x"866244",x"805d3f",x"876344",x"856143",x"825f40",x"825f41",x"825f41",x"7e5a3d",x"815d3e",x"866141",x"886342",x"805c3e",x"8b6745",x"896444",x"8f6949",x"886446",x"825f41",x"886444",x"8a6545",x"8a6544",x"8a6646",x"936e4d",x"936e4c",x"946f4d",x"605145",x"605145",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"473a2f",x"473a2f",x"3d220f",x"3d220f",x"371e0d",x"361d0c",x"3a200e",x"361e0d",x"311c0c",x"39200e",x"371f0e",x"472912",x"2d190b",x"251509",x"251509",x"323232",x"333333",x"323232",x"333333",x"333333",x"313131",x"323232",x"323232",x"323232",x"303030",x"333333",x"323232",x"323232",x"343434",x"313131",x"2f2f2f",x"2e2e2e",x"2e2e2e",x"2b2b2b",x"313131",x"2d2d2d",x"303030",x"333333",x"2e2e2e",x"323232",x"313131",x"323231",x"333333",x"323232",x"313131",x"2f2f2f",x"333333",x"323232",x"333333",x"2e2e2e",x"3a3835",x"44413d",x"413d3a",x"333332",x"323232",x"333333",x"323232",x"313131",x"313131",x"303030",x"323232",x"3d3c3b",x"4e4a46",x"5d5751",x"605851",x"615a52",x"5a544d",x"534f4b",x"3b3938",x"333232",x"424242",x"343434",x"323232",x"343434",x"333333",x"442510",x"1d1108",x"2a180a",x"341c0c",x"321b0b",x"3c2310",x"3c210f",x"3a200e",x"2f1c0d",x"371e0d",x"3b210f",x"351e0d",x"4e2b14",x"331c0c",x"351d0d",x"2e190b",x"432712",x"39200e",x"311a0b",x"150e07",x"371f0e",x"452712",x"150e07",x"3c3c3c",x"3c3c3c",x"1d1d1d",x"282828",x"313131",x"2f2f2f",x"333333",x"323232",x"323232",x"323232",x"323232",x"2d2d2d",x"2d2e2e",x"323232",x"313131",x"303030",x"323232",x"333333",x"323232",x"313131",x"2f2f2f",x"343434",x"323232",x"333333",x"313131",x"313131",x"333333",x"323232",x"333333",x"313131",x"323232",x"323232",x"312a25",x"313131",x"323232",x"323232",x"333333",x"323232",x"303030",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"41332a",x"41332a",x"2c190c",x"402411",x"3f2410",x"391f0e",x"39200e",x"351e0d",x"3e2310",x"381f0e",x"3a210f",x"150e07",x"150e07",x"000000",x"000000",x"29190e",x"29190e",x"311e10",x"331f11",x"301d0f",x"2b1a0e",x"28180c",x"27180b",x"18110a",x"311b0c",x"584335",x"452815",x"412816",x"3d2413",x"321e10",x"331d0f",x"25150a",x"91674a",x"835d41",x"916547",x"986b4b",x"956747",x"8a6042",x"7a553c",x"986c4d",x"906546",x"825c40",x"885e41",x"996c4c",x"9b704f",x"9a6f4f",x"966d4d",x"8e6446",x"986e4f",x"976d4e",x"9e7251",x"8a6041",x"936849",x"956a4a",x"976b4b",x"94694a",x"9a6f4f",x"8e6547",x"7d5238",x"95694a",x"966c4c",x"906646",x"865c40",x"916647",x"80593c",x"906647",x"926849",x"906648",x"8a6144",x"956b4c",x"8e6445",x"8b6446",x"7f5a3f",x"5f422c",x"4d3726",x"4d3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2511",x"3f2511",x"150e07",x"150e07",x"150e07",x"4d433a",x"4d433a",x"40342a",x"55331c",x"55331c",x"321c0d",x"150e07",x"150e07",x"150e07",x"472814",x"3f230f",x"412511",x"472a14",x"3c210f",x"391f0e",x"3e2310",x"3f2310",x"3f2310",x"3f2410",x"381e0d",x"1e1208",x"8e6649",x"8e6647",x"936949",x"976a4a",x"8b6043",x"986b4a",x"966948",x"8f6545",x"8b6143",x"9b6f4d",x"9a6f4e",x"986d4e",x"8b6041",x"96694a",x"885e3f",x"8e6446",x"8e6344",x"946849",x"81593e",x"8d6245",x"876143",x"8e6344",x"7d583d",x"93694a",x"a17452",x"855c40",x"8b6143",x"996f4f",x"976d4d",x"966b4c",x"906647",x"8b6243",x"926748",x"8a6143",x"8d6446",x"805a3e",x"6a4931",x"432e1e",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533929",x"533929",x"472813",x"3a210f",x"361d0d",x"361d0c",x"3b200e",x"3b210f",x"3c220f",x"3c210e",x"3d2310",x"422611",x"482912",x"331c0c",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"170f07",x"160f07",x"180f07",x"181007",x"2b180b",x"2b180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412411",x"412411",x"5f493a",x"2a1b11",x"4c4238",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"1a1008",x"321d0e",x"312116",x"40372e",x"40372e",x"000000",x"574638",x"574638",x"37200f",x"28180b",x"2d1b0c",x"2b190c",x"301c0d",x"2f1b0c",x"2e1b0c",x"2c1a0c",x"29180b",x"2a180b",x"25160a",x"27170a",x"2a190b",x"26160a",x"211409",x"211409",x"1f1309",x"24150a",x"2a180b",x"29180b",x"2a180b",x"28170b",x"27170b",x"1c1208",x"1f1309",x"27170b",x"2d1a0c",x"211409",x"2a180b",x"27160a",x"2a190b",x"2c1a0b",x"26170a",x"2c1a0c",x"29180b",x"26160a",x"26160a",x"241509",x"26160a",x"26160a",x"24150a",x"27170a",x"221409",x"27170a",x"24150a",x"25160a",x"27170a",x"2a180b",x"24150a",x"24150a",x"211409",x"221409",x"29170b",x"26160a",x"241509",x"341d0d",x"150e07",x"825d40",x"815d3f",x"805e40",x"7f5b3c",x"7b593a",x"805c3e",x"7c5a3c",x"7d5b3d",x"7c593c",x"7a593b",x"765438",x"7a593c",x"846141",x"7e5b3e",x"886545",x"7e5c3f",x"7a593c",x"846243",x"866345",x"876345",x"815e3f",x"815d3f",x"7f5d3f",x"866343",x"886546",x"886445",x"815f41",x"815e41",x"7d5b3d",x"735336",x"805b3e",x"7f5c3d",x"805c3f",x"78573a",x"846042",x"7e5b3c",x"7a583a",x"7d5a3d",x"7b593b",x"845f40",x"846041",x"815d3e",x"835f41",x"8c6746",x"866242",x"876242",x"8d6848",x"896444",x"876343",x"8d6847",x"926c4c",x"8e6949",x"8a6444",x"886443",x"8c6746",x"6a5444",x"6a5444",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d3c2f",x"4d3c2f",x"3f2310",x"442813",x"341d0c",x"39200e",x"341c0c",x"311c0c",x"3c2310",x"3e2310",x"361e0d",x"41230f",x"2e1a0c",x"27160a",x"27160a",x"333130",x"393939",x"303030",x"323232",x"323232",x"303030",x"303030",x"323232",x"2e2e2e",x"323232",x"323232",x"2d2d2d",x"30302f",x"313131",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"303030",x"313131",x"333333",x"32312f",x"515151",x"313131",x"323232",x"313131",x"323232",x"323232",x"323232",x"2f2f2f",x"303030",x"313131",x"3f3f3f",x"525252",x"484747",x"4b4b4b",x"404040",x"323232",x"323232",x"323232",x"333333",x"313131",x"3a3a3a",x"565656",x"5c5c5c",x"505050",x"505050",x"545454",x"555351",x"4f4f4f",x"505050",x"525252",x"545454",x"636363",x"393939",x"2f2f2f",x"323232",x"333333",x"482811",x"251509",x"28170a",x"361d0c",x"361d0c",x"3c210f",x"371f0d",x"311c0c",x"3a210f",x"3b220f",x"3f2411",x"3e220f",x"512e15",x"331c0c",x"3a200e",x"150e07",x"3a210f",x"2d190b",x"2f190b",x"150e07",x"2e1a0c",x"422511",x"150e07",x"494949",x"484848",x"313131",x"323232",x"2f2f2f",x"313131",x"333333",x"333333",x"363535",x"43403d",x"353434",x"313131",x"262626",x"323232",x"333333",x"323232",x"343434",x"2d2d2d",x"303030",x"303030",x"323232",x"343434",x"323232",x"333333",x"323232",x"323232",x"323232",x"303030",x"323232",x"333333",x"303030",x"353535",x"313131",x"313232",x"333333",x"313131",x"323232",x"363636",x"323232",x"323232",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e3027",x"3e3027",x"2e1a0c",x"452914",x"402411",x"150e07",x"361e0d",x"371f0e",x"311c0c",x"38200e",x"361e0d",x"150e07",x"150e07",x"000000",x"000000",x"2a190e",x"2a190e",x"331f11",x"341f10",x"2f1c0f",x"301d0f",x"2a1a0e",x"21150b",x"181009",x"3b210f",x"5c4333",x"432716",x"3b2314",x"3a2312",x"372012",x"2e1a0e",x"2d190c",x"8e6649",x"986c4d",x"8f6445",x"976948",x"936747",x"8d6143",x"976c4b",x"976b4c",x"906547",x"8c6245",x"92694b",x"936746",x"976b4c",x"906647",x"8e6548",x"8b6144",x"956c4e",x"a07452",x"9a6d4b",x"8d6243",x"976c4c",x"8c6244",x"926748",x"94694a",x"9d7150",x"906648",x"8c6142",x"996e4d",x"976b4b",x"976c4b",x"946a4a",x"875f43",x"8f6547",x"8d6445",x"8d6346",x"926849",x"805a3f",x"9b7151",x"8f6546",x"875f43",x"7e5a3f",x"5d402c",x"4f3625",x"4f3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"382110",x"382110",x"150e07",x"150e07",x"150e07",x"4c4339",x"4c4339",x"3e3127",x"52331e",x"52331e",x"341d0d",x"150e07",x"150e07",x"150e07",x"472913",x"3c210f",x"442813",x"442813",x"391f0e",x"3d2310",x"422511",x"402410",x"412511",x"412410",x"391f0d",x"1a1008",x"966d4f",x"906547",x"936849",x"986d4c",x"906647",x"9a6e4e",x"926645",x"956949",x"845c40",x"9b6f4e",x"a37756",x"9b7151",x"8a5f42",x"936746",x"865a3e",x"8a5f41",x"8e6445",x"946849",x"906547",x"976c4c",x"9d7351",x"885f41",x"976b4c",x"916646",x"976e4d",x"8c6345",x"875e42",x"946a4c",x"936749",x"926849",x"94684a",x"96694b",x"916748",x"906648",x"8e6647",x"7e593e",x"704e36",x"402c1d",x"442f1e",x"442f1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533827",x"533827",x"4a2b14",x"3c220f",x"381e0d",x"381f0d",x"391f0e",x"3c210f",x"3f2410",x"39200e",x"452812",x"472913",x"472812",x"301b0b",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"201308",x"201309",x"150e07",x"150e07",x"1a1008",x"281609",x"000000",x"201208",x"150e07",x"150e07",x"150e07",x"150e07",x"402411",x"402411",x"5e4332",x"2a1d14",x"51473d",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"150e07",x"150e07",x"150e07",x"150e07",x"311d0e",x"322218",x"42382e",x"42382e",x"000000",x"544134",x"544134",x"321d0d",x"24150a",x"301c0d",x"2b190c",x"2f1b0c",x"2c190b",x"2b190b",x"1f1309",x"2e1a0c",x"241509",x"28170a",x"231409",x"1b0f07",x"180f07",x"201208",x"201309",x"211309",x"221409",x"211309",x"251509",x"25150a",x"221409",x"28170b",x"1d1108",x"1f1309",x"241509",x"211409",x"1a1008",x"251509",x"29170a",x"27170a",x"29170a",x"251509",x"251509",x"211308",x"211309",x"231509",x"29170a",x"28170a",x"27170b",x"201309",x"25160a",x"27170a",x"26160a",x"241509",x"27160a",x"25160a",x"24150a",x"1d1208",x"27170b",x"28180b",x"24150a",x"25160a",x"201409",x"221509",x"412611",x"150e07",x"876241",x"836141",x"876343",x"835f40",x"856141",x"866242",x"886442",x"805d40",x"886443",x"835e3d",x"725235",x"765536",x"815d3d",x"846042",x"846244",x"76563a",x"77573b",x"7e5c3e",x"8b6749",x"8b6748",x"896647",x"886546",x"7e5a3d",x"7d5a3d",x"805c3e",x"845f42",x"7f5c3e",x"886446",x"866243",x"8a6647",x"8b6748",x"856242",x"7e5c3d",x"856242",x"856141",x"805d3e",x"825f3f",x"846041",x"866341",x"886445",x"8d6746",x"846040",x"7a5837",x"86613f",x"8a6441",x"876345",x"946f4d",x"846142",x"856143",x"916a48",x"95704e",x"926d4c",x"926c4c",x"916c4c",x"896343",x"644f41",x"644f41",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a3b2f",x"4a3b2f",x"40230f",x"452813",x"381e0d",x"3f230f",x"3e230f",x"3b210f",x"3f2411",x"3e2410",x"3c220f",x"3e210e",x"2b180b",x"241409",x"241409",x"323232",x"323232",x"333333",x"3e3f3f",x"323232",x"343434",x"313131",x"323232",x"323232",x"393736",x"544e47",x"423f3b",x"3f3c39",x"3e3b38",x"323232",x"323232",x"2f2f2f",x"292929",x"323232",x"2e2e2d",x"2f2f2e",x"353231",x"5a524a",x"5d554e",x"57514a",x"544d46",x"544d47",x"5e564e",x"5d554d",x"5d564e",x"5d554d",x"5d564e",x"5b534b",x"5f574f",x"5e564e",x"595148",x"5b534b",x"605951",x"514b44",x"333333",x"302e2c",x"312721",x"313131",x"313131",x"323232",x"5e5e5e",x"5c5c5a",x"504d4a",x"5c5651",x"544b42",x"585047",x"625c55",x"58534e",x"565454",x"504f4e",x"605f5f",x"323232",x"323232",x"323232",x"333333",x"40230f",x"221409",x"2d190b",x"2f180a",x"371e0c",x"402410",x"371f0e",x"391f0e",x"39210f",x"3c220f",x"412511",x"402310",x"4f2d15",x"331c0c",x"341c0c",x"27170b",x"3d2310",x"150e07",x"291609",x"1f1208",x"341d0d",x"3b210f",x"150e07",x"4c4c4c",x"484848",x"343434",x"323232",x"333333",x"333333",x"323232",x"343434",x"393838",x"54514e",x"444343",x"333333",x"2d2d2d",x"333333",x"323232",x"323232",x"333333",x"333333",x"323232",x"323232",x"313131",x"333333",x"333333",x"323232",x"3c3c3c",x"333333",x"343434",x"323232",x"323232",x"333333",x"303030",x"353535",x"313131",x"313232",x"333333",x"313131",x"323232",x"363636",x"323232",x"323232",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e3127",x"3e3127",x"301c0d",x"472a14",x"331e0e",x"180f07",x"321c0d",x"3a200e",x"201309",x"150e07",x"3a200e",x"191008",x"191008",x"000000",x"000000",x"2d1c10",x"2d1c10",x"372314",x"351f10",x"2e1a0e",x"2f1c0f",x"2a1a0e",x"29190e",x"181009",x"341d0d",x"5a4334",x"432715",x"3d2414",x"3a2313",x"382212",x"311b0e",x"28170b",x"865e42",x"966b4d",x"8a6143",x"9d714e",x"906445",x"865d3f",x"9a6f4e",x"9d7152",x"8e6346",x"8e6346",x"9e7250",x"885e40",x"94694a",x"91684a",x"986f4f",x"9b6f4e",x"986e4f",x"9a6f4f",x"916646",x"8d6345",x"986d4b",x"8e6345",x"916646",x"926849",x"966c4d",x"916748",x"926748",x"9a6f4d",x"936849",x"956949",x"926647",x"8d6345",x"966a4a",x"926849",x"966a4b",x"986d4c",x"936748",x"9a7051",x"8b6144",x"8a6244",x"805b40",x"5a3e29",x"4e3726",x"4e3726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200f",x"38200f",x"150e07",x"150e07",x"150e07",x"4e453c",x"4e453c",x"41352b",x"4f2f19",x"4f2f19",x"271609",x"150e07",x"150e07",x"150e07",x"442612",x"3d220f",x"482a14",x"422612",x"3e2310",x"402410",x"422611",x"442712",x"442711",x"3e220f",x"3c200e",x"211309",x"956c4d",x"8f6447",x"926748",x"996d4c",x"8d6243",x"986d4e",x"926646",x"8a6044",x"8f6447",x"906647",x"9d7150",x"9c704e",x"8d6343",x"805a3e",x"8d6342",x"875b3f",x"8e6444",x"8b6447",x"845d41",x"996c4c",x"9b7150",x"835b3d",x"956a4b",x"93694a",x"9c7251",x"936849",x"8b6245",x"916747",x"8f6546",x"8d6346",x"9a6f4e",x"946949",x"946a4c",x"906749",x"8b6447",x"835e42",x"6f4e36",x"483221",x"483221",x"483221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583b29",x"583b29",x"4c2d15",x"3b200e",x"3e220f",x"3a200e",x"351d0d",x"39200e",x"3a210f",x"3c210e",x"412511",x"432711",x"40220e",x"301c0d",x"25150a",x"150e07",x"150e07",x"150e07",x"000000",x"29160a",x"29160a",x"150e07",x"160f07",x"281609",x"281609",x"201208",x"201208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"412410",x"593922",x"35251b",x"50453a",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"191008",x"2a190c",x"34251b",x"443a30",x"443a30",x"000000",x"503b2e",x"503b2e",x"311c0c",x"241509",x"231409",x"251509",x"28160a",x"231409",x"251509",x"211309",x"241509",x"2c190b",x"2c190b",x"2b190b",x"2a180b",x"2a180b",x"27160a",x"28170a",x"25160a",x"221409",x"231409",x"231509",x"231509",x"241509",x"1d1208",x"231509",x"25160a",x"211409",x"25150a",x"231409",x"2d1a0b",x"27170a",x"2c1a0b",x"28170a",x"1e1208",x"28170a",x"201208",x"241509",x"27170a",x"25160a",x"241509",x"27170a",x"251509",x"26160a",x"221409",x"241509",x"231509",x"211409",x"1d1108",x"211409",x"25160a",x"27170a",x"1b1108",x"27170a",x"27170a",x"201309",x"180f07",x"3c200e",x"150e07",x"7e5b3d",x"815d3f",x"825d3f",x"805c3e",x"856143",x"805c3f",x"805d3f",x"815d3f",x"805d3f",x"825c3d",x"785838",x"765436",x"735335",x"79583c",x"735336",x"775639",x"765438",x"77573b",x"7c593c",x"846243",x"805d3f",x"825f41",x"805d3e",x"805c3e",x"7d5a3d",x"775539",x"775639",x"7c5a3d",x"7f5c3e",x"7e5b3d",x"7a583a",x"7f5b3e",x"79583a",x"815d3f",x"805d3e",x"815d3f",x"876243",x"7e5c3d",x"825f40",x"805c3e",x"836040",x"825d3c",x"7c5a39",x"815e3c",x"835e3d",x"825f40",x"825e3f",x"805d3d",x"7b573a",x"846042",x"8a6444",x"886545",x"815d3f",x"876343",x"876241",x"5b4b3f",x"5b4b3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"493b2f",x"493b2f",x"3b200e",x"432612",x"381f0d",x"3d220f",x"3c210f",x"371e0d",x"3f2411",x"3c230f",x"402410",x"422410",x"2d190b",x"241509",x"241509",x"32302f",x"333333",x"313131",x"313131",x"323232",x"636363",x"5d5d5c",x"313131",x"5a5a5a",x"3f3933",x"66625e",x"595756",x"39332d",x"241d17",x"3d3c3a",x"4a4a4a",x"2f2f2f",x"303030",x"454545",x"585858",x"535252",x"4c4c4b",x"564e45",x"52493f",x"4d443b",x"59514a",x"635c57",x"564d43",x"6c6660",x"6a635c",x"605750",x"665e56",x"6d6660",x"6d6660",x"6d6760",x"696159",x"675f57",x"676059",x"59524b",x"2f2d2c",x"313131",x"2f2f2f",x"313131",x"323232",x"323232",x"383838",x"4a4948",x"534f4c",x"605a55",x"645e58",x"645d57",x"5d5852",x"55514e",x"474645",x"3b3a3a",x"4e4e4e",x"2f2f2f",x"323232",x"333333",x"303030",x"492812",x"221409",x"251509",x"351c0b",x"341c0c",x"3b210f",x"371f0e",x"311b0c",x"371f0e",x"331c0d",x"3e2310",x"3e220f",x"4f2d15",x"361e0d",x"351d0d",x"311d0d",x"3b210f",x"150e07",x"2a160a",x"2b180b",x"331d0d",x"3d220f",x"150e07",x"150e07",x"565656",x"4e4e4e",x"313131",x"3e3e3e",x"323232",x"313131",x"333333",x"3a3837",x"595654",x"4c4c4c",x"373737",x"2f2f2f",x"333333",x"323232",x"333333",x"323232",x"333333",x"313131",x"333333",x"333333",x"313131",x"323232",x"3c3c3c",x"404040",x"343434",x"323232",x"333333",x"333333",x"5c544d",x"605851",x"615952",x"625b54",x"655e57",x"675f59",x"69625c",x"6a635c",x"645d56",x"615a52",x"5d554c",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"43362c",x"43362c",x"29180b",x"442813",x"3c2311",x"331e0e",x"3a210f",x"3b200f",x"2b190b",x"2f1b0c",x"381f0d",x"180f07",x"180f07",x"000000",x"000000",x"301d11",x"301d11",x"372213",x"321e10",x"362011",x"2d1b0e",x"2c1a0e",x"28190e",x"18110a",x"351d0d",x"594131",x"452a16",x"402716",x"3e2414",x"352012",x"321b0e",x"27170b",x"7b5438",x"886044",x"855c3f",x"9c6f4d",x"895e41",x"8b6141",x"9d7151",x"9e7251",x"8f6445",x"8d6143",x"9b714f",x"896042",x"8c6344",x"926849",x"986c4c",x"9a704f",x"916748",x"936848",x"916647",x"78533a",x"8d6345",x"855b3f",x"875d3f",x"8a6043",x"976b4b",x"976d4c",x"936747",x"946849",x"976b4b",x"8d6345",x"875d3f",x"906547",x"8e6445",x"8a6144",x"906648",x"906648",x"916748",x"986e4e",x"916647",x"79543b",x"6f4e34",x"61432e",x"503827",x"503827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2210",x"3d2210",x"150e07",x"150e07",x"150e07",x"4f453c",x"4f453c",x"382f26",x"533117",x"533117",x"28170a",x"150e07",x"150e07",x"150e07",x"482913",x"3f230f",x"472913",x"432712",x"422611",x"3e2310",x"402410",x"432611",x"432611",x"3c210e",x"3b200e",x"1d1108",x"986f50",x"8e6446",x"8c6242",x"946847",x"976c4c",x"9b704f",x"9b7050",x"8e6443",x"926745",x"976a47",x"956947",x"986b4b",x"8e6445",x"896043",x"8b6142",x"83593d",x"906748",x"896345",x"84593e",x"8c6243",x"986e4d",x"885f40",x"966a4b",x"986d4e",x"986d4c",x"996e4e",x"976d4c",x"996e4d",x"8d6345",x"8c6244",x"8f6546",x"936849",x"8f6647",x"906647",x"896143",x"835d40",x"714f37",x"432d1d",x"432d1d",x"432d1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e3423",x"4e3423",x"462813",x"361e0d",x"3c220f",x"39200e",x"381f0e",x"402511",x"39200e",x"341c0c",x"422611",x"422611",x"43240f",x"2b180b",x"1d1108",x"150e07",x"181009",x"181009",x"000000",x"1f1208",x"2c1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"351f0e",x"351f0e",x"24150a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"52321d",x"32261d",x"574d43",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0c",x"150e07",x"150e07",x"150e07",x"1a1008",x"28170b",x"35261c",x"453c33",x"453c33",x"000000",x"5a3f2d",x"5a3f2d",x"331e0e",x"2a180b",x"24150a",x"27170a",x"24150a",x"321e0e",x"2d1c0d",x"27170a",x"1d1208",x"27170a",x"2a190b",x"231509",x"29180b",x"28170a",x"26170a",x"26160a",x"28170b",x"1b1108",x"24150a",x"29180b",x"23150a",x"211409",x"25160a",x"25160a",x"241509",x"211409",x"1e1208",x"211309",x"221409",x"201309",x"24150a",x"25150a",x"1f1309",x"27170a",x"211309",x"1e1208",x"25150a",x"29180b",x"1f1208",x"1e1208",x"231409",x"231409",x"1e1108",x"241509",x"201309",x"211309",x"1d1108",x"241509",x"211409",x"211409",x"231409",x"1a1008",x"1c1108",x"201309",x"201309",x"3d210f",x"150e07",x"815d3f",x"7b593c",x"745439",x"765439",x"7d5a3e",x"765439",x"66462d",x"7c5a3c",x"7b583b",x"785637",x"815d3c",x"805c3d",x"715236",x"79573a",x"7a593a",x"7f5b3d",x"846142",x"7d5b3d",x"815e41",x"7d5c3e",x"715136",x"77573a",x"735337",x"765539",x"78563a",x"755438",x"805d3e",x"805d3e",x"805c3e",x"815e3f",x"7b593c",x"7a583c",x"7b593c",x"7a583b",x"7a583b",x"765439",x"7d5b3e",x"765438",x"64442b",x"7d5a3d",x"735337",x"755335",x"86603e",x"8a6441",x"7d5b3d",x"805c3e",x"805d3c",x"866141",x"8e6947",x"896442",x"8e6948",x"836041",x"815d3f",x"856140",x"7f5b3d",x"604e41",x"604e41",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a3b2f",x"4a3b2f",x"422510",x"462812",x"3d220f",x"391f0d",x"39200e",x"391f0d",x"422511",x"3c230f",x"422611",x"412310",x"301b0c",x"25150a",x"25150a",x"333333",x"323232",x"333333",x"313131",x"323232",x"373636",x"323232",x"323232",x"474747",x"676562",x"6a6764",x"4a4846",x"4e4b48",x"5f5e5e",x"535353",x"323232",x"313131",x"303030",x"2f2f2f",x"3f3f3e",x"40403f",x"41403f",x"5e5751",x"5a544e",x"59524c",x"5d5852",x"655f59",x"6c6761",x"68625c",x"675f59",x"635b54",x"605951",x"655e56",x"5e564e",x"615a52",x"605850",x"5d554d",x"5e564e",x"514b45",x"2b2b2b",x"323232",x"313131",x"333333",x"323232",x"323232",x"434343",x"50504f",x"52504f",x"5b5752",x"645e57",x"68615a",x"645d57",x"5d5853",x"4a4947",x"434343",x"545454",x"313131",x"303030",x"313131",x"333333",x"492812",x"27160a",x"221309",x"321a0b",x"311b0b",x"2f1a0b",x"321c0d",x"2b180a",x"361e0d",x"3c220f",x"3f2411",x"3a1f0d",x"522f15",x"331b0b",x"3b210f",x"27170a",x"3a220f",x"150e07",x"281609",x"341d0d",x"3b2210",x"29170a",x"150e07",x"150e07",x"454545",x"5c5c5c",x"4e4e4e",x"323232",x"323232",x"333333",x"313131",x"3c3a37",x"3f3c3a",x"414140",x"323232",x"333333",x"303030",x"323232",x"323232",x"323232",x"313131",x"333333",x"333333",x"2e2e2e",x"323232",x"333333",x"343434",x"323232",x"333333",x"323232",x"323232",x"5d564e",x"5c544d",x"605851",x"615952",x"625b54",x"655e57",x"675f59",x"69625c",x"6a635c",x"645d56",x"615a52",x"5d554c",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"47382e",x"47382e",x"1f1209",x"3c2310",x"412612",x"331d0d",x"402511",x"3d220f",x"1d1208",x"2d190b",x"341c0c",x"190f07",x"190f07",x"000000",x"000000",x"301e11",x"301e11",x"352012",x"382313",x"362113",x"301d11",x"2b1a0d",x"27180d",x"181009",x"3b210f",x"503e31",x"4d2e18",x"3f2614",x"392212",x"392212",x"371f0f",x"301c0e",x"6c4931",x"8c6446",x"906446",x"9b6d4c",x"976a4b",x"81563b",x"9e7151",x"9d704f",x"865d40",x"855c40",x"956c4c",x"916646",x"996d4c",x"986d4d",x"976c4d",x"966c4d",x"966a4a",x"936849",x"916748",x"94694a",x"946748",x"8f6648",x"8a5f41",x"8f6647",x"956a4b",x"956a4b",x"986b4b",x"936847",x"956949",x"80583d",x"845a3d",x"7a553b",x"815c3f",x"976d4d",x"7c563b",x"8f6545",x"95694b",x"9c7252",x"896043",x"745139",x"7d593e",x"593d29",x"4f3826",x"4f3826",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2411",x"3f2411",x"150e07",x"150e07",x"150e07",x"4c4339",x"4c4339",x"3c3027",x"51301a",x"51301a",x"381f0e",x"150e07",x"150e07",x"150e07",x"512d15",x"3d220f",x"422511",x"472914",x"432612",x"3d220f",x"3d220f",x"40240f",x"432511",x"3f230e",x"3b200d",x"201309",x"936b4d",x"906547",x"956948",x"956b4a",x"966b4a",x"996d4d",x"9b6f4e",x"8d6341",x"8d6242",x"986b48",x"916644",x"a17554",x"895e41",x"906647",x"8a5f41",x"80563c",x"9b6f4e",x"9a7050",x"8d6345",x"8b6143",x"9c6f4f",x"885f41",x"95694b",x"845c40",x"9e7451",x"986d4d",x"865d40",x"8f6547",x"9e7150",x"956a4a",x"956c4c",x"8a5f42",x"835c3f",x"906647",x"845d41",x"876145",x"6b4a32",x"493221",x"473120",x"473120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583a28",x"583a28",x"452812",x"341c0c",x"412611",x"361e0d",x"3e2310",x"3b210f",x"3f2410",x"31190a",x"3b200e",x"39200e",x"3b210e",x"2c190b",x"1b1008",x"150e07",x"170f08",x"170f08",x"000000",x"27160a",x"25150a",x"150e07",x"150e07",x"1b1108",x"150e07",x"361e0d",x"361d0d",x"371e0d",x"150e07",x"150e07",x"1c1108",x"150e07",x"150e07",x"55351f",x"36291f",x"584d43",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"150e07",x"1c1108",x"2f1b0e",x"37291e",x"453c32",x"453c32",x"000000",x"624330",x"624330",x"331d0d",x"29180b",x"1e1209",x"2b1a0c",x"2d1b0c",x"321d0d",x"29180b",x"2a190c",x"27170a",x"2c1a0c",x"2a180b",x"28170b",x"1e1208",x"25160a",x"1d1108",x"2b190b",x"2d1a0c",x"191008",x"23150a",x"25160a",x"2e1b0d",x"24150a",x"201309",x"24150a",x"211409",x"27160a",x"221409",x"201309",x"1b1108",x"1b1008",x"2a180b",x"27160a",x"2d190b",x"27170a",x"231409",x"221409",x"221409",x"29180b",x"27170a",x"25160a",x"27160a",x"241509",x"251509",x"241509",x"26160a",x"25150a",x"221409",x"27160a",x"241509",x"28170a",x"241509",x"211309",x"241509",x"27160a",x"221309",x"452712",x"150e07",x"815d3f",x"7d5a3d",x"7b593c",x"856141",x"835f40",x"805d3f",x"7b583a",x"785438",x"765336",x"8a6445",x"886544",x"866243",x"815f3f",x"825f41",x"866243",x"856344",x"856344",x"826041",x"7f5c3d",x"7a583b",x"7a583b",x"805d3e",x"7f5b3e",x"7f5b3d",x"7b593c",x"815d3f",x"815d3f",x"845f40",x"79583a",x"7d5b3d",x"805c3f",x"7d5b3d",x"7c5a3c",x"7a583b",x"805b3e",x"78573a",x"805d3f",x"815e3f",x"7a583a",x"755236",x"775436",x"886444",x"8b6748",x"8c6746",x"8c6645",x"8e6847",x"8f6a47",x"936d4c",x"886547",x"8f6948",x"896342",x"866142",x"876142",x"856040",x"886343",x"5f4e41",x"5f4e41",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d3e32",x"4d3e32",x"432611",x"412410",x"3c210f",x"381f0d",x"391f0e",x"2f1a0b",x"3f2310",x"3e2310",x"3f2410",x"462711",x"2e1a0c",x"241409",x"241409",x"313131",x"34302d",x"313131",x"333333",x"2b2b2b",x"5b5b5b",x"525252",x"333333",x"585858",x"505050",x"565656",x"5e5e5e",x"5c5c5c",x"606060",x"5c5c5c",x"414141",x"313131",x"4f4f4f",x"545454",x"5a5a5a",x"5a5a5a",x"535353",x"5c5b5b",x"5e5d5c",x"5f5f5f",x"616161",x"5e5d5c",x"626161",x"606060",x"666564",x"666464",x"636363",x"5e5e5e",x"5a5a5a",x"5c5c5c",x"5b5a59",x"5d5c5a",x"5a5a59",x"454545",x"333333",x"333333",x"313131",x"313131",x"313131",x"323232",x"323232",x"3a3938",x"4b4845",x"57514c",x"5d554e",x"645d55",x"615a54",x"595551",x"3b3938",x"333232",x"4b4b4b",x"313131",x"2f2f2f",x"323232",x"343434",x"492912",x"27160a",x"241308",x"321a0b",x"311b0b",x"361e0d",x"39200e",x"361d0d",x"3c210f",x"412612",x"3a210f",x"361c0c",x"4a2912",x"331c0c",x"2c190b",x"3f2411",x"3f2410",x"351d0c",x"150e07",x"27160a",x"321c0d",x"29170a",x"150e07",x"150e07",x"383838",x"484848",x"3b3b3b",x"333333",x"323232",x"323232",x"343434",x"323232",x"323232",x"313131",x"5d554d",x"4c4843",x"3e3b38",x"504a43",x"323232",x"333333",x"323232",x"313131",x"323232",x"313131",x"343333",x"333333",x"5d564e",x"5c554d",x"564f47",x"565049",x"565049",x"5d554e",x"645e56",x"625b53",x"5c544c",x"665f58",x"645d56",x"686159",x"676059",x"6a645e",x"645d56",x"615951",x"5c554c",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3e33",x"4d3e33",x"26160a",x"412511",x"39210f",x"3f2411",x"412511",x"361e0d",x"150e07",x"190f07",x"341c0c",x"150e07",x"150e07",x"000000",x"000000",x"332011",x"332011",x"311d10",x"352013",x"301d10",x"341f11",x"321e11",x"2d1b0e",x"181009",x"321b0b",x"564132",x"452916",x"3e2513",x"392212",x"331d10",x"3d2312",x"2b190b",x"926745",x"885f3f",x"8e6446",x"986b4b",x"9b6e4d",x"8a6042",x"916749",x"906649",x"906545",x"95694a",x"996e4e",x"8f6445",x"9a714f",x"976c4c",x"926749",x"986d4e",x"855e42",x"986e4f",x"936a4a",x"8f6546",x"936f4f",x"9d7151",x"895e41",x"906648",x"8f6647",x"906647",x"956848",x"976b4b",x"95694a",x"926747",x"895e3f",x"906647",x"93694b",x"986d4e",x"906446",x"8c6345",x"916748",x"9a704f",x"8e6446",x"704e36",x"7c583f",x"5d3f2a",x"4e3625",x"4e3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2210",x"3d2210",x"150e07",x"150e07",x"150e07",x"4d443a",x"4d443a",x"3e3228",x"50311d",x"50311d",x"331d0d",x"150e07",x"150e07",x"150e07",x"452612",x"3b200e",x"432712",x"432712",x"402511",x"3d220f",x"3e220f",x"3d210e",x"432510",x"391f0d",x"3a200e",x"211409",x"906749",x"855f42",x"936849",x"966d4d",x"936747",x"9b6e4e",x"976b4b",x"976946",x"8f6443",x"835a3c",x"966947",x"916643",x"906646",x"966948",x"8e6345",x"845c3e",x"936949",x"9e7352",x"916647",x"895f40",x"916749",x"946848",x"9f7554",x"906646",x"996e4e",x"986c4c",x"906547",x"986e4d",x"865e42",x"966a4a",x"916f4f",x"9d7251",x"875e41",x"8b6244",x"7d583f",x"755239",x"704e36",x"483221",x"473221",x"473221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543826",x"543826",x"452812",x"341c0c",x"3f2411",x"351d0d",x"391f0e",x"3e2310",x"412410",x"2f180a",x"371d0d",x"3d230f",x"432510",x"2c190b",x"170f07",x"150e07",x"160f08",x"160f08",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"25150a",x"2b190b",x"000000",x"341d0d",x"2d1a0b",x"150e07",x"150e07",x"311c0c",x"150e07",x"150e07",x"543521",x"37281d",x"51473d",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"150e07",x"150e07",x"150e07",x"191008",x"2f1d0f",x"33261d",x"453b32",x"453b32",x"000000",x"604430",x"604430",x"2f1a0b",x"201309",x"1d1108",x"190f07",x"1f1208",x"221409",x"150e07",x"28180b",x"25160a",x"28170a",x"2c190b",x"231409",x"201208",x"25150a",x"211409",x"23150a",x"26170b",x"26170b",x"22150a",x"26170b",x"28170b",x"28170b",x"1b1108",x"221409",x"28170b",x"231509",x"201309",x"27170a",x"211309",x"27160a",x"211309",x"251509",x"211309",x"231409",x"201208",x"1c1108",x"221409",x"201309",x"221409",x"231409",x"211309",x"1c1008",x"1c1008",x"1d1108",x"221409",x"231509",x"201309",x"221309",x"221309",x"211309",x"201309",x"1f1209",x"1b1008",x"1b1008",x"1d1108",x"472812",x"150e07",x"846041",x"856041",x"815d3f",x"835f41",x"845f41",x"846142",x"825e40",x"886444",x"886543",x"815e3f",x"835f3f",x"815d3e",x"7d5a3b",x"785639",x"7c593c",x"7e5d3e",x"7b593c",x"79573a",x"64442c",x"765639",x"7a593c",x"856143",x"836042",x"846244",x"7f5e41",x"825f41",x"856242",x"896645",x"8a6747",x"846041",x"825e40",x"876343",x"7a583c",x"7e5b3d",x"7f5b3d",x"825e41",x"7c593c",x"815f40",x"886341",x"886444",x"866343",x"845f40",x"886342",x"876241",x"845f3f",x"805c3c",x"866041",x"846141",x"825e40",x"825e3f",x"69462d",x"7f5d3f",x"886343",x"8b6646",x"8a6646",x"564436",x"564436",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"47382d",x"47382d",x"402410",x"381e0c",x"371e0d",x"3e230f",x"391f0d",x"381f0d",x"3f2410",x"38200e",x"3e2310",x"4a2a13",x"2a170a",x"231409",x"231409",x"313131",x"34302d",x"313131",x"333333",x"2b2b2b",x"5b5b5b",x"525252",x"333333",x"585858",x"505050",x"565656",x"5e5e5e",x"5c5c5c",x"606060",x"5c5c5c",x"414141",x"313131",x"4f4f4f",x"545454",x"5a5a5a",x"5a5a5a",x"535353",x"5c5b5b",x"5e5d5c",x"5f5f5f",x"616161",x"5e5d5c",x"626161",x"606060",x"666564",x"666464",x"636363",x"5e5e5e",x"5a5a5a",x"5c5c5c",x"5b5a59",x"5d5c5a",x"5a5a59",x"454545",x"323333",x"333333",x"2c2c2c",x"323232",x"333333",x"323232",x"343434",x"454442",x"54504c",x"5e5852",x"665f58",x"68615b",x"5b554f",x"55524e",x"484746",x"383838",x"545454",x"333333",x"313131",x"2b2b2b",x"313131",x"4b2912",x"28170a",x"261509",x"341c0b",x"331a0b",x"381e0d",x"3a210f",x"381e0d",x"3e2310",x"402511",x"3e2310",x"331a0b",x"4a2811",x"311b0c",x"351e0d",x"3e2410",x"39200e",x"351d0c",x"301a0b",x"150e07",x"361e0e",x"2c190b",x"150e07",x"341d0d",x"323232",x"313131",x"313131",x"313131",x"333333",x"323232",x"484848",x"313131",x"333333",x"545452",x"6f6963",x"605d5a",x"4e4a47",x"696561",x"5d5d5d",x"616161",x"323232",x"313131",x"353535",x"3e3e3d",x"464646",x"383838",x"5d564e",x"5d5650",x"65605a",x"5d5752",x"5f5954",x"6e6862",x"655e57",x"665f59",x"645d56",x"655e58",x"6b635c",x"625b54",x"605851",x"6e6760",x"69615a",x"675f58",x"5e564e",x"343434",x"323232",x"323232",x"462813",x"482913",x"442713",x"3b2210",x"482913",x"26160a",x"5e5044",x"25150a",x"4a2c15",x"3f2411",x"351d0d",x"39200e",x"351e0d",x"371e0d",x"150e07",x"311b0b",x"150e07",x"150e07",x"000000",x"000000",x"321f12",x"321f12",x"2d1b10",x"372111",x"362011",x"352011",x"2b1b0f",x"28190d",x"18110a",x"391f0d",x"543f32",x"442714",x"412615",x"3d2514",x"362011",x"3a2111",x"301c0d",x"855d3e",x"906443",x"886043",x"9a6d4c",x"9a6e4d",x"8f6445",x"9d704f",x"a07352",x"966a4b",x"996d4d",x"a37756",x"966b4a",x"a27755",x"95694a",x"906648",x"966a4a",x"946a4b",x"9e7453",x"946a4b",x"926748",x"946d4d",x"986c4c",x"8f6446",x"926749",x"7e583d",x"936849",x"966b4a",x"906444",x"986b4b",x"926646",x"946847",x"855d42",x"926748",x"916748",x"8c6344",x"996d4c",x"8e6447",x"92694a",x"866144",x"7b563c",x"825d42",x"543a26",x"503926",x"503926",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"331d0c",x"331d0c",x"150e07",x"150e07",x"150e07",x"4a4037",x"4a4037",x"3e332b",x"51311a",x"51311a",x"2b190b",x"150e07",x"150e07",x"150e07",x"462712",x"3b1f0d",x"472913",x"442813",x"402511",x"3e2310",x"351d0d",x"381f0d",x"41240f",x"381d0c",x"3a200e",x"1d1208",x"78533b",x"966e4e",x"926748",x"8e6547",x"8a6041",x"9d714e",x"9c7050",x"895f3f",x"986b48",x"865d3d",x"996c48",x"895f3f",x"966a4b",x"986b4b",x"906445",x"8c6243",x"8c6547",x"916a4d",x"825c3f",x"8d6345",x"976c4d",x"956b4b",x"976e4d",x"8b6142",x"976a4b",x"94694a",x"946849",x"996d4e",x"966b4b",x"835b3f",x"946949",x"926849",x"8c6344",x"91684a",x"875f42",x"80593f",x"704e35",x"442f1e",x"46301f",x"46301f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513623",x"513623",x"412511",x"351d0c",x"3d2210",x"361e0d",x"3c210f",x"412511",x"3e230f",x"361d0c",x"3a1f0d",x"3b200e",x"452611",x"311b0d",x"1c1008",x"1a0f08",x"171009",x"171009",x"000000",x"170f07",x"170f07",x"150e07",x"150e07",x"26160a",x"2a190b",x"000000",x"28170a",x"29180a",x"1c1108",x"150e07",x"2d1a0b",x"150e07",x"150e07",x"523423",x"37281d",x"564d43",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1d11",x"332319",x"3f352d",x"3f352d",x"000000",x"5a422f",x"5a422f",x"271609",x"1f1208",x"1f1309",x"1f1208",x"1c1008",x"1b1008",x"150e07",x"2d1a0c",x"27160a",x"2a190b",x"2d1a0c",x"2a190b",x"28170a",x"25160a",x"25150a",x"1e1208",x"25150a",x"201309",x"1d1208",x"27170a",x"221409",x"28170a",x"29170a",x"211309",x"25150a",x"231409",x"26160a",x"29170a",x"241509",x"27160a",x"28180b",x"1b1108",x"241509",x"26160a",x"24150a",x"27170a",x"1e1209",x"2a190b",x"28170b",x"201309",x"28170b",x"23150a",x"25160a",x"231409",x"27160a",x"2b190b",x"27170a",x"29180b",x"2d1a0c",x"231409",x"231409",x"211309",x"231509",x"1f1208",x"1f1309",x"442611",x"150e07",x"775437",x"705135",x"7b593b",x"6f4f33",x"815d3f",x"876343",x"876243",x"815e3f",x"866141",x"7d593b",x"835e3f",x"866142",x"845f40",x"7b593a",x"7c583a",x"7c5a3c",x"7e5b3d",x"846143",x"846244",x"7d5b3f",x"7c5b3c",x"805d3e",x"826041",x"7d593c",x"79573b",x"7d5a3c",x"7e5b3d",x"7d5b3d",x"825e3f",x"7b593b",x"775538",x"725136",x"6f4d33",x"755437",x"7c593b",x"765536",x"805c3e",x"866141",x"846041",x"805d3e",x"7f5b3d",x"7c593b",x"825e3e",x"876243",x"846040",x"815d3e",x"805b3c",x"866041",x"846040",x"8f6a49",x"8d6949",x"856243",x"896543",x"866142",x"896445",x"58463a",x"58463a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"322921",x"322921",x"3b210e",x"3e2310",x"361d0c",x"3f2310",x"381f0d",x"3b200e",x"3d220f",x"3d220f",x"3f2410",x"4a2a13",x"271609",x"231409",x"231409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"303030",x"323232",x"333333",x"2c2c2c",x"323232",x"505050",x"575756",x"545352",x"52514f",x"595756",x"51504f",x"514f4d",x"414141",x"4c4c4c",x"4f4f4f",x"606060",x"313131",x"323232",x"303030",x"333332",x"472711",x"27160a",x"27160a",x"321a0b",x"321a0b",x"331c0c",x"3c210f",x"2f1a0c",x"3a210f",x"3a210f",x"39200e",x"391f0d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a200e",x"2f1b0c",x"282828",x"2d2d2d",x"323232",x"343434",x"323232",x"2f2f2f",x"323232",x"323232",x"333333",x"4d4c4b",x"6f6862",x"4b4946",x"4b4642",x"5c5955",x"505050",x"4b4b4b",x"323232",x"323232",x"333333",x"393938",x"3d3d3c",x"3d3c3c",x"645d55",x"5c554f",x"5c5650",x"59534c",x"5a544f",x"67615b",x"665f5a",x"676059",x"68615a",x"635b53",x"5d554e",x"5f5750",x"625a52",x"625a52",x"5d554d",x"5f5750",x"605850",x"333333",x"333333",x"462812",x"462813",x"482913",x"442713",x"3c2310",x"462812",x"472913",x"4b2b14",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"301f13",x"301f13",x"362214",x"321e11",x"372011",x"2f1c10",x"321e11",x"301d0f",x"181009",x"351d0b",x"564235",x"3d2312",x"452a17",x"3c2312",x"382112",x"331e0f",x"24150a",x"704c33",x"80593b",x"966a4a",x"986b4b",x"966b4b",x"8c6041",x"a07555",x"9e7352",x"94694a",x"946949",x"a37656",x"996c4c",x"a27655",x"926747",x"916648",x"936849",x"926748",x"9e7251",x"966a4a",x"8a6043",x"8e694a",x"906648",x"885f41",x"8e6447",x"956a4b",x"926749",x"906647",x"8d6242",x"885f41",x"936747",x"8c6446",x"8b6143",x"92694b",x"8f6445",x"926749",x"956a4b",x"8e6546",x"80593f",x"8e6648",x"815a3f",x"7d5a3f",x"523825",x"4b3523",x"4b3523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a210f",x"3a210f",x"150e07",x"150e07",x"150e07",x"4c4239",x"4c4239",x"3a2f26",x"532f17",x"532f17",x"28160a",x"150e07",x"150e07",x"150e07",x"4f2d15",x"371d0d",x"442813",x"3e2410",x"402511",x"3a200e",x"351d0d",x"3a200d",x"3f230f",x"3c210e",x"371d0c",x"211409",x"896144",x"996e4d",x"8f6546",x"9d714f",x"875a3f",x"966a48",x"9a6f4e",x"8b6145",x"936745",x"906544",x"81593b",x"8f6442",x"986c4c",x"926646",x"8a6143",x"865d3f",x"926a4b",x"9e7555",x"8a6142",x"976b4b",x"966b4d",x"916747",x"a07454",x"885e41",x"926849",x"896043",x"8d6446",x"906648",x"936b4b",x"946949",x"936849",x"8e6445",x"8b6243",x"936a4b",x"8b6245",x"815b3f",x"6f4e34",x"46311f",x"473120",x"473120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2f1d",x"4b2f1d",x"442611",x"321b0c",x"3e2310",x"351d0d",x"3c210f",x"3b220f",x"3b200e",x"381f0d",x"381f0d",x"391f0e",x"3e220f",x"2d1a0b",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"36200f",x"150e07",x"150e07",x"150e07",x"2d1b0c",x"2e1a0c",x"000000",x"000000",x"1c1108",x"1c1108",x"150e07",x"2b190b",x"150e07",x"150e07",x"543522",x"36291f",x"554c41",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"150e07",x"150e07",x"150e07",x"150e07",x"291d13",x"322317",x"3b3229",x"3b3229",x"000000",x"5e4431",x"5e4431",x"2f1a0b",x"1c1108",x"150e07",x"201309",x"1f1208",x"1e1208",x"150e07",x"2c1a0c",x"25160a",x"29180b",x"27170a",x"2a180b",x"231509",x"26160a",x"211409",x"211409",x"241509",x"231509",x"26160a",x"26160b",x"1e1209",x"25160a",x"24150a",x"1e1208",x"1f1309",x"24150a",x"221409",x"231409",x"191008",x"29180b",x"26160a",x"26160a",x"25150a",x"2e1a0c",x"27160a",x"25150a",x"211309",x"201309",x"221409",x"231409",x"231509",x"211409",x"23150a",x"231509",x"27170b",x"25160a",x"27170a",x"27170b",x"2a180b",x"26160a",x"26160a",x"1f1208",x"211409",x"1d1108",x"1d1108",x"442712",x"150e07",x"846041",x"7b593c",x"7c593c",x"7f5b3d",x"856141",x"886545",x"8b6646",x"825f41",x"886444",x"826040",x"815e3f",x"8c6746",x"866242",x"815e3e",x"7e5b3d",x"735337",x"755537",x"765538",x"825e41",x"7d5b3d",x"75553a",x"745437",x"58381d",x"745437",x"725236",x"775639",x"77563a",x"7a593b",x"7e5b3d",x"7e5b3d",x"805d40",x"7a593c",x"805d3e",x"7e5c3e",x"7e5b3e",x"815d3e",x"866242",x"886444",x"876343",x"825f41",x"856242",x"825e40",x"815d3f",x"8a6645",x"815e3f",x"876241",x"825d3f",x"7b593b",x"7f5c3c",x"835f40",x"896344",x"856141",x"7f5c3f",x"7c593b",x"613e20",x"4f4237",x"4f4237",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"412d1e",x"412d1e",x"361e0d",x"412611",x"3a200d",x"3f2410",x"39200e",x"3c220f",x"3a200e",x"391f0e",x"432712",x"452611",x"2c190b",x"221409",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"303030",x"323232",x"333333",x"2c2c2c",x"323232",x"505050",x"575756",x"545352",x"52514f",x"595756",x"51504f",x"514f4d",x"414141",x"4c4c4c",x"4f4f4f",x"606060",x"313131",x"323232",x"303030",x"442c1d",x"4f2c13",x"26160a",x"2d190b",x"351d0c",x"331a0b",x"39200e",x"3b210f",x"3a200e",x"331d0e",x"371f0e",x"3d220f",x"402410",x"59341a",x"432713",x"311c0d",x"432713",x"462a14",x"3d2411",x"150e07",x"37200f",x"3d2411",x"452914",x"422612",x"4a2d16",x"462813",x"4a2b15",x"4a2b15",x"4c2d16",x"482913",x"432511",x"422511",x"462712",x"482813",x"472813",x"452712",x"412511",x"452611",x"452612",x"442611",x"462812",x"412611",x"492a14",x"452712",x"3e220f",x"462812",x"4c2d15",x"492b15",x"452813",x"452713",x"442713",x"462813",x"482a14",x"492a14",x"492a14",x"482b14",x"4a2c15",x"492b15",x"472a15",x"452814",x"402511",x"442813",x"462914",x"412511",x"3d220f",x"3e2310",x"3b210f",x"442813",x"432712",x"412511",x"462813",x"3c210f",x"3b210f",x"3b210f",x"3a200e",x"3b210f",x"331d0d",x"422511",x"3f2411",x"402511",x"3c2310",x"27160a",x"3d2410",x"150e07",x"150e07",x"000000",x"000000",x"2f1e12",x"2f1e12",x"342013",x"2f1c10",x"352011",x"331e11",x"321e11",x"29190d",x"181009",x"311b0b",x"524135",x"4a2a15",x"3e2413",x"402615",x"3a2313",x"382110",x"2f1b0d",x"845c3d",x"674733",x"996d4d",x"966a4a",x"8e6444",x"8e6243",x"8d6345",x"a17554",x"966b4b",x"926648",x"a07453",x"986c4c",x"a37857",x"95694a",x"996c4b",x"8c6345",x"906647",x"956b4c",x"986e4f",x"825b40",x"9d7554",x"8d6345",x"8e6547",x"875e42",x"825b40",x"8d6445",x"956949",x"835b3f",x"704c33",x"946848",x"946849",x"8b6243",x"946a49",x"906548",x"93684a",x"835c40",x"916747",x"926646",x"906749",x"855d42",x"7f5a40",x"452d1c",x"4d3625",x"4d3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381e0d",x"381e0d",x"150e07",x"150e07",x"150e07",x"473f35",x"473f35",x"3c3128",x"4b2d19",x"4b2d19",x"331c0c",x"150e07",x"150e07",x"150e07",x"502e16",x"3b210e",x"3f2511",x"3e2411",x"3f2410",x"3b200e",x"381f0e",x"3b210f",x"3c230f",x"3b200e",x"361d0c",x"1b1108",x"8a6346",x"966d4d",x"8d6344",x"986d4c",x"774d33",x"9b6e4c",x"986d4d",x"926546",x"95694a",x"8b6141",x"855d3d",x"986d4d",x"976b4b",x"8d6447",x"8b6245",x"8b6344",x"9e7252",x"9b6f51",x"8e6447",x"80593e",x"8e6547",x"936949",x"a07554",x"8d6446",x"9a6e4d",x"8d6346",x"8f6445",x"9d7251",x"936849",x"906445",x"9a6f4f",x"8b6143",x"8d6346",x"6c4b34",x"845d41",x"7f5a3e",x"6d4c34",x"432e1e",x"462f1f",x"462f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462916",x"462916",x"40230f",x"361e0d",x"3f2410",x"39200e",x"3b210f",x"402410",x"3a200e",x"3a200d",x"3a200e",x"3b200e",x"442511",x"2f1a0c",x"150e07",x"27160a",x"150e07",x"150e07",x"000000",x"351e0d",x"351e0d",x"231509",x"221409",x"2e1a0c",x"2e1a0c",x"000000",x"000000",x"170f07",x"170f07",x"150e07",x"2d1a0b",x"180f07",x"150e07",x"503320",x"3a291f",x"584e43",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1d14",x"2f2015",x"383028",x"383028",x"000000",x"554233",x"554233",x"2e190a",x"1e1208",x"1e1209",x"1e1208",x"1e1208",x"1d1108",x"150e07",x"28170a",x"2a180b",x"2a180b",x"2d1a0c",x"27170a",x"28170a",x"26160a",x"25160a",x"26160a",x"28180b",x"25160a",x"26170b",x"26160a",x"211409",x"29180b",x"2a1a0c",x"24160a",x"24160a",x"26170b",x"24150a",x"27180b",x"221409",x"24160a",x"1e1208",x"311c0d",x"25160a",x"28180b",x"23150a",x"221409",x"231409",x"201309",x"201309",x"1f1209",x"1f1309",x"231409",x"211409",x"211409",x"26160a",x"25160a",x"24150a",x"27170a",x"27160a",x"25150a",x"150e07",x"1d1108",x"25150a",x"1c1108",x"1d1108",x"452812",x"150e07",x"896544",x"835f40",x"7f5c3d",x"815e3f",x"846142",x"8b6748",x"8e6949",x"8b6647",x"906b4a",x"8e6a4a",x"8e6949",x"886546",x"856241",x"815c3e",x"876243",x"8b6647",x"876445",x"815e41",x"805e3f",x"805e40",x"7e5c3f",x"816040",x"7d5a3c",x"7d5b3e",x"7a583b",x"795739",x"7c593c",x"815e40",x"825e3f",x"825d3f",x"805c3e",x"835f3f",x"846141",x"7f5c3e",x"7e5c3d",x"805e3e",x"745539",x"926c4b",x"8d6949",x"896646",x"8f6a49",x"8b6748",x"8d6849",x"886546",x"846141",x"866041",x"8c6646",x"906a4a",x"805e41",x"906a48",x"8c6646",x"886445",x"876343",x"8a6544",x"886342",x"57473a",x"57473a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"372418",x"372418",x"3a200e",x"3e2411",x"3d2310",x"3d2310",x"3e2310",x"381f0e",x"381f0d",x"3b210e",x"3c2310",x"4a2a13",x"2b1a0c",x"201208",x"201208",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"43250f",x"381f0c",x"4e392b",x"4e2b12",x"29180b",x"2a180b",x"391f0d",x"331b0b",x"3b200e",x"3b210f",x"3c210f",x"37200f",x"3e2310",x"3d2310",x"3e220f",x"553119",x"442813",x"3e2411",x"472914",x"452914",x"412511",x"351d0d",x"341d0d",x"381f0e",x"432712",x"432713",x"442713",x"3c210f",x"3c210f",x"3e220f",x"3c210f",x"3d210f",x"3d210f",x"3a200e",x"381f0d",x"381e0d",x"3b200e",x"391e0d",x"3b200e",x"3b200e",x"3b200f",x"3a200f",x"3a200f",x"3f230f",x"3d220f",x"3e2310",x"3f2511",x"432712",x"462813",x"402511",x"402511",x"3e2411",x"3e2411",x"3f2411",x"39200e",x"3f2512",x"422613",x"442813",x"3f2410",x"402411",x"432612",x"412612",x"412512",x"3f2511",x"422713",x"3f2310",x"3c210e",x"3a210f",x"381f0e",x"351d0d",x"3a210f",x"412511",x"3b210f",x"3d2310",x"3f2410",x"432612",x"39200e",x"412612",x"371f0e",x"402411",x"39200e",x"361f0e",x"39200f",x"211409",x"371f0e",x"150e07",x"150e07",x"000000",x"000000",x"2f1d12",x"2f1d12",x"352114",x"301e12",x"341f11",x"341f11",x"2d1b0f",x"29190e",x"181009",x"391f0d",x"524338",x"452714",x"3c2312",x"3b2312",x"3d2312",x"3f2513",x"321d0e",x"835d43",x"9a7050",x"906647",x"9a6d4d",x"936747",x"916648",x"a37654",x"a37856",x"9c6f50",x"936748",x"956b4c",x"966c4d",x"9e7452",x"986c4c",x"976b4b",x"9b7150",x"8f6547",x"93694a",x"966c4c",x"916748",x"946d4f",x"916748",x"8e6447",x"9b6f4f",x"8d6446",x"906646",x"986d4d",x"845c3e",x"8d6343",x"906445",x"6d4933",x"966b4b",x"906547",x"8f6547",x"976b4c",x"8a6143",x"8d6445",x"7d563b",x"906748",x"7e573d",x"7b573d",x"5a3d29",x"4b3423",x"4b3423",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"391f0e",x"391f0e",x"150e07",x"150e07",x"150e07",x"463e35",x"463e35",x"3c3128",x"4c2f1d",x"4c2f1d",x"311b0c",x"150e07",x"150e07",x"150e07",x"472712",x"402411",x"3d2410",x"3e2410",x"3c210f",x"3c210f",x"3d220f",x"402510",x"3d2310",x"3a210e",x"331b0b",x"201309",x"8a6344",x"8e6647",x"8d6344",x"986b4b",x"7f5639",x"966b4a",x"95694a",x"906545",x"8f6546",x"906647",x"976c4c",x"916648",x"94694a",x"9b7051",x"8d6344",x"896043",x"926748",x"8e6649",x"916749",x"926849",x"916748",x"946a4b",x"956c4c",x"956a4a",x"996f4d",x"996e4f",x"946849",x"996e4e",x"906646",x"8f6648",x"9b7251",x"906648",x"8b6346",x"91684b",x"825b3e",x"7b573c",x"6e4e36",x"402b1c",x"402b1c",x"402b1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472916",x"472916",x"402310",x"321b0b",x"412611",x"371e0d",x"3b210f",x"3f2410",x"3b210e",x"371e0c",x"3d220f",x"3b200e",x"452611",x"321c0d",x"2b190b",x"2b190b",x"150e07",x"150e07",x"000000",x"351e0d",x"351e0d",x"231509",x"25150a",x"2e1a0c",x"2e1a0c",x"000000",x"000000",x"1e1208",x"191008",x"150e07",x"150e07",x"1b1008",x"150e07",x"543623",x"38291f",x"574d43",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1e14",x"2d2017",x"382e26",x"382e26",x"000000",x"584538",x"584538",x"2f1a0a",x"1f1208",x"201308",x"170f07",x"1e1208",x"211309",x"150e07",x"24160a",x"27170b",x"29180b",x"29170b",x"2c190c",x"241509",x"241509",x"231409",x"221409",x"24150a",x"28170b",x"2d1a0c",x"1d1209",x"1e1209",x"1d1209",x"1f1309",x"2b190b",x"1e1208",x"201309",x"221409",x"2b190b",x"211409",x"27170b",x"27160a",x"251509",x"201309",x"1d1108",x"251509",x"231509",x"201309",x"211309",x"1f1208",x"191008",x"201208",x"1d1108",x"1e1208",x"211409",x"1c1108",x"211309",x"1e1208",x"1f1208",x"25150a",x"25150a",x"1d1108",x"190f08",x"1c1108",x"1d1108",x"150e07",x"4d2c15",x"150e07",x"7c5a3b",x"775337",x"7c5b3b",x"765436",x"7f5c3e",x"805d40",x"805d3e",x"8b6746",x"886344",x"886344",x"836041",x"836043",x"835f41",x"856142",x"836041",x"815e40",x"805e3f",x"7b593c",x"815e40",x"815e40",x"7e5c3d",x"7a583b",x"7a593b",x"7a593c",x"815e3f",x"79573b",x"7a593a",x"7a583c",x"815c3f",x"855f41",x"815d3f",x"79583a",x"79583a",x"775537",x"7a593a",x"775537",x"775639",x"835f41",x"7f5d3e",x"866243",x"856243",x"886344",x"886444",x"906a4a",x"896444",x"8a6545",x"866243",x"8c6646",x"8a6445",x"866142",x"846042",x"8a6645",x"876242",x"815d3f",x"846041",x"5a473a",x"5a473a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3f291a",x"3f291a",x"3d220f",x"402512",x"3e2310",x"3e2310",x"3c210f",x"3b210f",x"3a200e",x"3c210f",x"3e230f",x"422510",x"24150a",x"3a1e0c",x"3d210f",x"28170a",x"3f2310",x"442611",x"492913",x"442510",x"432510",x"40230f",x"3f230e",x"452711",x"432610",x"4f2d15",x"4d2d16",x"4c2c16",x"4e2d16",x"4b2b14",x"4c2d15",x"543117",x"4a2a14",x"4b2b14",x"4e2d15",x"492913",x"452711",x"472712",x"482812",x"452712",x"442611",x"3f220f",x"3e220f",x"41240f",x"422510",x"3f230f",x"442610",x"462711",x"452711",x"452710",x"472811",x"472811",x"432510",x"4a2a14",x"4a2a14",x"4b2b14",x"4a2a14",x"462711",x"452611",x"462711",x"472712",x"422410",x"442511",x"422510",x"442611",x"472812",x"462812",x"462812",x"442712",x"432611",x"3f2410",x"3f220f",x"3e220e",x"452610",x"533118",x"4d2a13",x"1f1309",x"211409",x"391f0d",x"331c0c",x"3d210e",x"3a200e",x"3f230f",x"432812",x"462913",x"371f0d",x"3c210f",x"512f16",x"38210f",x"452914",x"3f2612",x"3f2411",x"422612",x"3a2310",x"1e1309",x"442914",x"442813",x"452813",x"432712",x"472a14",x"442712",x"432611",x"3e220f",x"3e220f",x"3d2310",x"3d2310",x"3f220f",x"3f230f",x"432611",x"412511",x"432611",x"402411",x"432611",x"3f2310",x"3f2410",x"3d220f",x"432611",x"472913",x"422612",x"3e220f",x"3d220f",x"3e2411",x"412411",x"3c210f",x"3f2411",x"3b220f",x"3f2410",x"3c2210",x"3d2310",x"412410",x"3f230f",x"381f0d",x"381e0d",x"281307",x"351c0c",x"391f0e",x"3b210e",x"391f0e",x"3c210f",x"3d210f",x"3a200f",x"3b210f",x"3d220f",x"3d2210",x"3f2410",x"3e2310",x"422611",x"402511",x"422611",x"3f2511",x"412612",x"3d2410",x"37200f",x"39210f",x"321d0d",x"150e07",x"341d0d",x"150e07",x"150e07",x"000000",x"000000",x"311e12",x"311e12",x"342013",x"311f12",x"351f11",x"342011",x"2f1d10",x"28190e",x"18110a",x"3a200d",x"534235",x"3f2513",x"362011",x"412715",x"341f11",x"3e2412",x"28180b",x"5f412e",x"9c7151",x"986d4d",x"976b4b",x"8f6545",x"9b7050",x"a27654",x"9c7050",x"986c4d",x"926749",x"9b6f4e",x"936849",x"a07454",x"976c4b",x"8e6345",x"9c7151",x"986c4d",x"966c4d",x"936949",x"8d6446",x"976d4d",x"7a553d",x"906547",x"825b41",x"906546",x"946949",x"9c6f4f",x"8c6142",x"926647",x"8c6143",x"966949",x"956a4a",x"986b4b",x"7d573b",x"966b4c",x"896042",x"885f43",x"8b6245",x"896144",x"7e5a3d",x"725036",x"553a27",x"4b3323",x"4b3323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"331d0d",x"331d0d",x"150e07",x"150e07",x"150e07",x"423a31",x"423a31",x"3d3128",x"462916",x"462916",x"29170a",x"150e07",x"150e07",x"150e07",x"432612",x"442813",x"412611",x"3a210f",x"3e2310",x"3b210f",x"3b210e",x"422611",x"3f2410",x"371f0d",x"341c0b",x"1d1108",x"90674b",x"906748",x"8c6143",x"916645",x"8a5d3f",x"966a4a",x"9c6f50",x"8a6041",x"8a6143",x"845a3e",x"a07352",x"95694a",x"9e7151",x"93694a",x"8c6345",x"876043",x"8e6648",x"986f50",x"8d6448",x"946a4a",x"946949",x"986d4d",x"946b4b",x"906547",x"9a6d4c",x"976d4d",x"956b4b",x"986c4c",x"966a4a",x"8d6546",x"9d7554",x"906648",x"8a6144",x"8f6649",x"845d41",x"775339",x"6f4d35",x"442e1d",x"432e1d",x"432e1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472815",x"472815",x"402410",x"311a0b",x"371f0e",x"361e0d",x"412511",x"412511",x"3d220f",x"361e0c",x"3e220f",x"391f0d",x"4a2913",x"2b180a",x"2f1b0c",x"2f1b0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"170e07",x"1f1208",x"150e07",x"5a3a24",x"392a1f",x"554b40",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"150e07",x"1d1108",x"2f2016",x"302219",x"342b23",x"342b23",x"000000",x"523e30",x"523e30",x"301a0b",x"170f07",x"1c1108",x"1d1108",x"201309",x"1a1008",x"150e07",x"26160a",x"27170b",x"301d0d",x"2c1a0c",x"2c1a0c",x"2a190b",x"2c190c",x"26160a",x"25160a",x"27170b",x"27170b",x"29180b",x"211409",x"24160a",x"25160a",x"26160a",x"26160a",x"2b190c",x"29180b",x"2a190c",x"29190b",x"27170b",x"27170b",x"27170b",x"28170b",x"24150a",x"251509",x"1c1108",x"211309",x"1f1309",x"1e1208",x"211309",x"190f08",x"26160a",x"26160a",x"231509",x"1c1108",x"211409",x"241509",x"1f1209",x"231509",x"27170b",x"211309",x"24150a",x"150e07",x"1c1108",x"1e1208",x"201309",x"402410",x"150e07",x"785639",x"7b593b",x"795538",x"765436",x"7d5b3b",x"7c593c",x"7f5c3e",x"835f41",x"805e40",x"7d5a3d",x"815d3f",x"7c593c",x"7e5c3e",x"846042",x"836143",x"876445",x"856142",x"7d5b3e",x"7a593c",x"755437",x"7a583b",x"765638",x"7c5b3c",x"815e40",x"775538",x"805d3e",x"825f41",x"78573a",x"7b593a",x"7a583a",x"79583a",x"805d3d",x"755438",x"7b583b",x"765336",x"775637",x"745436",x"7c593c",x"7b593c",x"805c3f",x"825f41",x"7f5b3e",x"815d3f",x"805c3e",x"846041",x"896545",x"8e6949",x"916c4b",x"8c6746",x"846140",x"815d3f",x"6b4d32",x"815e3f",x"7d5b3c",x"825f3f",x"57473a",x"57473a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"342418",x"342418",x"3b200e",x"3c210f",x"38200e",x"3b210e",x"3b200e",x"39200e",x"3a200e",x"3b200e",x"3d210e",x"371e0d",x"3a200d",x"3c210e",x"3c200e",x"2c190b",x"3f2310",x"442611",x"492913",x"442510",x"432510",x"40230f",x"3f230e",x"452711",x"432610",x"4f2d15",x"4d2d16",x"4c2c16",x"4e2d16",x"4b2b14",x"4c2d15",x"543117",x"4a2a14",x"4b2b14",x"4e2d15",x"492913",x"452711",x"472712",x"482812",x"452712",x"442611",x"3f220f",x"3e220f",x"41240f",x"422510",x"3f230f",x"442610",x"462711",x"452711",x"452710",x"472811",x"472811",x"432510",x"4a2a14",x"4a2a14",x"4b2b14",x"4a2a14",x"462711",x"452611",x"462711",x"472712",x"422410",x"442511",x"422510",x"442611",x"472812",x"462812",x"462812",x"442712",x"432611",x"3f2410",x"402310",x"40230f",x"4a2b15",x"4a2b15",x"462913",x"462913",x"482a14",x"462914",x"4a2c15",x"422612",x"432711",x"432711",x"3c220f",x"422611",x"442812",x"472a14",x"563419",x"442813",x"442814",x"150e07",x"3a2210",x"1f1309",x"150e07",x"150e07",x"38200f",x"3b220f",x"3e220f",x"402411",x"402410",x"3d220f",x"3d220f",x"3c210f",x"3f2410",x"3c220f",x"3c200e",x"432611",x"422510",x"3f230f",x"3e220f",x"3c210e",x"39200d",x"3b200e",x"3a1f0d",x"3b200e",x"391f0d",x"381f0d",x"361d0c",x"3c200e",x"3d210e",x"3a200e",x"3c210f",x"3c210f",x"3b210e",x"3d220f",x"3e2310",x"3e230f",x"371e0d",x"381e0d",x"3a1f0d",x"3f2410",x"452712",x"3b210f",x"381f0d",x"381f0d",x"3c220f",x"412511",x"3c210f",x"3c220f",x"3c220f",x"3a210f",x"3a210e",x"3e230f",x"3f2410",x"3e220f",x"3f2410",x"412511",x"412511",x"432612",x"412511",x"3f2511",x"150e07",x"29170a",x"2d190b",x"150e07",x"150e07",x"331d0d",x"150e07",x"150e07",x"000000",x"000000",x"301e13",x"301e13",x"342013",x"362113",x"362011",x"321e11",x"321e11",x"28190e",x"17110a",x"351d0c",x"574538",x"3a2312",x"351f10",x"3f2615",x"382212",x"3a2112",x"321d0e",x"90674a",x"845f46",x"9d7151",x"94694a",x"9c7050",x"9a6f50",x"815b41",x"9f7252",x"986d4e",x"95694a",x"96694b",x"956a4b",x"a07453",x"93694b",x"8c6244",x"9a6f4f",x"906647",x"916647",x"906647",x"986e4f",x"845d43",x"976c4e",x"8e6344",x"886145",x"895f42",x"815b3f",x"926747",x"7f563b",x"8f6446",x"8e6443",x"8f6646",x"8f6444",x"966c4b",x"8f6446",x"9b7050",x"835c41",x"855d41",x"926a4b",x"896041",x"7e593d",x"745138",x"533a26",x"4c3624",x"4c3624",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0c",x"311c0c",x"150e07",x"150e07",x"150e07",x"3f372e",x"3f372e",x"3b3027",x"4a2b17",x"4a2b17",x"2a180b",x"150e07",x"150e07",x"150e07",x"512e16",x"472a14",x"3d220f",x"3c210f",x"3d2311",x"3a210f",x"39200e",x"432611",x"412511",x"3b200e",x"2e180a",x"1c1108",x"8d6648",x"8b6143",x"8a6041",x"8f6546",x"8a6041",x"875e40",x"8f6445",x"8b6142",x"8b6143",x"885e3f",x"936849",x"855d42",x"815c41",x"936a4a",x"755138",x"996e4e",x"956b4d",x"936a4d",x"93694b",x"92694a",x"916747",x"9e7352",x"976d4d",x"94694a",x"7f593f",x"946b4c",x"8c6547",x"9b6f4e",x"9d7251",x"8c6244",x"a17757",x"91674a",x"885f43",x"8b6447",x"80593d",x"79543a",x"65452e",x"422d1c",x"432d1d",x"432d1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492a15",x"492a15",x"462812",x"361d0d",x"3a200e",x"3a200e",x"402511",x"3e230f",x"381e0d",x"3a200e",x"39200e",x"3f230f",x"3c210e",x"2c180a",x"351f0e",x"351f0e",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"27160a",x"27160a",x"150e07",x"23150a",x"150e07",x"150e07",x"563823",x"392b21",x"595045",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"1c1108",x"312117",x"332319",x"352b22",x"352b22",x"000000",x"543e31",x"543e31",x"321c0b",x"1f1208",x"1f1208",x"211409",x"231409",x"1d1208",x"150e07",x"23150a",x"26160a",x"2f1c0d",x"29180b",x"2c1a0c",x"211409",x"24150a",x"25160a",x"27170a",x"29180b",x"26170b",x"29180b",x"23150a",x"27170b",x"24160a",x"29180b",x"27170b",x"211409",x"26170a",x"28170b",x"24150a",x"25160a",x"25150a",x"25160a",x"211409",x"221409",x"1f1209",x"1d1108",x"201309",x"1f1208",x"201309",x"231409",x"150e07",x"211309",x"211309",x"211309",x"211309",x"1d1108",x"201308",x"1f1208",x"1f1208",x"201208",x"150e07",x"1b1108",x"191008",x"1a1008",x"150e07",x"1d1108",x"412410",x"150e07",x"856043",x"805d3f",x"805d3f",x"7e5a3d",x"7b593c",x"7e5b3e",x"775639",x"7d5a3d",x"815e41",x"805f41",x"805d3e",x"825f41",x"866443",x"886546",x"856242",x"826041",x"815d3f",x"765538",x"705033",x"755537",x"7c5a3b",x"815e40",x"7e5c3e",x"815c3e",x"815e41",x"866143",x"866343",x"856242",x"7d5b3e",x"825e3f",x"755536",x"7d5a3d",x"846142",x"805d3e",x"7f5b3e",x"7c593c",x"7c593b",x"7e5b3e",x"775639",x"7e5b3e",x"815f41",x"825f42",x"7d5b3d",x"866243",x"8a6745",x"886546",x"896544",x"886545",x"896343",x"7d5b3c",x"775637",x"7c5a3a",x"835f40",x"846142",x"805d3f",x"484037",x"484037",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"32251b",x"32251b",x"3c200d",x"3a200d",x"381e0d",x"351c0c",x"341c0c",x"341c0b",x"341c0c",x"341c0b",x"341c0b",x"361d0c",x"361d0c",x"371e0c",x"381e0d",x"3c210e",x"391f0e",x"361e0d",x"301a0b",x"331b0b",x"391f0d",x"3a200e",x"3f2411",x"3e2411",x"391f0e",x"3f2410",x"3a200f",x"3b200e",x"412612",x"472a14",x"402612",x"432713",x"452813",x"472a14",x"462914",x"442712",x"3a200e",x"3c220f",x"412612",x"442813",x"412712",x"402512",x"3d2310",x"3e2310",x"3e2411",x"412611",x"3d2410",x"3f2511",x"3a210f",x"3c2310",x"402511",x"3b2210",x"3d2411",x"3b2311",x"3f2512",x"412612",x"442813",x"3e2411",x"3a2210",x"3d2311",x"3e2310",x"442712",x"3f2411",x"3c210f",x"3b210f",x"412511",x"412511",x"3c220f",x"361e0e",x"402410",x"412511",x"412511",x"402511",x"432712",x"412511",x"412411",x"3e230f",x"3f2410",x"412510",x"3f240f",x"3f2510",x"432812",x"4b2c15",x"462913",x"422712",x"412612",x"462913",x"4f2d15",x"38200f",x"3b210f",x"321c0c",x"311c0c",x"29170a",x"2e1a0b",x"150e07",x"301b0c",x"371f0e",x"3b210f",x"39200e",x"3e2310",x"3c220f",x"3e2310",x"3e2310",x"3c210f",x"391f0e",x"391e0d",x"361d0d",x"371d0c",x"371d0c",x"371d0c",x"351c0c",x"341c0b",x"371d0c",x"361d0c",x"361d0c",x"361d0c",x"391e0d",x"3a200d",x"3a200e",x"39200e",x"381e0d",x"361d0c",x"381e0d",x"3a200e",x"3e2310",x"472813",x"412511",x"3d220f",x"402410",x"3c210f",x"462813",x"4b2c15",x"4b2c16",x"492b15",x"432713",x"482a15",x"462914",x"432713",x"3e220f",x"3d210f",x"432713",x"442813",x"492b15",x"452813",x"412511",x"422611",x"412612",x"402511",x"412511",x"412511",x"3d2310",x"361f0f",x"341e0e",x"331d0e",x"2b190b",x"150e07",x"341f0f",x"150e07",x"150e07",x"000000",x"000000",x"311f12",x"311f12",x"352114",x"382114",x"362012",x"2d1c0f",x"2c1b0f",x"27180d",x"181009",x"361e0c",x"544134",x"3a2211",x"372011",x"3d2514",x"392113",x"382112",x"27170b",x"946a4a",x"7a573e",x"986e4f",x"926849",x"966c4d",x"9a6d4c",x"74513a",x"a47957",x"9a6e4e",x"986c4c",x"986b4b",x"996d4d",x"9f7353",x"9e7353",x"956a4b",x"986e4e",x"926749",x"996d4e",x"996e4d",x"93694a",x"a17555",x"9f7352",x"93684a",x"865f44",x"956a4b",x"593928",x"996c4b",x"8e6345",x"8d6343",x"926646",x"845c3f",x"906747",x"896043",x"8c6344",x"8f6749",x"926749",x"7f593d",x"8f6748",x"855d41",x"765137",x"714e36",x"5e422d",x"503827",x"503827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"3d230f",x"150e07",x"150e07",x"150e07",x"403830",x"403830",x"352c23",x"4e2d18",x"4e2d18",x"301a0b",x"150e07",x"150e07",x"150e07",x"4c2a14",x"432612",x"432612",x"3b200e",x"412512",x"3b2210",x"3d230f",x"412611",x"462913",x"3b210e",x"341b0b",x"1f1208",x"876044",x"8e6647",x"845c3f",x"906647",x"896043",x"906546",x"94694a",x"936849",x"8e6345",x"875d3f",x"906747",x"916748",x"8b6447",x"8b6345",x"906648",x"966d4d",x"9a7050",x"90674a",x"8d6649",x"93694a",x"926648",x"996e4e",x"906748",x"976a4b",x"8c6345",x"986c4c",x"996e4e",x"976c4c",x"946949",x"996e4d",x"a07957",x"805b40",x"8b6145",x"90684a",x"7f5a3d",x"78543a",x"6b4a32",x"45301f",x"45301f",x"45301f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482915",x"482915",x"462812",x"3b200e",x"3c220f",x"3c220f",x"3c210f",x"3e230f",x"351d0c",x"3c210f",x"3a200d",x"3b200e",x"391e0c",x"271509",x"2f1b0b",x"2f1b0b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b190b",x"2b190b",x"150e07",x"221409",x"2b180a",x"150e07",x"55351f",x"312319",x"584e44",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"191008",x"372519",x"332317",x"312921",x"312921",x"000000",x"543e2f",x"543e2f",x"311b0b",x"251509",x"1e1208",x"1e1209",x"1f1208",x"27170a",x"150e07",x"25160a",x"27160a",x"26160a",x"2b180b",x"2c190b",x"2f1c0d",x"2d1a0c",x"24160a",x"28180b",x"24150a",x"28180b",x"27170a",x"26160a",x"25160a",x"27160a",x"25160a",x"26160a",x"241509",x"251609",x"211409",x"231509",x"24150a",x"241509",x"25150a",x"231509",x"26160a",x"27160a",x"1f1208",x"211309",x"1c1108",x"1d1108",x"1d1108",x"1a1008",x"1b1008",x"1e1208",x"170f07",x"231409",x"211308",x"1e1108",x"1a1008",x"150e07",x"1c1108",x"201309",x"1b1108",x"1a1008",x"150e07",x"191008",x"1a1008",x"412410",x"150e07",x"805d3f",x"866142",x"77563a",x"7b583b",x"7b593b",x"7d5a3c",x"856243",x"815d3e",x"886444",x"805c3e",x"7a5839",x"775337",x"835e3f",x"846041",x"805d3f",x"7a593b",x"7b5a3c",x"815d3f",x"7f5c3e",x"7e5c3e",x"805e3f",x"856242",x"856243",x"8a6747",x"866343",x"7f5b3e",x"825e3f",x"856141",x"7d5b3d",x"7b5a3b",x"7e5a3a",x"7d5a3b",x"7b593c",x"79583a",x"7c5a3c",x"7d5a3c",x"7d5a3c",x"735237",x"7f5d3f",x"7f5c3d",x"876343",x"815d3f",x"7d5a3b",x"705033",x"835f3f",x"876343",x"876343",x"7f5c3e",x"856141",x"825e3f",x"876342",x"825f41",x"826040",x"876343",x"896544",x"4c3a2d",x"4c3a2d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452f20",x"452f20",x"3e220f",x"3e220f",x"351d0c",x"351d0c",x"371d0c",x"371e0c",x"381e0c",x"331c0b",x"361d0d",x"371e0d",x"3a200e",x"3a1f0d",x"3a200d",x"391f0d",x"3c210f",x"3c220f",x"3c230f",x"361e0d",x"3d220f",x"371e0d",x"361d0c",x"3b210e",x"371f0e",x"341d0d",x"311c0c",x"351d0d",x"391f0d",x"391f0e",x"351e0d",x"321b0b",x"311a0b",x"351d0d",x"3e2411",x"39200e",x"331c0c",x"311b0b",x"321c0c",x"371f0d",x"341c0d",x"341d0c",x"321c0c",x"361e0e",x"3e2411",x"3a2210",x"3a2210",x"39210f",x"371f0e",x"331c0d",x"2e1a0b",x"39200f",x"38200e",x"2f1b0c",x"351e0e",x"371f0e",x"3e2311",x"3c2311",x"331d0e",x"38200f",x"39200f",x"3b220f",x"39200e",x"432713",x"432712",x"442813",x"462914",x"3e2511",x"36200f",x"3e2411",x"422713",x"432813",x"492b15",x"492b15",x"462914",x"462a14",x"432713",x"442713",x"452913",x"472913",x"452813",x"402512",x"442713",x"442713",x"3e2310",x"432712",x"4d2d16",x"5a351b",x"402612",x"3e2511",x"331d0d",x"150e07",x"150e07",x"2f1b0c",x"150e07",x"311c0d",x"3c220f",x"39200e",x"3c220f",x"3f2410",x"3b210f",x"3f240f",x"3b210f",x"391f0d",x"381f0d",x"3b200e",x"381f0d",x"3a200e",x"381f0c",x"351d0c",x"331b0b",x"341c0b",x"371e0d",x"391f0d",x"3a1f0d",x"3c210e",x"3b200e",x"3a200e",x"3f220f",x"422510",x"422611",x"3e230f",x"3c220f",x"3e220f",x"3a200d",x"3e220f",x"3f230f",x"3d220f",x"3d220f",x"3b210f",x"3e230f",x"3d210f",x"3c210e",x"3a1f0d",x"361d0c",x"371e0d",x"432611",x"462813",x"381e0d",x"361d0c",x"351d0c",x"3c210f",x"3f220f",x"361e0d",x"391f0d",x"412411",x"412511",x"402511",x"412511",x"3d2410",x"3b2210",x"371f0e",x"150e07",x"150e07",x"29180b",x"150e07",x"341d0d",x"150e07",x"150e07",x"000000",x"000000",x"322013",x"322013",x"332013",x"342013",x"2f1c10",x"341f10",x"2a1b0f",x"2c1a0f",x"181009",x"341d0c",x"513f33",x"422613",x"301d10",x"422816",x"382112",x"3d2413",x"311d0e",x"876043",x"8c6448",x"9d7150",x"986e4e",x"9a6d4d",x"936749",x"986d4d",x"a37856",x"8b6345",x"976b4b",x"835c41",x"996e4f",x"996e4f",x"a07352",x"996e4d",x"a07453",x"8c6144",x"896144",x"936b4b",x"9a6f4e",x"9c7252",x"9f7352",x"936748",x"9e7252",x"906747",x"7b553c",x"865e41",x"926647",x"8b6041",x"946847",x"8b6043",x"976c4c",x"895e41",x"885f42",x"93694b",x"94694b",x"8e6647",x"92694a",x"8b6244",x"79563b",x"704f35",x"5b3f2c",x"4d3626",x"4d3626",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a210f",x"3a210f",x"150e07",x"150e07",x"150e07",x"383129",x"383129",x"2f241b",x"4d2d17",x"4d2d17",x"251509",x"150e07",x"150e07",x"150e07",x"482813",x"412611",x"422612",x"391f0d",x"402511",x"3b200e",x"3c220f",x"432612",x"452712",x"3e220f",x"30190a",x"190f07",x"74523a",x"8b6345",x"8f6545",x"906747",x"896142",x"825b40",x"825b40",x"78533a",x"8f6345",x"875f41",x"956a4b",x"91684a",x"91684a",x"875e42",x"996f4f",x"946a4b",x"986f4f",x"966c4f",x"886043",x"8b6345",x"896144",x"936a4b",x"95694a",x"9a6f50",x"875e41",x"8c6245",x"956b4b",x"8c6246",x"966c4d",x"865d40",x"8d674a",x"8f6649",x"8b6245",x"8e6649",x"825b40",x"75533a",x"6c4b32",x"442f1f",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472814",x"472814",x"442611",x"39200e",x"3f2310",x"3e220f",x"3b210e",x"361d0c",x"331c0c",x"3c220f",x"3a200e",x"3b200e",x"3c200d",x"311b0b",x"2a180b",x"2a180b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2a180b",x"2a180b",x"150e07",x"221409",x"291609",x"150e07",x"51311c",x"2f2017",x"52473d",x"150e07",x"150e07",x"150e07",x"150e07",x"211308",x"150e07",x"150e07",x"150e07",x"150e07",x"312319",x"302117",x"352a22",x"352a22",x"000000",x"554032",x"554032",x"301a0b",x"231409",x"1e1208",x"241509",x"251509",x"26160a",x"150e07",x"2d1a0c",x"2d1a0c",x"27170b",x"2e1b0c",x"2b190c",x"27170b",x"2a190b",x"28180b",x"24150a",x"28170b",x"2f1c0d",x"27170b",x"27170b",x"24160a",x"221409",x"2a190b",x"201309",x"26160a",x"27170a",x"241509",x"231509",x"241509",x"211309",x"24150a",x"26160a",x"211409",x"221409",x"1a1008",x"211309",x"231409",x"1d1108",x"1d1108",x"1c1108",x"1b1008",x"1a1008",x"211308",x"1c1108",x"201208",x"191008",x"150e07",x"191008",x"211309",x"25160a",x"180f08",x"1b1008",x"1c1108",x"150e07",x"201309",x"351d0d",x"150e07",x"825e3f",x"805d3e",x"7d5b3d",x"7f5b3d",x"805d3e",x"836041",x"836041",x"876343",x"876343",x"825e3f",x"7f5b3c",x"825d3f",x"7f5b3d",x"805c3e",x"7d5a3b",x"866243",x"856243",x"866343",x"7e5c3d",x"77573a",x"836040",x"825f41",x"886444",x"8b6746",x"8a6442",x"886443",x"845f3f",x"825f3f",x"8b6645",x"8b6645",x"7a5839",x"7c593b",x"815d3e",x"805d3e",x"7b593c",x"7b583b",x"7f5c3d",x"836042",x"836041",x"846042",x"7f5c3f",x"815c3e",x"7f5b3d",x"825f3f",x"725136",x"815d3e",x"7f5b3b",x"8a6545",x"8b6745",x"8f6a47",x"876243",x"835f41",x"876343",x"825f41",x"8b6846",x"45362a",x"45362a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"473427",x"473427",x"41230f",x"3c200e",x"3b200d",x"3c210e",x"3c210e",x"39200e",x"3f230f",x"351c0c",x"311a0b",x"331c0c",x"3b210f",x"402410",x"412511",x"422611",x"3a210f",x"412511",x"3e220f",x"381f0d",x"381f0d",x"371f0d",x"3b200e",x"361e0d",x"351d0d",x"311c0d",x"331e0d",x"331d0d",x"341d0d",x"371f0e",x"381f0e",x"221409",x"1d1208",x"150e07",x"2c190b",x"351e0e",x"1a1008",x"341e0d",x"351f0e",x"2e1b0d",x"1f1309",x"150e07",x"150e07",x"2b190c",x"37200f",x"311d0e",x"160e07",x"2a190b",x"1a1008",x"180f07",x"3c2310",x"2d1a0c",x"201409",x"191008",x"150e07",x"36200f",x"392210",x"361f0f",x"2d1a0c",x"311c0d",x"1f1309",x"150e07",x"27160a",x"341d0d",x"3a2210",x"39210f",x"351e0d",x"2d1a0b",x"2d190b",x"311b0c",x"331d0d",x"3b2210",x"412713",x"432713",x"432712",x"412612",x"452914",x"462a14",x"442913",x"472914",x"462913",x"4a2c15",x"422712",x"422712",x"472a14",x"432813",x"4e2e16",x"573319",x"371f0e",x"402511",x"402511",x"2e1b0c",x"2b190b",x"2f1b0c",x"150e07",x"321d0d",x"39200f",x"3b2210",x"402511",x"3e220f",x"381f0d",x"3b200e",x"3c210e",x"361e0d",x"3b200e",x"381e0d",x"3e220e",x"3f230f",x"3a200d",x"412410",x"3b210e",x"3b200e",x"341b0b",x"361d0c",x"3e220f",x"3f2410",x"412511",x"432711",x"442712",x"432611",x"402410",x"3e230f",x"3c210e",x"3a200e",x"3c210f",x"3b210e",x"3e220f",x"371f0d",x"412611",x"3f2410",x"3f230f",x"412410",x"412411",x"432611",x"402410",x"412511",x"442712",x"412411",x"422511",x"3d2310",x"3d2310",x"432713",x"462913",x"472a14",x"3f2512",x"482a15",x"452914",x"482b15",x"472a14",x"3b2210",x"402612",x"442713",x"321d0d",x"301c0d",x"3a2210",x"150e07",x"311d0e",x"1b1108",x"1b1108",x"000000",x"000000",x"311f13",x"311f13",x"322013",x"362113",x"372112",x"341f11",x"2e1c10",x"23160d",x"18100a",x"311b0b",x"514034",x"452813",x"392111",x"3f2614",x"3f2614",x"3d2312",x"26160b",x"886145",x"78553d",x"9c7252",x"9b6f50",x"976b4b",x"9a6d4d",x"9d7251",x"805b41",x"9b7150",x"906647",x"875f43",x"8a6144",x"9c7152",x"9d7152",x"966b4a",x"976d4e",x"966a4b",x"6d4a35",x"896246",x"966c4b",x"9b7050",x"9b6f4f",x"8f6445",x"956a4a",x"906547",x"8e6346",x"8e6343",x"8b6040",x"895e40",x"956949",x"8c6142",x"95694a",x"8a6043",x"8a6143",x"8e6446",x"936a4b",x"906548",x"936b4b",x"8a6144",x"815a3f",x"745138",x"5d422d",x"4a3524",x"4a3524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412511",x"412511",x"150e07",x"150e07",x"150e07",x"29221b",x"29221b",x"291e15",x"4a2914",x"4a2914",x"271509",x"150e07",x"150e07",x"150e07",x"452612",x"402511",x"432612",x"391f0d",x"442712",x"402410",x"3a200e",x"432611",x"442712",x"412510",x"361d0c",x"1d1108",x"78543a",x"886043",x"906445",x"835d42",x"8a6144",x"8a6246",x"8a6043",x"76523a",x"8b6043",x"8a5f42",x"886145",x"8a6144",x"9a7051",x"8f6347",x"91674a",x"956b4d",x"9b7152",x"91684a",x"835b3f",x"8c6446",x"805a3f",x"936b4c",x"916748",x"966d4d",x"885e40",x"956a4c",x"986d4d",x"8d6244",x"986e4d",x"885e40",x"926a4d",x"956b4c",x"7a553b",x"8c6447",x"7f5a3f",x"684732",x"6c4b32",x"422d1c",x"412c1c",x"412c1c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492a15",x"492a15",x"452712",x"371e0d",x"381f0d",x"371e0d",x"3c210f",x"331c0b",x"341c0c",x"3c210f",x"341c0b",x"3c200e",x"41240f",x"2a170a",x"2f1a0b",x"2f1a0b",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29170a",x"29170a",x"150e07",x"1f1309",x"2c180a",x"150e07",x"52331e",x"2f2015",x"554c41",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1108",x"150e07",x"150e07",x"150e07",x"170f07",x"362418",x"312216",x"2b2119",x"2b2119",x"000000",x"594131",x"594131",x"2e190a",x"241509",x"221409",x"201309",x"221409",x"1f1209",x"150e07",x"211409",x"2c1a0c",x"24160a",x"29180b",x"2c1a0c",x"2d1b0d",x"2c1a0c",x"29190b",x"26170b",x"2c1a0c",x"2a190c",x"2e1b0c",x"221409",x"1e1209",x"23150a",x"29180b",x"211409",x"1b1108",x"26160a",x"27170a",x"231509",x"24150a",x"211409",x"231509",x"261609",x"211409",x"221409",x"1f1208",x"251509",x"201208",x"201208",x"251509",x"1c1108",x"1f1208",x"1d1108",x"1e1208",x"1d1108",x"1d1108",x"1e1208",x"211409",x"221409",x"150e07",x"1d1208",x"201309",x"1a1008",x"1a1008",x"1c1108",x"1c1108",x"3b210f",x"150e07",x"825f40",x"7f5d3f",x"846142",x"856343",x"825f40",x"825f3f",x"896546",x"886243",x"8b6646",x"856141",x"845f3f",x"846040",x"825f3f",x"815c3e",x"7a573a",x"765437",x"725035",x"785438",x"7d593d",x"7d5a3d",x"7f5c3d",x"7d5a3c",x"825e40",x"856142",x"805c3e",x"805d3e",x"815e3e",x"7d5a3b",x"7f5b3c",x"815d3f",x"805c3f",x"7c593d",x"825f40",x"7c5b3d",x"836041",x"846242",x"825f41",x"825e3f",x"846244",x"846041",x"856243",x"876243",x"7e5c3c",x"835f3f",x"856140",x"866041",x"7a583a",x"7b5739",x"7a5639",x"7b5639",x"825f40",x"835f40",x"846040",x"805c3e",x"825f3f",x"4a3628",x"4a3628",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"382f27",x"382f27",x"381e0c",x"371d0c",x"391e0d",x"3a200d",x"3f220f",x"3b200e",x"3a200e",x"3d220f",x"3c210f",x"391f0e",x"361e0d",x"3c210f",x"3f230f",x"3f2410",x"381f0d",x"3c210f",x"3b210f",x"3b220f",x"412611",x"412411",x"38200e",x"3a210f",x"1d1209",x"2d1a0c",x"150e07",x"180f08",x"2d190b",x"311c0d",x"331d0e",x"3b2210",x"402511",x"351f0e",x"201309",x"3a2110",x"38200f",x"150e07",x"3d2310",x"3d2411",x"150e07",x"150e07",x"150e07",x"38200f",x"2a190c",x"412712",x"3a2210",x"402612",x"39220f",x"3f2612",x"432813",x"150e07",x"150e07",x"150e07",x"39210f",x"150e07",x"150e07",x"38200f",x"150e07",x"3b2310",x"150e07",x"150e07",x"462914",x"150e07",x"26160a",x"462a14",x"412612",x"412612",x"3f2511",x"3e2411",x"150e07",x"2f1c0d",x"442813",x"462a14",x"462a14",x"492b15",x"452913",x"412612",x"402511",x"452813",x"432713",x"412511",x"3f2511",x"412512",x"3d2310",x"442712",x"4a2b14",x"573319",x"39210f",x"442712",x"3e2310",x"361f0d",x"391f0e",x"2e1a0c",x"150e07",x"2d190b",x"3e2410",x"381f0d",x"39200e",x"3b200e",x"381f0d",x"3b200d",x"381f0d",x"3a1f0d",x"391e0d",x"361d0c",x"351d0c",x"381f0d",x"3e220e",x"3f230f",x"3b200e",x"3e230f",x"3f230f",x"3d220f",x"3b200e",x"3d210f",x"3d220f",x"412410",x"422510",x"3b200e",x"412410",x"412511",x"452812",x"432611",x"412410",x"432611",x"452813",x"422712",x"402511",x"442713",x"422611",x"3f230f",x"432712",x"472914",x"462914",x"452813",x"492a13",x"482a14",x"472914",x"452914",x"402511",x"452813",x"462914",x"442813",x"422712",x"432712",x"432813",x"472a14",x"432813",x"422713",x"452913",x"452913",x"402612",x"462a15",x"402713",x"150e07",x"351f0e",x"191008",x"191008",x"000000",x"000000",x"301f12",x"301f12",x"352013",x"382214",x"321e11",x"341f11",x"2e1a0d",x"2b1a0e",x"181009",x"2f1a0b",x"534033",x"3c2311",x"422614",x"412715",x"3c2313",x"3e2412",x"27170b",x"805a3f",x"94694b",x"9d7453",x"956a4b",x"9b6e4d",x"9d7151",x"9f7352",x"966a4c",x"9a6f50",x"956b4b",x"92684a",x"8d6344",x"956c4e",x"8e6648",x"8e6546",x"996c4c",x"986c4c",x"865e42",x"a47856",x"946848",x"9c7453",x"93694a",x"966a4b",x"9b7151",x"93684a",x"9a6d4d",x"976b4b",x"8d6143",x"895f41",x"7d563b",x"976b4b",x"936749",x"896042",x"875f41",x"875f41",x"865f42",x"855e42",x"8d6445",x"8b6345",x"805b40",x"75533b",x"5e422e",x"493323",x"493323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b210e",x"3b210e",x"150e07",x"150e07",x"150e07",x"28221b",x"28221b",x"2b1f17",x"492a14",x"492a14",x"29160a",x"150e07",x"150e07",x"150e07",x"432511",x"3f2411",x"412511",x"3b200e",x"452812",x"3c210f",x"371e0d",x"442712",x"422611",x"412510",x"331a0b",x"190f07",x"926a4c",x"8d6446",x"855c41",x"8e6546",x"845c40",x"75523a",x"835c3f",x"916748",x"916646",x"94694a",x"8b6447",x"966d4d",x"926a4b",x"8e6748",x"956a4c",x"976b4c",x"8d664a",x"8e6649",x"664530",x"986d4d",x"835b40",x"956b4b",x"986e4f",x"956a4c",x"8a6143",x"8d6546",x"8e6546",x"865d40",x"9a714f",x"906747",x"8c664a",x"90674a",x"7e593d",x"8b6548",x"7d583c",x"755138",x"65462f",x"422d1d",x"452f1e",x"452f1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482a15",x"482a15",x"432611",x"361e0d",x"3a200e",x"3a200e",x"3c210f",x"3a1f0d",x"371e0d",x"361e0d",x"341c0b",x"3b200e",x"3f230f",x"2b180a",x"2a170a",x"2a170a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"261609",x"261609",x"150e07",x"1c1109",x"2a180b",x"150e07",x"4f3019",x"312015",x"5a4f45",x"150e07",x"150e07",x"150e07",x"150e07",x"241409",x"150e07",x"150e07",x"150e07",x"1a1008",x"2d2017",x"291c12",x"261c13",x"261c13",x"000000",x"523d2f",x"523d2f",x"361e0d",x"201208",x"241509",x"26160a",x"231509",x"26160a",x"150e07",x"29180b",x"221409",x"2c1a0c",x"29180b",x"29180b",x"2a190b",x"2d1b0c",x"2a180b",x"27170a",x"2a190b",x"2c1a0c",x"29180b",x"25160a",x"23150a",x"241509",x"241509",x"231409",x"1d1208",x"231409",x"201309",x"24150a",x"211409",x"231409",x"201309",x"211309",x"1e1208",x"211309",x"221309",x"211308",x"211308",x"201208",x"1f1208",x"241509",x"221409",x"211309",x"170f07",x"1f1208",x"1c1108",x"1f1208",x"1f1208",x"1f1309",x"1f1209",x"1c1108",x"180f07",x"191008",x"191008",x"211409",x"201309",x"39200e",x"150e07",x"7f5c3d",x"7a583c",x"815e41",x"846042",x"846042",x"856141",x"835f41",x"845f41",x"896444",x"7f5c3e",x"7f5c3d",x"825e3f",x"7e5c3d",x"855f40",x"7a583a",x"805c3d",x"7f5b3b",x"785637",x"815e3f",x"7f5c3e",x"835f40",x"83603f",x"856243",x"825f3f",x"815f40",x"876343",x"896545",x"8e6949",x"8d6949",x"866242",x"805e3f",x"836041",x"7f5b3e",x"745439",x"7c5b3e",x"7d5b3e",x"825f41",x"7b5a3d",x"805d3f",x"815d3f",x"866243",x"7b593c",x"7c5a3b",x"846140",x"876241",x"856040",x"7c593b",x"856040",x"825d3d",x"745335",x"896443",x"7f5b3d",x"876343",x"866241",x"8c6746",x"413328",x"413328",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"413429",x"413429",x"41230f",x"3e220f",x"3d210e",x"412410",x"422611",x"412511",x"3d230f",x"3b210f",x"412410",x"3c210f",x"3c210f",x"3d220f",x"3a200e",x"3c210f",x"371f0e",x"3e220f",x"391f0e",x"321c0c",x"3f2511",x"402411",x"3d2310",x"351d0d",x"3f2410",x"3b210f",x"371f0d",x"3a200e",x"3c210f",x"150e07",x"3a200e",x"150e07",x"361f0e",x"150e07",x"28170b",x"221409",x"341c0c",x"402310",x"422612",x"321d0d",x"2f1b0c",x"38200e",x"150e07",x"321c0d",x"180f08",x"2f1d0a",x"2b1b09",x"311f0a",x"311f0a",x"584b3e",x"361f0e",x"170f07",x"150e07",x"201309",x"2d1a0c",x"201309",x"3d2410",x"3d220f",x"371e0d",x"150e07",x"1c1108",x"251509",x"150e07",x"331b0b",x"361d0c",x"150e07",x"150e07",x"402410",x"3e2310",x"3f2410",x"3f2310",x"150e07",x"3d2310",x"3b200e",x"3e220f",x"412411",x"402511",x"422612",x"3f2411",x"3f2410",x"3c210f",x"3a200e",x"39200e",x"39200e",x"3a210f",x"402511",x"4b2c15",x"563318",x"482811",x"4c2a13",x"4a2b14",x"512e16",x"472811",x"4c2a13",x"502e15",x"4e2c14",x"4c2a13",x"4c2a13",x"4a2912",x"4f2d15",x"482d16",x"4f2e15",x"4e2e15",x"4c2b14",x"4f2e16",x"513017",x"54331a",x"4e2e16",x"533319",x"58361b",x"5a361b",x"563319",x"5b361b",x"58351b",x"523118",x"57331a",x"57361b",x"5b361c",x"522f17",x"4f2e16",x"482812",x"4b2a12",x"4d2c14",x"512f16",x"563218",x"4b2b14",x"4c2a13",x"442611",x"4a2913",x"4e2d15",x"563218",x"512f16",x"512e16",x"512e15",x"4e2b14",x"4e2c14",x"4f2d15",x"4d2b13",x"4d2b14",x"502c14",x"4d2c14",x"482711",x"442510",x"492912",x"4e2c15",x"43240f",x"3e210d",x"482810",x"40230d",x"4c2911",x"40230e",x"4d2c14",x"4e2d15",x"4a2913",x"4b2a13",x"4c2b14",x"492812",x"3d200e",x"3d200e",x"150e07",x"000000",x"301f12",x"301f12",x"362213",x"351f11",x"382112",x"321f10",x"2f1c0f",x"25180d",x"181009",x"2f1a0b",x"4e3e32",x"432614",x"412815",x"402614",x"432815",x"412713",x"341f0f",x"8b6549",x"956b4c",x"926a4d",x"946949",x"9f7252",x"a07454",x"9d7151",x"9d7050",x"9d7050",x"966c4c",x"8c6345",x"885e41",x"a37756",x"966a4a",x"8e6345",x"8a6043",x"8c6447",x"9a6f4f",x"a27553",x"a27554",x"936d4e",x"996e4d",x"926749",x"886043",x"966a49",x"8e6344",x"956847",x"95694a",x"885f42",x"886044",x"916648",x"94694b",x"8b6345",x"744f36",x"755138",x"8a6145",x"835c40",x"946a4b",x"8b6346",x"7c573d",x"7c5b41",x"634531",x"473121",x"473121",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311b0d",x"311b0d",x"150e07",x"150e07",x"150e07",x"28221a",x"28221a",x"2b1f16",x"492d1b",x"492d1b",x"371e0d",x"150e07",x"150e07",x"150e07",x"4e2c15",x"402511",x"3e2310",x"3b200e",x"432712",x"3c210e",x"381f0d",x"412511",x"442712",x"40230f",x"261106",x"1b1008",x"8d664a",x"8d6447",x"896043",x"936b4d",x"926648",x"7d593f",x"845c40",x"916848",x"8f6547",x"916648",x"815a3f",x"996f4e",x"986e4f",x"866042",x"91674a",x"966c4d",x"896144",x"825b3f",x"8c6243",x"90674a",x"875f42",x"7e573e",x"976d4d",x"956b4d",x"916748",x"93694a",x"8a6143",x"906647",x"92694b",x"8d6448",x"976e4f",x"986d4d",x"855d42",x"876043",x"724e36",x"7e593c",x"714f36",x"442e1e",x"452f1f",x"452f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462815",x"462815",x"452611",x"3c210f",x"3c210f",x"39200e",x"3a200e",x"3f230f",x"381f0d",x"39200e",x"341c0c",x"3c220f",x"41230f",x"301b0b",x"2b190b",x"2b190b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"29170a",x"29170a",x"150e07",x"1a1008",x"331c0d",x"150e07",x"502f18",x"2f2015",x"52493f",x"150e07",x"150e07",x"150e07",x"150e07",x"241409",x"150e07",x"150e07",x"150e07",x"170f07",x"322116",x"2b1b10",x"261b12",x"261b12",x"000000",x"553f31",x"553f31",x"2a1709",x"241509",x"221409",x"231409",x"211309",x"24150a",x"150e07",x"26160a",x"25160a",x"2a180b",x"26160a",x"28170a",x"241509",x"231409",x"211309",x"231409",x"29180b",x"2d1a0c",x"2b190b",x"231409",x"1e1208",x"25160a",x"29180b",x"241509",x"26160a",x"26160a",x"27170b",x"23150a",x"27170b",x"23150a",x"1c1108",x"1f1208",x"221409",x"1f1208",x"221409",x"221409",x"231409",x"1e1208",x"241509",x"241509",x"25150a",x"211309",x"221409",x"1f1209",x"201309",x"231409",x"1f1308",x"1a1008",x"201309",x"27160a",x"1d1108",x"170f07",x"1a1008",x"1b1108",x"1a1008",x"3d210f",x"150e07",x"876242",x"7c593c",x"825f40",x"825f41",x"7d5b3d",x"7a593a",x"805d3f",x"805e40",x"866243",x"825e40",x"876344",x"805d40",x"805d3e",x"7b593c",x"7c593c",x"7a593b",x"846040",x"7d5a3d",x"765637",x"785738",x"815e3f",x"7b593c",x"7a583b",x"755438",x"755236",x"7c593c",x"7a593c",x"886445",x"856143",x"79583a",x"7f5b3d",x"755438",x"7d5c3d",x"7a583b",x"7b5a3d",x"805e40",x"79573a",x"795839",x"825e40",x"815f41",x"7e5c3e",x"7d5b3d",x"8e6848",x"876344",x"805d3e",x"845f3f",x"815d3f",x"7c5a3c",x"846041",x"815e3f",x"7b573a",x"7b593a",x"815d3f",x"815d3f",x"7c5a3c",x"382c23",x"382c23",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"493a30",x"493a30",x"3f230f",x"3c200e",x"3b200d",x"3a200d",x"3d210e",x"3b220f",x"391f0d",x"371e0d",x"381f0d",x"3a200e",x"3c220f",x"3c210f",x"3e220f",x"3f2310",x"3c210f",x"381f0e",x"3f2511",x"3b210f",x"3b200e",x"3c210e",x"3f2410",x"39200e",x"301b0c",x"1c1108",x"150e07",x"39200e",x"2c1a0b",x"150e07",x"24150a",x"321d0d",x"311c0d",x"24150a",x"150e07",x"38200e",x"150e07",x"331d0d",x"170f07",x"231409",x"1a1008",x"381f0e",x"150e07",x"150e07",x"29180b",x"412511",x"371f0e",x"3b2310",x"412611",x"3d2411",x"3f2411",x"211409",x"38200f",x"150e07",x"150e07",x"39200f",x"3c230f",x"1e1208",x"2f1b0c",x"341c0c",x"201309",x"361e0e",x"391f0e",x"3b210f",x"432712",x"2b190b",x"3a220f",x"39200f",x"301b0c",x"251509",x"211309",x"321b0b",x"371f0d",x"3d220f",x"3f2310",x"3d220f",x"3d2310",x"3e2410",x"3f2411",x"432713",x"412611",x"432612",x"432712",x"3d2310",x"412611",x"432712",x"452812",x"201508",x"3a1f0c",x"472610",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1408",x"1d1208",x"1d1208",x"1f1408",x"1f1408",x"1c1208",x"221508",x"211508",x"211508",x"221608",x"201508",x"1b1108",x"1e1408",x"201408",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"301f13",x"301f13",x"362215",x"372113",x"362012",x"331f11",x"2f1d10",x"28190e",x"181009",x"321c0b",x"4e3e32",x"452916",x"3d2413",x"3c2414",x"422714",x"3f2412",x"2c1a0c",x"8a6245",x"9b7150",x"976c4d",x"976d4d",x"996f51",x"a67a58",x"9d7253",x"5d3e2c",x"8b6144",x"9c7050",x"94694a",x"865e41",x"9e7554",x"996c4c",x"845c40",x"94694b",x"8f6547",x"956a4a",x"a07957",x"a27656",x"a27756",x"8f6442",x"8e6341",x"906445",x"9b6f50",x"8a5f42",x"966a4a",x"8b6142",x"936949",x"896042",x"936848",x"966b4c",x"875e41",x"865d40",x"7f593d",x"865f42",x"855e40",x"865d41",x"8f6748",x"876245",x"78563d",x"5f422f",x"422b1d",x"422b1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3a200f",x"3a200f",x"150e07",x"150e07",x"150e07",x"322a23",x"322a23",x"2d231b",x"4a2c19",x"4a2c19",x"2c180b",x"150e07",x"150e07",x"150e07",x"4b2b14",x"432612",x"442713",x"3a200e",x"412511",x"3c210e",x"361d0c",x"3e220f",x"432711",x"3b210e",x"301809",x"1b1007",x"92694b",x"8a6346",x"90674a",x"8b6447",x"855c41",x"916b4c",x"865d40",x"956b4c",x"956a4b",x"936a4b",x"895f42",x"8d6447",x"8b6447",x"825d42",x"946c4c",x"91684a",x"8d6346",x"936c4c",x"896345",x"8f6547",x"8d6648",x"8c6445",x"7b573f",x"9b7051",x"966a4a",x"7f583e",x"8a6143",x"966d4d",x"967251",x"80583c",x"876043",x"8b6041",x"80593b",x"7e573d",x"75513a",x"745036",x"6f4e35",x"483221",x"473120",x"473120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472915",x"472915",x"3f2310",x"3a200e",x"3b210e",x"3a200e",x"3c210f",x"3d220f",x"341d0c",x"381f0e",x"361e0d",x"3b210e",x"3f230f",x"271609",x"2e190a",x"2e190a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1b0c",x"2f1b0c",x"231509",x"150e07",x"331d0c",x"191008",x"523119",x"302015",x"413830",x"150e07",x"150e07",x"150e07",x"150e07",x"221309",x"150e07",x"150e07",x"150e07",x"150e07",x"322217",x"27190f",x"231910",x"231910",x"000000",x"533d2f",x"533d2f",x"351e0d",x"241509",x"28170a",x"211409",x"1d1108",x"231409",x"150e07",x"2d1a0b",x"2a180b",x"26170a",x"2d1a0c",x"2b190c",x"211409",x"231509",x"25160a",x"27170a",x"2b190c",x"27170a",x"241509",x"221409",x"211309",x"221409",x"28170a",x"28170a",x"221409",x"221409",x"251509",x"251509",x"1f1208",x"211309",x"1f1208",x"1e1208",x"1d1108",x"201309",x"1e1208",x"251609",x"1f1208",x"221409",x"1d1108",x"1c1108",x"201208",x"201309",x"1a1008",x"1d1108",x"150e07",x"28170a",x"231409",x"1d1108",x"201309",x"201309",x"180f07",x"1a1008",x"170f07",x"1b1108",x"1b1108",x"3b210e",x"150e07",x"815f41",x"7f5d3f",x"7e5b3e",x"825f41",x"815e40",x"805e40",x"866343",x"7e5c3e",x"815d3f",x"896645",x"866243",x"835f41",x"7e5c3f",x"815e3f",x"866241",x"8b6646",x"846142",x"846041",x"856143",x"846143",x"765436",x"846142",x"7c5a3d",x"785739",x"765337",x"765438",x"715036",x"78583a",x"7c5a3d",x"7d5a3e",x"7d5b3d",x"7e5c3e",x"805e40",x"7b5a3d",x"77563a",x"76563a",x"7a593c",x"805e3f",x"805d3f",x"815e3f",x"7d5b3d",x"846343",x"876344",x"836041",x"886445",x"876242",x"886344",x"8a6545",x"886445",x"866242",x"8a6545",x"886545",x"7b5838",x"866243",x"7e5b3e",x"302921",x"302921",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a3e34",x"4a3e34",x"381e0d",x"3a200d",x"381e0d",x"361c0c",x"351c0b",x"371d0c",x"351d0d",x"39200e",x"2e180a",x"371e0d",x"381f0e",x"381f0e",x"3a200e",x"3e230f",x"3c210f",x"38200e",x"38200e",x"3d230f",x"412410",x"3c210e",x"361e0d",x"3a210f",x"38200e",x"301a0b",x"351f0e",x"311b0c",x"341e0e",x"361f0e",x"371f0e",x"3b2210",x"3c2311",x"351f0f",x"29180b",x"311c0d",x"331d0d",x"3a2110",x"38200f",x"39210f",x"412612",x"2b190b",x"191008",x"311c0c",x"371f0e",x"2c180b",x"221409",x"2e1b0c",x"301c0d",x"25160a",x"341e0e",x"311b0c",x"301a0b",x"2d190b",x"2e1b0c",x"351f0e",x"392110",x"3b2210",x"412612",x"301c0d",x"39200f",x"39200e",x"29170b",x"37200f",x"3a2110",x"402612",x"412712",x"412612",x"3f2410",x"371f0e",x"361e0d",x"381f0d",x"351d0c",x"3d220f",x"422611",x"432711",x"402511",x"412611",x"3e2411",x"402511",x"402612",x"432712",x"412511",x"402410",x"3d220f",x"3f2310",x"422611",x"1b1108",x"56493e",x"4b2a12",x"3d210e",x"3b200e",x"3c200e",x"3a200d",x"351d0c",x"381f0d",x"3b200e",x"381f0d",x"351d0d",x"3a200e",x"371d0d",x"3b200e",x"3f230f",x"3c210e",x"3f220f",x"391f0d",x"391f0d",x"361d0c",x"361c0c",x"371d0c",x"3a200e",x"40230f",x"371d0c",x"3b210e",x"3e230f",x"391f0e",x"3a200e",x"3e220f",x"422510",x"412310",x"422611",x"462812",x"41250f",x"44260f",x"40240f",x"422711",x"442811",x"472911",x"482b13",x"40240f",x"4c2c15",x"492a12",x"4a2a13",x"472912",x"422611",x"472a14",x"452813",x"442712",x"422611",x"452813",x"452712",x"422611",x"472914",x"452813",x"462913",x"452712",x"422511",x"3b210f",x"432611",x"432712",x"452812",x"462813",x"432713",x"3b210e",x"39200e",x"3c210f",x"3e220f",x"432611",x"150e07",x"1a1008",x"1a1008",x"2f1e13",x"2f1e13",x"362214",x"372112",x"382112",x"372113",x"2d1b0e",x"2f1c0f",x"181009",x"38200f",x"4d3f35",x"472916",x"452a17",x"422716",x"3f2514",x"442814",x"311c0e",x"8b6447",x"92684b",x"986d4e",x"9a6f4f",x"a37857",x"a07352",x"986d4e",x"916748",x"976b4c",x"966b4c",x"9d7150",x"865e40",x"a27655",x"865d41",x"81593d",x"8f6749",x"6c4832",x"92694b",x"a47a58",x"986e4e",x"976c4e",x"986b48",x"906544",x"8a6040",x"9b6f4e",x"9c7050",x"986b4b",x"966a4a",x"956a4b",x"926647",x"926748",x"94694b",x"896141",x"825b3f",x"7b563a",x"896244",x"845d40",x"8b6346",x"896143",x"876247",x"7a573e",x"5e422e",x"483223",x"483223",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381f0e",x"381f0e",x"150e07",x"150e07",x"150e07",x"362f27",x"362f27",x"31261d",x"4a2a15",x"4a2a15",x"29170a",x"150e07",x"150e07",x"150e07",x"4d2d15",x"422612",x"442713",x"3c210f",x"422611",x"3b200e",x"3c210e",x"3f230f",x"3d220f",x"371d0c",x"361c0b",x"1a1008",x"845b3f",x"8d6445",x"90694b",x"946a4b",x"906748",x"8b6648",x"6f4b33",x"8b6243",x"936a4b",x"996f50",x"926849",x"90674a",x"8d6648",x"986f50",x"876047",x"976d4e",x"8b6447",x"8b674a",x"855d42",x"866143",x"875f43",x"896044",x"986e4e",x"8f6549",x"906748",x"946a4a",x"8d6344",x"966c4d",x"8d6c4d",x"936b4c",x"896144",x"855c3e",x"7d5739",x"7e573a",x"815b41",x"745138",x"6a4a32",x"432d1d",x"442e1d",x"442e1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2b15",x"4c2b15",x"422510",x"381f0d",x"39200e",x"3a200e",x"412511",x"3c210e",x"341c0c",x"39200e",x"341c0c",x"381f0d",x"3d220e",x"2d190b",x"301b0c",x"301b0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"432511",x"432511",x"1d1208",x"180f07",x"150e07",x"2d190b",x"150e07",x"160e07",x"3b210f",x"150e07",x"543119",x"312015",x"41372f",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"150e07",x"150e07",x"150e07",x"1a1008",x"352316",x"291a0f",x"22170f",x"22170f",x"000000",x"544135",x"544135",x"341d0d",x"221409",x"1d1108",x"25150a",x"211309",x"1a1008",x"150e07",x"2e1b0c",x"27170a",x"301c0d",x"2c1a0c",x"2a190b",x"2a190b",x"27170b",x"25160a",x"231409",x"27160a",x"29180a",x"26160a",x"231409",x"231409",x"1e1208",x"231409",x"1f1208",x"211309",x"231409",x"211309",x"1f1208",x"261609",x"221409",x"211309",x"201208",x"1d1108",x"1d1108",x"201309",x"1f1208",x"211309",x"1e1108",x"1e1208",x"1d1108",x"1c1108",x"1d1108",x"201308",x"150e07",x"1f1208",x"201308",x"211309",x"1e1208",x"251509",x"1e1208",x"1a1008",x"211409",x"1e1208",x"1e1208",x"201308",x"391f0d",x"150e07",x"8b6646",x"836144",x"856142",x"856243",x"7f5d3e",x"815e41",x"7a593a",x"805d3e",x"7d5b3d",x"815e3f",x"835f41",x"886444",x"825f41",x"856243",x"836142",x"825f40",x"7f5c3f",x"7e5d3f",x"78563a",x"825d3c",x"815d3e",x"815f41",x"7e5c3e",x"805d3f",x"826040",x"896545",x"886444",x"856143",x"826041",x"836042",x"846143",x"825e41",x"846042",x"805e42",x"7c5b3d",x"805e40",x"78573a",x"7b5a3e",x"735438",x"805c3e",x"835f41",x"815e3f",x"866343",x"886444",x"866243",x"866343",x"866344",x"846041",x"835f41",x"815e41",x"7b593c",x"835d3e",x"85603f",x"886445",x"835f40",x"3b2e24",x"3b2e24",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"54473c",x"54473c",x"381e0d",x"3a200d",x"391f0d",x"3b200e",x"3a200e",x"331c0c",x"3d210f",x"351d0c",x"361e0d",x"361e0d",x"3a200e",x"3c220f",x"3b220f",x"3e2310",x"3b210f",x"3a210f",x"3d2310",x"3b210f",x"39200f",x"371f0d",x"39200f",x"2f190a",x"412511",x"341d0d",x"341d0d",x"341d0d",x"3c2310",x"37200f",x"38200e",x"3d230f",x"3d2310",x"351f0e",x"3d2310",x"3f2411",x"38200f",x"3b220f",x"3e2411",x"3e2310",x"331c0c",x"371f0e",x"3a210f",x"351d0d",x"3b210f",x"3d220f",x"371f0e",x"3b210f",x"3b2210",x"3d2411",x"3b2311",x"3d2411",x"3a210f",x"3b220f",x"3b220f",x"3c220f",x"3f2310",x"3d2310",x"361f0e",x"3c210f",x"311c0c",x"311c0c",x"3d2310",x"3c220f",x"3e230f",x"3f2411",x"402512",x"402511",x"402511",x"3d2310",x"402511",x"3c220f",x"391f0e",x"3b210e",x"3d220f",x"3e2410",x"3f2310",x"412511",x"3c210f",x"3d220f",x"3f2411",x"3b2210",x"432712",x"402410",x"3d220f",x"3a220f",x"462813",x"231608",x"493b2f",x"593318",x"553118",x"4a2a13",x"4d2a13",x"472711",x"432410",x"422410",x"3f220e",x"452610",x"452611",x"422410",x"4a2a13",x"492a13",x"472812",x"452611",x"41230e",x"43240f",x"442510",x"442510",x"462711",x"472711",x"472711",x"4b2913",x"4b2912",x"4d2b14",x"4a2912",x"4a2913",x"4e2d15",x"4f2d15",x"4f2c15",x"4f2d15",x"512d15",x"502e15",x"4c2b13",x"432511",x"522f16",x"3c1f0d",x"512f15",x"4f2c13",x"502d14",x"532f15",x"513015",x"533016",x"512f16",x"4d2c14",x"4d2c15",x"4f2d15",x"4e2d15",x"533117",x"4b2a14",x"4d2c14",x"543117",x"502e16",x"4a2912",x"472711",x"533117",x"4e2c14",x"4d2a13",x"4c2b13",x"512f15",x"4f2d15",x"512e15",x"553118",x"573419",x"523017",x"4e2d16",x"4f2e15",x"512f16",x"4e2d15",x"4b2b14",x"150e07",x"150e07",x"321f13",x"321f13",x"362214",x"382212",x"372011",x"372112",x"2f1c0f",x"321e10",x"191109",x"412612",x"564336",x"452915",x"432715",x"382112",x"432715",x"452915",x"29180b",x"815a3f",x"936849",x"946949",x"986e4e",x"a47957",x"986b4c",x"9e7251",x"956a4b",x"966b4c",x"9a6d4d",x"986e4e",x"93694a",x"9d7251",x"9c704e",x"926647",x"90684a",x"885e43",x"91694c",x"9d7856",x"986d4e",x"9c7050",x"93684a",x"8f6443",x"906443",x"976a48",x"916647",x"996d4e",x"956b4a",x"936847",x"8a5f41",x"926748",x"8c6547",x"8c6243",x"936a4a",x"8b6243",x"78543a",x"8a6144",x"8c6546",x"916749",x"8a6448",x"7a583d",x"5d422e",x"473222",x"473222",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"301b0b",x"301b0b",x"150e07",x"150e07",x"150e07",x"3a332b",x"3a332b",x"2d231b",x"462915",x"462915",x"261509",x"150e07",x"150e07",x"150e07",x"4c2c15",x"452913",x"452712",x"3d220f",x"3f2410",x"3a200e",x"3d220f",x"3e230f",x"3c210f",x"381e0d",x"331a0b",x"1d1108",x"8c6244",x"825c40",x"966c4e",x"8f6647",x"886043",x"916c4e",x"845c41",x"896143",x"8b6244",x"906748",x"896044",x"956c4c",x"936a4b",x"986f50",x"966e4e",x"8c6548",x"866042",x"8b6347",x"8d6445",x"865f43",x"835d40",x"7b563c",x"966b4d",x"886043",x"8c6548",x"976c4e",x"8c6445",x"8d674a",x"8b6446",x"977151",x"8b6347",x"8f6749",x"8b6141",x"7a5438",x"755135",x"714f35",x"6f5037",x"46301f",x"432e1e",x"432e1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"502f18",x"502f18",x"412410",x"351d0c",x"371e0d",x"361d0c",x"3f2411",x"3a200e",x"351c0c",x"3a200d",x"351d0c",x"3b200e",x"3a1f0d",x"28160a",x"2b180a",x"2b180a",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"432511",x"432511",x"2a180b",x"180f07",x"150e07",x"25150a",x"201309",x"26160a",x"3a200e",x"150e07",x"4c2c17",x"2c2017",x"40382f",x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"150e07",x"150e07",x"150e07",x"211309",x"342216",x"29190f",x"1f160f",x"1f160f",x"000000",x"564134",x"564134",x"3d2411",x"26160a",x"201309",x"150e07",x"25160a",x"1d1208",x"150e07",x"29180b",x"2d1a0b",x"28170a",x"221409",x"2b190b",x"2c190c",x"29180b",x"221409",x"231409",x"27160a",x"2a190b",x"25160a",x"27160a",x"27170a",x"221409",x"25160a",x"251509",x"231409",x"251509",x"251509",x"221409",x"241509",x"211309",x"211309",x"26160a",x"27160a",x"221409",x"1e1208",x"1c1108",x"221409",x"201309",x"1e1208",x"1c1108",x"150e07",x"150e07",x"1c1108",x"1d1108",x"211409",x"201309",x"211409",x"24150a",x"26160a",x"221409",x"211409",x"1a1008",x"1c1108",x"1e1208",x"150e07",x"3b200e",x"150e07",x"8a6545",x"856243",x"7f5d3e",x"846142",x"825f40",x"835f40",x"856142",x"8a6747",x"825f40",x"805b3e",x"846041",x"815f41",x"846243",x"856243",x"8b6646",x"886344",x"836041",x"7d5b3d",x"866242",x"815c3d",x"7d5b3c",x"7f5b3e",x"7f5c3e",x"835f40",x"846041",x"815e3f",x"805c3e",x"7b593c",x"7f5c3d",x"765536",x"805d3d",x"755436",x"7c5a3e",x"805e40",x"7d5b3d",x"846142",x"78583b",x"7e5c3e",x"7f5d3f",x"896647",x"805e3f",x"805b3e",x"815e40",x"856143",x"876344",x"886444",x"876344",x"866143",x"846142",x"805d3e",x"856141",x"7f5b3c",x"7a593d",x"7b5a3c",x"815e3f",x"342c23",x"342c23",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"5e4f43",x"5e4f43",x"432611",x"432511",x"412511",x"422611",x"412511",x"412511",x"3e230f",x"3c220f",x"381f0e",x"3f2411",x"3a200e",x"331c0b",x"2f1a0a",x"331c0b",x"361d0c",x"3a200d",x"3a200e",x"3f2310",x"351e0e",x"3a210f",x"3c2310",x"38200e",x"371f0e",x"361e0e",x"381f0e",x"371f0e",x"361f0e",x"39200f",x"39200f",x"3c220f",x"3d2310",x"3f2410",x"3f2410",x"3f2410",x"3f2411",x"402511",x"3e2410",x"3b210f",x"351e0e",x"3e2410",x"3c220f",x"3b2210",x"3d2310",x"3e2310",x"3e2310",x"3e2411",x"3f2511",x"402612",x"432712",x"381f0d",x"371e0d",x"3c210f",x"3c210f",x"3b210f",x"3e220f",x"3f2410",x"412410",x"3c210f",x"39200f",x"3e2411",x"442713",x"432712",x"3e2310",x"402511",x"482b15",x"452913",x"492c15",x"452913",x"442813",x"432712",x"432712",x"462913",x"432712",x"472a14",x"452913",x"412511",x"452712",x"472914",x"402511",x"3f2410",x"3d2210",x"3c210f",x"3a200e",x"472914",x"462914",x"1c1208",x"4d3728",x"3e220f",x"29170a",x"241509",x"28160a",x"241509",x"1e1208",x"1c1108",x"201208",x"1e1208",x"1f1209",x"221409",x"1b1108",x"1e1209",x"211309",x"170f07",x"1d1208",x"1f1209",x"1e1208",x"201309",x"190f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"241708",x"281909",x"281909",x"261809",x"1c1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"150e07",x"150e07",x"150e07",x"170f07",x"170f07",x"180f07",x"180f07",x"191008",x"1d1208",x"190f08",x"1e1209",x"27170b",x"25160a",x"26160a",x"211409",x"221309",x"1f1209",x"1d1208",x"1f1208",x"231409",x"28170b",x"28170b",x"342114",x"342114",x"362113",x"352012",x"372111",x"2e1a0f",x"321d0f",x"2e1b0e",x"1a1109",x"3e2310",x"534133",x"452917",x"3f2615",x"3e2614",x"402715",x"442815",x"29180b",x"875e41",x"95694b",x"986d4d",x"9c7051",x"9e7554",x"a07453",x"9f7352",x"a07352",x"9e7251",x"9a6f4e",x"95694a",x"926748",x"a37756",x"9b7050",x"906648",x"8c6446",x"734e36",x"825d42",x"977051",x"9b7150",x"976b4b",x"956b4c",x"8f6649",x"765136",x"906543",x"906547",x"996d4d",x"94694a",x"8c6244",x"875d3f",x"906647",x"946a4a",x"8c6243",x"8c6446",x"7e583c",x"845d40",x"845c3f",x"906648",x"8d6548",x"866043",x"7d593e",x"5f432f",x"4f3826",x"4f3826",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200e",x"38200e",x"150e07",x"150e07",x"150e07",x"3b332b",x"3b332b",x"231c15",x"492a17",x"492a17",x"331c0c",x"150e07",x"150e07",x"150e07",x"462813",x"442813",x"432712",x"3f2411",x"3f2410",x"391f0d",x"3d210f",x"3c210e",x"3e220f",x"3e220e",x"361d0c",x"190f07",x"896043",x"8e6547",x"996f4f",x"93694b",x"8f6748",x"91694b",x"7d573b",x"7d573c",x"745036",x"8f6647",x"8b6245",x"91674a",x"906748",x"966b4c",x"8d674a",x"8e684a",x"936a4b",x"8e6547",x"875f43",x"805a3e",x"8b6245",x"876043",x"886144",x"845d41",x"8a6345",x"936a4b",x"8f6546",x"9a6f4f",x"8b6345",x"946d4e",x"90694a",x"875f42",x"8f6649",x"7e583b",x"735035",x"5f3e2b",x"694932",x"422e1e",x"432e1e",x"432e1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2c16",x"4a2c16",x"422511",x"361d0d",x"2f180a",x"361d0c",x"3d220f",x"391f0d",x"361d0c",x"381f0d",x"381f0d",x"412510",x"40230e",x"281609",x"301c0c",x"301c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"4e2c15",x"4e2c15",x"512e16",x"201309",x"150e07",x"150e07",x"27160a",x"231509",x"2c180a",x"3e2410",x"150e07",x"4c2c16",x"2f2017",x"40372e",x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"150e07",x"150e07",x"150e07",x"170f07",x"322116",x"2b1b10",x"21170f",x"21170f",x"000000",x"584334",x"584334",x"351e0e",x"27160a",x"27160a",x"221308",x"25160a",x"201309",x"150e07",x"2c1a0c",x"2d1a0c",x"2a190b",x"2b190c",x"2d1a0c",x"26160a",x"2b180b",x"26160a",x"1e1208",x"27170b",x"2d1a0c",x"2d1a0c",x"2a190b",x"29180b",x"25150a",x"241509",x"241509",x"251509",x"211309",x"231409",x"201208",x"1b1108",x"211409",x"27170a",x"26160a",x"25160a",x"24150a",x"29170b",x"211409",x"211409",x"241509",x"28170a",x"211409",x"24150a",x"241509",x"1f1208",x"221409",x"211409",x"221409",x"231409",x"221409",x"1e1208",x"221409",x"211309",x"201309",x"150e07",x"150e07",x"170f07",x"361d0c",x"150e07",x"8b6746",x"7e5b3d",x"7e5b3c",x"7e5b3d",x"7f5d3e",x"7d5b3d",x"8a6747",x"825f3f",x"896545",x"8a6645",x"825d3f",x"825e3f",x"896647",x"8d6a4a",x"8a6748",x"7b593c",x"725136",x"704f34",x"67482d",x"825f3f",x"805d40",x"846143",x"8d694a",x"896445",x"896443",x"846042",x"8f6b4b",x"886546",x"8a6647",x"805d3e",x"805c3b",x"7c593a",x"846142",x"7a583b",x"745336",x"725236",x"7b5a3c",x"7a583b",x"836244",x"7e5c3d",x"815f40",x"8b6545",x"835e40",x"815e3f",x"8b6849",x"8f6c4c",x"926d4c",x"7b593d",x"7b573a",x"735135",x"6f4c31",x"825e40",x"836042",x"8b6646",x"8b6748",x"3c2f26",x"3c2f26",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"522f16",x"522f16",x"4d2c14",x"4a2912",x"4b2b14",x"4c2b13",x"4f2d15",x"4e2d16",x"4b2a14",x"4a2912",x"482812",x"4a2913",x"492a13",x"4e2d15",x"4b2b13",x"472711",x"462611",x"482812",x"462711",x"523017",x"513018",x"57331a",x"533119",x"4b2a14",x"55341a",x"4d2d16",x"513017",x"4e2d15",x"533219",x"4b2b14",x"4a2a13",x"502d15",x"482913",x"4d2c14",x"3f220f",x"492812",x"4f2e16",x"4c2c15",x"472812",x"432611",x"402410",x"472812",x"41230f",x"41240f",x"412410",x"4c2c15",x"4b2c15",x"432611",x"4b2a14",x"4a2a14",x"482812",x"432510",x"482811",x"4a2b12",x"452711",x"3a1e0a",x"492a11",x"472811",x"472911",x"492a12",x"472811",x"442611",x"482912",x"442711",x"442710",x"42240f",x"422510",x"462711",x"4a2913",x"482913",x"4b2b14",x"4c2c15",x"4b2b15",x"4b2b15",x"4b2c15",x"4d2e16",x"502f16",x"4e2e15",x"4d2d14",x"4c2c13",x"4d2d14",x"4a2b12",x"512f15",x"513015",x"4a2c12",x"4d2c13",x"522f16",x"311c0d",x"3b3128",x"4c2c15",x"422612",x"3d2310",x"371f0e",x"39200e",x"381f0d",x"341c0c",x"311a0b",x"281509",x"2f190b",x"3e2411",x"351e0e",x"331c0c",x"39200e",x"351f0e",x"3d2310",x"3c2310",x"3b2210",x"3a2210",x"2f1b0c",x"150e07",x"150e07",x"150e07",x"150e07",x"211308",x"150e07",x"2e1a0b",x"301b0b",x"150e07",x"150e07",x"150e07",x"201308",x"2c180a",x"251509",x"150e07",x"28170a",x"37200f",x"3a220f",x"361f0d",x"38210d",x"281809",x"2b1a0a",x"331c0b",x"2d190b",x"311c0c",x"150e07",x"211409",x"351f0f",x"150e07",x"37210f",x"301b0c",x"201309",x"150e07",x"2f1b0d",x"38210f",x"28180b",x"1f1209",x"2e1a0c",x"38200f",x"3a2210",x"442914",x"422813",x"422712",x"3e2411",x"3e2310",x"3b220f",x"39200e",x"3b210f",x"3b2210",x"3c2310",x"231409",x"231409",x"322013",x"322013",x"311e12",x"362011",x"3a2212",x"2e1b0f",x"311d0f",x"2e1c0f",x"1a110a",x"3b210f",x"503d32",x"432815",x"402715",x"3e2615",x"412615",x"3e2412",x"331e0e",x"7e583d",x"94694b",x"976c4d",x"9b7150",x"9a7051",x"996f4f",x"9d7353",x"a07453",x"996e4d",x"977050",x"9a6e4d",x"95694a",x"a47857",x"9b7151",x"94694a",x"906648",x"8b6244",x"8b6549",x"8b6647",x"876044",x"8c6344",x"906646",x"8f6546",x"765139",x"734f38",x"7a5339",x"9d7150",x"936747",x"855e40",x"8d6243",x"8c6244",x"885f41",x"8d6546",x"876144",x"805a3f",x"855e41",x"79553b",x"8d6445",x"8b6447",x"845d42",x"745338",x"614530",x"4b3625",x"4b3625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d2310",x"3d2310",x"150e07",x"150e07",x"150e07",x"453d35",x"453d35",x"2c221a",x"4b2a16",x"4b2a16",x"2a180a",x"150e07",x"150e07",x"150e07",x"4c2b15",x"472a14",x"452813",x"402511",x"3c210f",x"3c210e",x"3e220f",x"3c220f",x"3b200e",x"3e220f",x"351c0c",x"1e1108",x"896042",x"8e6547",x"906748",x"815b3f",x"876043",x"876447",x"755138",x"7e583d",x"825b3f",x"906748",x"8a6245",x"9a7151",x"8c6447",x"926a4b",x"9e7553",x"9c7252",x"90694b",x"8c6447",x"886044",x"855d42",x"805a3e",x"865f42",x"8c6447",x"865e42",x"896245",x"8b6447",x"90674a",x"8e6649",x"8c6546",x"8b6547",x"825d41",x"7d583d",x"815b3f",x"6d4b34",x"755138",x"684630",x"674731",x"412d1d",x"432e1e",x"432e1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"52321c",x"52321c",x"442611",x"361d0c",x"361e0d",x"381e0d",x"3d220f",x"3d210e",x"3a1f0d",x"361d0c",x"331c0c",x"412410",x"432410",x"28160a",x"301c0c",x"301c0c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"4d2b14",x"482a13",x"492b14",x"150e07",x"321c0d",x"4a2a14",x"2a190b",x"301d0d",x"251509",x"3c2310",x"150e07",x"4c2d16",x"312217",x"473e36",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2015",x"281a0f",x"1e160f",x"1e160f",x"000000",x"524135",x"524135",x"38200f",x"29180b",x"211309",x"211409",x"241509",x"231509",x"150e07",x"2d1a0c",x"2a180b",x"2a190c",x"2a190b",x"2a190b",x"28180b",x"2b190c",x"2a190b",x"24160a",x"201309",x"1c1108",x"26160a",x"25150a",x"26160a",x"27170b",x"27170a",x"2b180b",x"251509",x"241509",x"221309",x"1f1208",x"1a1008",x"201208",x"27170b",x"24150a",x"211409",x"231509",x"25160a",x"201309",x"25160a",x"201309",x"231509",x"211409",x"221409",x"1d1108",x"221409",x"1c1108",x"1f1208",x"1d1108",x"231409",x"241509",x"1e1208",x"201309",x"1c1108",x"1b1008",x"150e07",x"170f07",x"190f07",x"371e0d",x"150e07",x"8c6848",x"866445",x"846142",x"846242",x"846042",x"805c3e",x"866242",x"825f41",x"815c3d",x"7d5a3d",x"866242",x"886444",x"856142",x"866243",x"886343",x"826040",x"8a6645",x"8d6848",x"846142",x"8d6b4a",x"896b4b",x"866445",x"8d6949",x"8b6848",x"8b6748",x"8d6949",x"8b6747",x"886545",x"886544",x"7a5a3c",x"876243",x"815e41",x"856344",x"826143",x"7b5a3d",x"79593c",x"7e5c3e",x"78563a",x"866242",x"805e40",x"7c593b",x"78573a",x"876343",x"876444",x"846041",x"886343",x"8b6645",x"846041",x"866443",x"8c6848",x"896544",x"8c6b4a",x"8d6d4c",x"906c4a",x"936d4c",x"5f4738",x"5f4738",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2a13",x"4a2a13",x"351d0d",x"3c210f",x"3d220f",x"3e2310",x"3b2310",x"3f2411",x"2b180a",x"2d190a",x"150e07",x"2c180a",x"2b180a",x"2d190a",x"341d0c",x"361e0c",x"301a0b",x"301a0a",x"381f0d",x"371e0c",x"3f220f",x"3d2310",x"351e0e",x"3b200f",x"3e2310",x"3c2210",x"3d2310",x"412511",x"3f2410",x"3b200e",x"381e0d",x"3b210e",x"3c210f",x"3c220f",x"361e0d",x"39200f",x"452914",x"452913",x"3e2511",x"3d2411",x"402512",x"412612",x"472914",x"452914",x"412411",x"3e220f",x"3b210f",x"432713",x"412511",x"402410",x"3c210f",x"3d220f",x"3e220f",x"3a200e",x"341d0c",x"371e0d",x"371e0d",x"381f0d",x"3e220f",x"402410",x"3f2410",x"3f230f",x"3c210f",x"40230f",x"3b200e",x"422611",x"432712",x"472a14",x"452712",x"3f220f",x"3d210f",x"3f230f",x"3f2410",x"472914",x"462914",x"452813",x"3e2411",x"3b220f",x"432712",x"452812",x"3f2410",x"321c0c",x"351d0d",x"321c0c",x"3c2310",x"150e07",x"422612",x"3b220f",x"3f3025",x"4a2a13",x"412511",x"3d230f",x"3c210f",x"3f230f",x"3c220f",x"422511",x"371f0d",x"331c0c",x"331c0c",x"3d2310",x"3c220f",x"3d230f",x"391f0e",x"3a200e",x"371e0d",x"381f0e",x"3b210f",x"341d0d",x"412611",x"462914",x"361e0d",x"2d190b",x"2e190a",x"150e07",x"2d190a",x"191007",x"2c180a",x"150e07",x"351d0c",x"2f1a0a",x"241509",x"301a0b",x"150e07",x"331e0e",x"231409",x"191007",x"26160a",x"38210e",x"5d5145",x"2f1b0c",x"331d0d",x"1a1007",x"311b0c",x"150e07",x"3b200e",x"3b200e",x"301b0c",x"150e07",x"24150a",x"191008",x"28180b",x"150e07",x"150e07",x"412612",x"402511",x"422612",x"402511",x"3a200e",x"3a200e",x"422612",x"3f2411",x"402410",x"3f230f",x"3a200e",x"3e220f",x"3a200e",x"39200e",x"341c0c",x"361e0d",x"2b180a",x"2b180a",x"311f13",x"311f13",x"392314",x"372111",x"3c2312",x"341e11",x"311c0f",x"301d0f",x"1a110a",x"3d230f",x"4f3f33",x"452915",x"432816",x"402615",x"472b17",x"3f2513",x"29180b",x"7f573c",x"956b4c",x"9d7351",x"9a7051",x"9b7252",x"986e50",x"976e4e",x"9e7454",x"956a4b",x"997150",x"8b6245",x"93694a",x"9d7353",x"9e7352",x"916748",x"986d4c",x"855d41",x"7a563c",x"8a6448",x"876145",x"8f6547",x"875d40",x"865d3f",x"926749",x"80573c",x"694631",x"896144",x"8a6144",x"8f6445",x"895f41",x"916747",x"8a6344",x"805a3e",x"865e41",x"896143",x"896244",x"765339",x"896043",x"8b6446",x"74523a",x"7b583e",x"5a3f2b",x"473121",x"473121",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2411",x"3f2411",x"150e07",x"150e07",x"150e07",x"423a31",x"423a31",x"31241a",x"492914",x"492914",x"281609",x"150e07",x"150e07",x"150e07",x"553016",x"402612",x"412612",x"422511",x"3c210f",x"3b200e",x"3b210e",x"3c220e",x"381f0d",x"3b200e",x"371d0c",x"1b1008",x"835a3f",x"8b6244",x"876044",x"7f5a3e",x"815c40",x"7a573c",x"714c34",x"775439",x"825c3f",x"845d41",x"785338",x"90694a",x"875f43",x"986f50",x"9f7654",x"8d6648",x"825e42",x"7e593e",x"8c6346",x"825d41",x"815b3e",x"926a4b",x"92694a",x"865e41",x"8b6145",x"8b6244",x"8b6447",x"966c4d",x"7e593f",x"7a583e",x"8f6749",x"7e583d",x"7a563b",x"6b4931",x"61402d",x"704d35",x"694a34",x"4c3524",x"4a3423",x"4a3423",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2f1b",x"4c2f1b",x"3e220f",x"3a200e",x"381f0d",x"341c0b",x"3d220f",x"3b210e",x"331c0c",x"321b0b",x"371e0d",x"3f230f",x"452611",x"271509",x"2a190b",x"2a190b",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"4c2b15",x"4c2b15",x"3c2311",x"150e07",x"311b0c",x"482914",x"2b180b",x"412510",x"2d190b",x"371e0d",x"191008",x"4e2d17",x"2f2015",x"433b32",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"150e07",x"150e07",x"150e07",x"150e07",x"2d2016",x"2a1a10",x"231811",x"231811",x"000000",x"513d2f",x"513d2f",x"341e0e",x"241509",x"231509",x"201308",x"23150a",x"211309",x"150e07",x"29180b",x"2b190b",x"27170a",x"29180b",x"27170a",x"2d1a0b",x"29170a",x"27160a",x"2b190b",x"27170b",x"1d1208",x"201309",x"231509",x"221409",x"1f1309",x"1c1108",x"26160a",x"251509",x"241509",x"26160a",x"241509",x"211309",x"211308",x"24150a",x"28170a",x"241509",x"221409",x"231409",x"251509",x"211409",x"221409",x"211409",x"1f1309",x"26170a",x"1d1108",x"1a1008",x"1d1108",x"251509",x"1f1208",x"1e1208",x"201308",x"221409",x"201309",x"1f1309",x"1d1208",x"1b1008",x"1f1208",x"170f07",x"351d0c",x"150e07",x"825e3f",x"79583a",x"7d5a3d",x"7a583a",x"765639",x"78563a",x"7c5a3c",x"805e3e",x"846041",x"7d5b3c",x"7f5c3e",x"805d3e",x"825f41",x"7e5c3e",x"835f40",x"805c3f",x"846041",x"815e40",x"846142",x"846042",x"825e40",x"866345",x"886446",x"825f41",x"8a6544",x"835f3f",x"7f5b3d",x"815e40",x"846143",x"7e5c3e",x"886443",x"836041",x"78573a",x"6e4f34",x"745338",x"745437",x"755438",x"79583a",x"805d3e",x"7f5d3e",x"7d5c3e",x"7d5b3c",x"77563a",x"7d5a3c",x"856243",x"7e5b3e",x"825e40",x"825e40",x"805d3f",x"7f5c3e",x"896544",x"8a6545",x"8b6545",x"8d694a",x"8f6a4a",x"5f4d40",x"5f4d40",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4f2e15",x"4f2e15",x"39210f",x"3e2411",x"3f2410",x"341d0d",x"2e1a0b",x"301a0b",x"311b0b",x"2f1a0b",x"150e07",x"2c180a",x"311b0b",x"351d0c",x"3a200d",x"3b200d",x"351d0c",x"371e0c",x"311b0b",x"3f230e",x"361d0c",x"3b220f",x"412612",x"3a210f",x"3e2310",x"432712",x"39200f",x"3c220f",x"3c220f",x"402410",x"452812",x"3e220f",x"3a1f0e",x"402511",x"422611",x"412511",x"432612",x"412512",x"3d2310",x"412612",x"432712",x"442813",x"422612",x"412511",x"412611",x"402411",x"412612",x"3f2410",x"371f0e",x"331c0c",x"321b0b",x"331b0c",x"321a0b",x"351b0b",x"2c1609",x"2e180a",x"2e180a",x"381f0d",x"3d220f",x"3c210f",x"391f0d",x"371e0d",x"361d0c",x"351d0c",x"321a0b",x"361d0c",x"3a200e",x"381f0d",x"391f0d",x"3a1f0d",x"3e230f",x"3b210f",x"3a210f",x"39200f",x"3f2310",x"3a200e",x"3a200e",x"3a200e",x"331c0d",x"3e220f",x"361d0c",x"28160a",x"2e1a0b",x"361e0d",x"371f0e",x"150e07",x"402410",x"371f0e",x"3d2f25",x"4b2a12",x"3e2310",x"3b210f",x"412511",x"412511",x"432611",x"422611",x"432612",x"3f2511",x"422611",x"3a200e",x"3c210e",x"3e220f",x"402410",x"3f2411",x"3e2411",x"422612",x"432712",x"422612",x"29180b",x"1d1108",x"2f1a0b",x"2d190a",x"301b0b",x"301a0b",x"341d0c",x"361e0d",x"2f1a0b",x"381f0d",x"1f1208",x"341c0c",x"2e190a",x"150e07",x"150e07",x"321c0b",x"34200e",x"432711",x"3f240f",x"3d2310",x"3e2310",x"301b0c",x"311c0d",x"150e07",x"3e2410",x"25150a",x"2c190b",x"3c220f",x"38200f",x"1b1108",x"150e07",x"3f2411",x"311d0d",x"1e1209",x"412612",x"412612",x"150e07",x"150e07",x"341e0e",x"3d2310",x"452712",x"402411",x"3e2310",x"381f0d",x"351d0c",x"361d0c",x"361c0c",x"361c0c",x"311a0a",x"2b1508",x"361c0c",x"29170a",x"29170a",x"331f12",x"331f12",x"392415",x"392212",x"3c2414",x"382112",x"341e0f",x"301c0d",x"1a110a",x"3a220f",x"4b3d32",x"4b2d18",x"402615",x"402615",x"432916",x"3b2312",x"352010",x"7f583c",x"946a4b",x"92694a",x"986d4c",x"9c7352",x"987050",x"946c4c",x"996f4f",x"92694b",x"986f4f",x"8f6647",x"815a40",x"a17654",x"90694a",x"946a4a",x"865e41",x"7a553b",x"866044",x"936a4b",x"936b4c",x"916647",x"886042",x"805a3e",x"835b3f",x"7a5338",x"7e593e",x"896043",x"8b6244",x"8f6649",x"7e573b",x"825c40",x"875f43",x"896043",x"896144",x"8b6244",x"835c3f",x"815a3e",x"896144",x"835d41",x"7b583e",x"755239",x"583e2a",x"4b3523",x"4b3523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"321c0d",x"321c0d",x"150e07",x"150e07",x"150e07",x"413830",x"413830",x"32271f",x"4a2b17",x"4a2b17",x"311a0b",x"150e07",x"150e07",x"150e07",x"552f16",x"39210f",x"3f2411",x"3d220f",x"391f0d",x"361e0d",x"3a200e",x"341c0c",x"361e0d",x"3a200e",x"351c0b",x"1c1108",x"845d40",x"815c40",x"90684a",x"7e583e",x"825d41",x"8f6749",x"765137",x"7c573c",x"8c6345",x"8e6647",x"755137",x"845c3f",x"835c41",x"966d4d",x"976f50",x"8a6447",x"8b6447",x"866044",x"815b3f",x"886345",x"785339",x"956e4e",x"835b3f",x"865e41",x"926848",x"91684a",x"79553a",x"936a4b",x"8b6143",x"7e593e",x"956b4c",x"7e583e",x"7e593f",x"815a3f",x"6c4830",x"78543a",x"64452e",x"453120",x"463120",x"463120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543520",x"543520",x"3d210e",x"321c0c",x"341c0c",x"321c0c",x"3a200e",x"341b0b",x"371e0d",x"351c0c",x"381f0d",x"412510",x"462711",x"2c190b",x"2c190c",x"2c190c",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"39200f",x"39200f",x"1b1108",x"150e07",x"150e07",x"27160a",x"2c180b",x"180f07",x"271609",x"321c0c",x"221409",x"4c2b16",x"2d1e14",x"453c32",x"150e07",x"150e07",x"150e07",x"150e07",x"231309",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2015",x"27190e",x"20170f",x"20170f",x"000000",x"4b372b",x"4b372b",x"341d0d",x"231409",x"231509",x"221409",x"201309",x"201308",x"150e07",x"26160a",x"26160a",x"2a180b",x"27160a",x"221409",x"261509",x"241509",x"28170a",x"25150a",x"26160a",x"1d1108",x"201309",x"231409",x"231409",x"221409",x"221409",x"24150a",x"24150a",x"27160a",x"221409",x"25160a",x"2a180b",x"27170a",x"241509",x"251509",x"221409",x"25150a",x"24150a",x"25160a",x"27170b",x"2b190c",x"29180b",x"231509",x"1f1208",x"201309",x"1c1108",x"251509",x"201208",x"1f1208",x"1d1108",x"221409",x"221409",x"25160a",x"1d1108",x"201309",x"1c1108",x"191008",x"1b1008",x"321b0b",x"150e07",x"755335",x"735135",x"5c3d24",x"785739",x"836140",x"846143",x"815d40",x"805e40",x"866343",x"866243",x"886545",x"826041",x"846042",x"8d6849",x"815f43",x"866445",x"8a6646",x"836041",x"805d3f",x"866343",x"846041",x"825e40",x"836041",x"78573b",x"815f41",x"876343",x"7e5d3e",x"78563a",x"79573b",x"7d5a3c",x"7c593c",x"775639",x"745236",x"6d4c32",x"5a3c22",x"775638",x"7e5d3e",x"7f5e40",x"7e5c3f",x"7f5d3f",x"856243",x"826041",x"846243",x"876244",x"835f41",x"946e4c",x"856245",x"8a6747",x"886445",x"876243",x"856141",x"8b6746",x"8a6545",x"8a6445",x"876343",x"615043",x"615043",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"492a13",x"492a13",x"39200f",x"351e0d",x"311c0c",x"2f1b0c",x"150e07",x"150e07",x"1d1108",x"2a180a",x"150e07",x"311b0b",x"2a180a",x"281609",x"2f1a0a",x"351d0b",x"391f0d",x"391f0d",x"2e190a",x"3c210e",x"351d0b",x"361e0e",x"3c210f",x"3c220f",x"3b210e",x"39200e",x"351d0d",x"371e0d",x"311b0b",x"391f0d",x"371e0d",x"3a200e",x"3c220f",x"3e230f",x"3c220f",x"432712",x"422611",x"3f2411",x"412511",x"402511",x"422612",x"412511",x"3b2210",x"3d2310",x"412511",x"371f0e",x"3d2310",x"3f2410",x"3b210f",x"3a210f",x"3e2310",x"3c220f",x"3d220f",x"3c220f",x"3f2410",x"3f2310",x"402511",x"3f2411",x"39200e",x"3a1f0e",x"371e0d",x"381e0d",x"361d0c",x"351d0c",x"371d0c",x"371e0c",x"3c210f",x"3c2210",x"432612",x"482914",x"462913",x"402511",x"3d2311",x"442713",x"3f2310",x"3f2410",x"402410",x"3c220f",x"3f2310",x"361e0d",x"351d0d",x"170f07",x"150e07",x"2c190b",x"341d0c",x"150e07",x"422511",x"3f2310",x"372b22",x"4e2d15",x"3c210f",x"3f2310",x"432611",x"432712",x"3a200e",x"3d210f",x"391f0d",x"39200f",x"3b2210",x"3d220f",x"3f2410",x"402411",x"3f2410",x"3f2411",x"3b210f",x"3d2310",x"3d210f",x"3e220f",x"412410",x"3d2310",x"321b0b",x"3a200d",x"301a0a",x"301b0b",x"311b0b",x"281609",x"2a1709",x"2c180a",x"341d0c",x"3a200d",x"341c0b",x"311b0b",x"2d190a",x"381f0d",x"39200e",x"38200e",x"39210e",x"361f0c",x"2d1a0b",x"170f07",x"321b0b",x"2a170a",x"2a180a",x"321c0c",x"381f0d",x"381f0e",x"39200f",x"361f0e",x"311c0d",x"351f0e",x"3a2210",x"3a2110",x"3a210f",x"3a210f",x"3d2310",x"3c2310",x"402410",x"402411",x"452712",x"412511",x"422511",x"412510",x"3f2410",x"432611",x"412511",x"442711",x"3e220f",x"432611",x"3c220f",x"27170a",x"27170a",x"301e12",x"301e12",x"3a2314",x"3a2212",x"3c2313",x"382010",x"341e0f",x"2d1b0d",x"1b1109",x"39200f",x"4e3d30",x"472915",x"412715",x"3a2312",x"412715",x"402614",x"2a190c",x"543015",x"91694b",x"855c40",x"966c4d",x"9d7453",x"92694a",x"8e6547",x"8b6547",x"8d6448",x"8d694c",x"885f42",x"926a4b",x"93694a",x"8c6448",x"6c4a34",x"886245",x"8e6547",x"7d583f",x"8e674a",x"815c40",x"7e5a3f",x"7b543a",x"7e583d",x"7d573c",x"67442f",x"78543b",x"7d573d",x"865e42",x"815a3f",x"735035",x"8b6345",x"815a3f",x"886244",x"865e42",x"785239",x"835c41",x"7a543a",x"7c573d",x"765238",x"7e5a3f",x"6e4c35",x"553b28",x"473221",x"473221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4a4138",x"4a4138",x"3b3129",x"4b2f1c",x"4b2f1c",x"311b0b",x"150e07",x"150e07",x"150e07",x"492913",x"3e2410",x"361f0e",x"39200e",x"3d230f",x"2d1609",x"361e0d",x"321b0b",x"351d0c",x"381f0e",x"321b0c",x"1c1108",x"815d41",x"7c573c",x"7a563c",x"7a553a",x"876145",x"886144",x"704d34",x"6e4c34",x"866042",x"8a6245",x"6c462e",x"865f43",x"835d42",x"825b3f",x"866145",x"7e593e",x"8b6345",x"825b40",x"805a3e",x"79583f",x"785339",x"8e6749",x"805c41",x"875f41",x"855e42",x"8f6749",x"815a40",x"886143",x"876144",x"91684a",x"8b6244",x"7b553b",x"7d583d",x"77533a",x"6e4a31",x"79563b",x"5c402c",x"412d1d",x"422e1e",x"422e1e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543622",x"543622",x"412310",x"361e0d",x"301a0b",x"351c0c",x"391f0d",x"3b200e",x"3c210e",x"351d0c",x"381e0c",x"3d220f",x"482812",x"2a180a",x"452610",x"452610",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"331d0d",x"2f1b0b",x"150e07",x"150e07",x"261509",x"24150a",x"150e07",x"261509",x"271509",x"150e07",x"482916",x"2d2018",x"4b4238",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2015",x"281a0f",x"201710",x"201710",x"000000",x"4e392c",x"4e392c",x"341d0d",x"211409",x"1e1208",x"241509",x"27170b",x"211409",x"150e07",x"28170b",x"27160a",x"29170b",x"29170a",x"251509",x"27160a",x"27160a",x"27160a",x"241509",x"231409",x"26160a",x"25160a",x"25150a",x"201309",x"1c1108",x"201309",x"241509",x"27170b",x"211409",x"26160a",x"231409",x"29170a",x"24150a",x"29180b",x"26160a",x"24150a",x"26160a",x"2a190b",x"27160a",x"26160a",x"251509",x"1d1108",x"26160a",x"1f1209",x"211308",x"1c1108",x"201308",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1f1208",x"1d1108",x"1b1108",x"150e07",x"1c1108",x"1d1108",x"150e07",x"331c0b",x"150e07",x"7c5a3d",x"856041",x"876445",x"846244",x"8e6c4a",x"8b6748",x"846042",x"866344",x"826041",x"846142",x"835f41",x"7f5b3d",x"7e5b3d",x"815e41",x"7a583c",x"836041",x"815f40",x"825f42",x"7d5c3f",x"7e5d3f",x"846143",x"805d40",x"7e5c3f",x"7b5a3d",x"805e41",x"825f42",x"66452b",x"745437",x"7c5a3c",x"815e41",x"78583b",x"815f41",x"7f5c3f",x"7c593c",x"866445",x"8d6949",x"896748",x"856345",x"805d40",x"815f41",x"846142",x"825f41",x"805d40",x"815d3e",x"845f40",x"846142",x"815d40",x"846041",x"815f41",x"836041",x"856244",x"846143",x"8a6545",x"876344",x"866244",x"5b4c40",x"5b4c40",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4c2b14",x"4c2b14",x"3a200e",x"3b210f",x"361e0d",x"28170a",x"150e07",x"1a1008",x"28160a",x"271609",x"231409",x"2c190a",x"311b0b",x"2c180a",x"2e190a",x"331c0b",x"391f0d",x"361e0c",x"2c190a",x"391f0d",x"361e0c",x"341c0c",x"341c0c",x"3b210f",x"361e0d",x"361d0c",x"351d0c",x"381e0d",x"3a200d",x"39200d",x"381f0d",x"391f0d",x"3b200e",x"3c210f",x"3a210f",x"39200f",x"371f0e",x"412411",x"412511",x"3a210f",x"39200f",x"3f2410",x"3f2410",x"3d2310",x"3e230f",x"3b210f",x"371e0d",x"361e0d",x"331d0d",x"3b220f",x"3b220f",x"361d0c",x"371d0c",x"3b220f",x"3c210f",x"3f2410",x"3c220f",x"3a200e",x"3b210f",x"3d220f",x"3b200e",x"3c210f",x"381f0d",x"361d0c",x"331c0c",x"3c210e",x"3c220f",x"3d220f",x"412411",x"3b200e",x"3d220f",x"3f2310",x"3c220f",x"3c210f",x"39200e",x"391f0d",x"3c210e",x"381f0d",x"3a200e",x"39200e",x"2f1a0b",x"150e07",x"1e1208",x"2e1a0b",x"331c0d",x"211409",x"3f2410",x"3b200e",x"34261c",x"4a2912",x"402410",x"3b200e",x"3c210e",x"3e2310",x"3d210f",x"412411",x"3e220f",x"3c210f",x"3a200f",x"3d220f",x"391f0d",x"3e2310",x"402310",x"3c220f",x"3c220f",x"3d220f",x"40230f",x"3d220f",x"3c210f",x"3e220e",x"351d0b",x"3b200d",x"341d0c",x"3a200d",x"331c0b",x"301a0a",x"301a0a",x"2f1a0a",x"381f0d",x"3a200d",x"301a0a",x"3b200e",x"311b0b",x"381f0d",x"3a210e",x"39200e",x"381f0d",x"361e0d",x"381f0d",x"381f0d",x"381f0d",x"3a200e",x"391f0d",x"39200e",x"39200d",x"3b210f",x"39200e",x"3f2310",x"402410",x"3b220f",x"3f2410",x"3c220f",x"3c2210",x"3d2310",x"3b220f",x"3b210f",x"3e230f",x"3f2310",x"3f240f",x"391f0e",x"3f2310",x"422611",x"402410",x"402410",x"371d0c",x"3e220f",x"3f230f",x"432611",x"402410",x"2f1b0c",x"2f1b0c",x"311f13",x"311f13",x"3a2314",x"3c2414",x"3c2313",x"3b2212",x"341f10",x"2c1a0d",x"180f07",x"38200e",x"533e30",x"462916",x"422816",x"3a2312",x"472b17",x"3a2211",x"2d1b0d",x"6a472f",x"8c674a",x"835b3f",x"815b3f",x"835e43",x"865e42",x"886145",x"815a3f",x"674731",x"7b5a41",x"7d573c",x"896347",x"8d684a",x"805b41",x"755339",x"805b40",x"7a543b",x"825e43",x"835e42",x"855e43",x"805b3f",x"785339",x"7a563a",x"765139",x"754f36",x"845f43",x"7e593e",x"725037",x"785439",x"5f3d27",x"79573d",x"6d4b34",x"7c583e",x"7f593f",x"765137",x"785339",x"7a563c",x"795539",x"765238",x"78543a",x"684932",x"553c29",x"422f1f",x"422f1f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"52483e",x"52483e",x"3f352b",x"4e2d18",x"4e2d18",x"271609",x"150e07",x"150e07",x"150e07",x"482811",x"3a210f",x"351e0e",x"331c0c",x"361f0d",x"241208",x"301a0b",x"371e0d",x"341c0b",x"3f230f",x"3d210e",x"1b1108",x"5e412e",x"735138",x"78543c",x"77553b",x"7c573d",x"714f36",x"78543a",x"715036",x"765138",x"845f43",x"704d35",x"76533a",x"77563c",x"7f5b40",x"7f5d42",x"704d36",x"805d41",x"78543a",x"7b573d",x"7c583e",x"77543a",x"7e593e",x"866246",x"805b3f",x"815c40",x"825e42",x"6c4c35",x"684833",x"78553c",x"6f4d36",x"76533b",x"7b553a",x"734f37",x"6d4c35",x"5b3d27",x"5c3d2b",x"5c402c",x"3e2b1c",x"3d2a1b",x"3d2a1b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50331f",x"50331f",x"412410",x"381f0d",x"381f0d",x"381f0d",x"331b0b",x"381f0d",x"3b200e",x"391f0e",x"371d0c",x"432611",x"472811",x"321c0c",x"553319",x"503017",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"2d190c",x"26160a",x"150e07",x"150e07",x"231509",x"211409",x"150e07",x"2e190b",x"251509",x"201309",x"472815",x"2f2118",x"4a4138",x"150e07",x"150e07",x"150e07",x"150e07",x"211208",x"150e07",x"150e07",x"150e07",x"150e07",x"322116",x"24170e",x"201810",x"201810",x"000000",x"48372b",x"48372b",x"341e0d",x"211409",x"1c1108",x"211409",x"211409",x"201309",x"150e07",x"231409",x"231409",x"27160a",x"27160a",x"29170a",x"28170a",x"27160a",x"27160a",x"25150a",x"231409",x"29180b",x"28170a",x"241509",x"231409",x"211409",x"1e1208",x"1d1108",x"1e1208",x"1f1208",x"241509",x"251509",x"241509",x"1f1208",x"221409",x"231409",x"211409",x"25150a",x"25160a",x"28170a",x"2a180b",x"28170a",x"241509",x"231509",x"251509",x"1f1208",x"1a1008",x"1a1008",x"1a1008",x"201308",x"201308",x"1d1108",x"1c1108",x"1f1309",x"1a1008",x"231409",x"1c1108",x"1d1208",x"1c1108",x"371e0d",x"150e07",x"886547",x"876445",x"876444",x"886445",x"876446",x"876446",x"836041",x"846142",x"7e5d40",x"7a583b",x"876445",x"896647",x"896547",x"8a6648",x"856345",x"795a3c",x"816042",x"8a6648",x"8e6b4b",x"846244",x"8c6747",x"896546",x"846244",x"816041",x"8a6747",x"866343",x"825f3f",x"815f41",x"75563a",x"7f5d40",x"7f5e41",x"7e5e41",x"826143",x"7d5c40",x"886444",x"836042",x"866345",x"886546",x"815e40",x"836041",x"815e41",x"79583b",x"886547",x"8d6949",x"896547",x"8e6949",x"8d694a",x"8a6745",x"866445",x"8e694a",x"8e6b4b",x"866445",x"8e6949",x"926c4c",x"8c6849",x"584639",x"584639",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452611",x"452611",x"351e0d",x"381f0e",x"351e0d",x"251509",x"2a170a",x"28160a",x"170f07",x"221409",x"1a1008",x"2d190b",x"341d0c",x"361d0c",x"351d0c",x"391f0d",x"3b200e",x"311b0b",x"351d0c",x"2e190a",x"371e0d",x"351d0d",x"351d0c",x"381f0d",x"341c0c",x"331c0c",x"381e0d",x"331b0b",x"3a200d",x"391f0d",x"3b200e",x"3a200e",x"3c210f",x"402410",x"402411",x"412511",x"3a200e",x"3b210e",x"412511",x"3a210f",x"39200f",x"341d0c",x"321c0c",x"3f2410",x"3d2210",x"341c0c",x"311b0b",x"301a0b",x"2e190b",x"2f1a0b",x"2e190b",x"2c180a",x"361e0d",x"361e0d",x"381f0e",x"3b210f",x"381e0d",x"331c0c",x"331c0c",x"321b0b",x"351b0b",x"331b0b",x"361d0d",x"361d0c",x"381e0c",x"311a0b",x"361e0d",x"3d210e",x"3b200e",x"3c210e",x"3a200e",x"3c210f",x"391f0d",x"391f0d",x"371f0e",x"39200e",x"3b210e",x"3b210e",x"351c0c",x"361d0c",x"28160a",x"2a170a",x"2a170a",x"241509",x"29170a",x"211308",x"3c210e",x"341c0c",x"30251d",x"3d200d",x"371e0c",x"391f0e",x"3a200e",x"3b210e",x"391f0d",x"3a210f",x"3a210f",x"381f0e",x"381f0e",x"3c210f",x"402310",x"3a200e",x"39200e",x"3a200e",x"3a200e",x"361e0d",x"3c220e",x"3c220f",x"38200e",x"39200e",x"3f2411",x"3b210f",x"371f0e",x"3e2310",x"3a210f",x"39200e",x"3b210e",x"3b210f",x"3a210f",x"39200e",x"371e0d",x"3b200e",x"3b200e",x"3c220f",x"381f0e",x"361d0c",x"351c0c",x"321b0b",x"3a200e",x"3b200f",x"3a200e",x"371d0c",x"381f0e",x"3e230f",x"3c220f",x"3a200e",x"361d0c",x"341c0b",x"361d0c",x"361e0d",x"381f0d",x"3f220f",x"3e230f",x"3d220f",x"3c220f",x"3c220f",x"3d220f",x"412310",x"3a200e",x"381e0c",x"391f0d",x"3a200d",x"381e0d",x"341c0c",x"3b200e",x"3d210f",x"412410",x"3f230f",x"3c210f",x"29170a",x"29170a",x"342014",x"342014",x"362011",x"3c2514",x"3d2414",x"3c2312",x"341f10",x"2b190c",x"180f07",x"38200e",x"503e30",x"482a17",x"382313",x"3d2413",x"462b18",x"3b2212",x"2f1c0e",x"472e1e",x"674934",x"63442f",x"6a4b34",x"6c4d36",x"634630",x"6c4d35",x"6b4c34",x"644631",x"6b4e37",x"684932",x"6b4d36",x"6c4e37",x"6d4e37",x"684933",x"644732",x"5c402c",x"60422d",x"674933",x"6f5139",x"694a32",x"5f422c",x"64452f",x"60422d",x"573a26",x"694a34",x"60432d",x"624530",x"593f2a",x"4a2e1d",x"5a3e2a",x"482f1f",x"634630",x"5e412b",x"61442e",x"5c3f2a",x"5f422d",x"5d412c",x"5a3e2a",x"5b402c",x"4c3624",x"372619",x"1d140d",x"1d140d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4f463d",x"4f463d",x"322821",x"4f2c14",x"4f2c14",x"271509",x"150e07",x"150e07",x"150e07",x"482711",x"3a220f",x"361e0d",x"311b0c",x"361e0d",x"2e190a",x"361e0d",x"3b200e",x"341c0c",x"3d220f",x"3d220f",x"1e1208",x"593e2b",x"593e2b",x"654934",x"5d422e",x"5e412d",x"593f2b",x"63442f",x"60422d",x"63442e",x"674833",x"62442e",x"6a4c35",x"5e432e",x"664832",x"6c4d36",x"5f422c",x"684a33",x"62432d",x"5e432d",x"61442e",x"674731",x"6a4a34",x"72513a",x"694a33",x"674932",x"684932",x"694a33",x"6e4f36",x"6c4d36",x"715138",x"5f412d",x"543826",x"674832",x"573c27",x"43281c",x"472e1f",x"45301f",x"1a1109",x"20150c",x"20150c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584e44",x"584f44",x"4f3422",x"41240f",x"3b200e",x"402410",x"3a200e",x"2f190b",x"331c0b",x"381f0d",x"3b210e",x"351c0c",x"432612",x"4a2a13",x"5d5349",x"584e44",x"574d43",x"564d42",x"564d42",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"211309",x"1e1208",x"150e07",x"231309",x"150e07",x"201308",x"452714",x"322116",x"494037",x"150e07",x"150e07",x"150e07",x"150e07",x"221208",x"150e07",x"150e07",x"150e07",x"150e07",x"301f14",x"2a1a0f",x"201811",x"201811",x"000000",x"50392a",x"50392a",x"301c0c",x"1e1208",x"221409",x"2b190b",x"1a1008",x"211409",x"150e07",x"1e1208",x"26160a",x"221409",x"241409",x"261509",x"221409",x"251509",x"231409",x"251509",x"201308",x"221409",x"201309",x"231409",x"211308",x"1f1208",x"1d1108",x"201208",x"1c1108",x"1e1208",x"1e1208",x"211309",x"231409",x"25150a",x"211309",x"25150a",x"221409",x"1e1208",x"241509",x"251509",x"28170a",x"28170a",x"25150a",x"221309",x"211309",x"1d1108",x"211309",x"1f1208",x"211309",x"1f1208",x"241509",x"1f1208",x"221409",x"201309",x"1d1208",x"201309",x"1e1208",x"150e07",x"1c1108",x"381f0d",x"150e07",x"886546",x"836144",x"896646",x"8e6b4a",x"8d6b4b",x"8c694a",x"836143",x"866443",x"846142",x"856141",x"836041",x"846142",x"815f40",x"815e3f",x"805d3e",x"7d5b3d",x"7a593c",x"7b593c",x"775538",x"7e5b3e",x"7f5b3e",x"825f40",x"876343",x"825f40",x"805d3f",x"7f5e41",x"7a593c",x"76563a",x"79593c",x"78573c",x"7c5c40",x"79593e",x"76573c",x"816042",x"866445",x"8d6a49",x"8a6749",x"8d6a49",x"876445",x"886444",x"866242",x"835f41",x"856242",x"846142",x"846142",x"815e3f",x"815d3f",x"815d3f",x"79573b",x"815d3f",x"7c5a3c",x"79573b",x"77563a",x"836140",x"8b6746",x"5d493b",x"5d493b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452510",x"452510",x"311b0c",x"361e0d",x"1c1108",x"201309",x"2e190b",x"2d190a",x"150e07",x"2b180a",x"190f07",x"331c0c",x"371e0d",x"361e0d",x"3a200d",x"351d0c",x"2f190a",x"351d0c",x"301a0b",x"361e0d",x"321b0b",x"311b0c",x"38200e",x"371e0d",x"371e0c",x"331b0b",x"351b0b",x"341c0c",x"3b200d",x"351d0d",x"3a200e",x"3f2310",x"3f2410",x"3f2310",x"402410",x"39200e",x"3b210f",x"3f2410",x"39200e",x"371f0e",x"3a200f",x"3a210f",x"37200f",x"39210f",x"3a210f",x"371f0e",x"341c0c",x"301a0b",x"2d180a",x"2f180a",x"2c170a",x"2a170a",x"351d0d",x"381f0e",x"3b200e",x"3c220f",x"412411",x"3a210e",x"38200e",x"3a200e",x"39200e",x"39200e",x"3f230f",x"412511",x"3d2410",x"432711",x"432611",x"412511",x"432611",x"422611",x"402410",x"39200e",x"391f0d",x"361e0d",x"391f0d",x"3a200e",x"3d220f",x"3a200e",x"3a200e",x"331d0c",x"191008",x"2f1a0b",x"2a170a",x"150e07",x"28160a",x"241409",x"3e230f",x"39200e",x"33251b",x"432410",x"3d220f",x"381f0e",x"3a200e",x"452914",x"3f2411",x"361e0d",x"361f0e",x"150e07",x"4a2a13",x"321c0c",x"170f07",x"3a200e",x"39200e",x"3a200e",x"3a200e",x"361e0d",x"3c220e",x"3c220f",x"38200e",x"39200e",x"3f2411",x"3b210f",x"371f0e",x"3e2310",x"3a210f",x"39200e",x"3b210e",x"3b210f",x"3a210f",x"321c0b",x"2d190b",x"261509",x"1c1108",x"241509",x"25160a",x"24150a",x"241409",x"221308",x"1e1108",x"29160a",x"2a180a",x"361d0d",x"351d0d",x"351d0d",x"321c0c",x"321c0d",x"361e0e",x"26150a",x"27160a",x"2e1b0b",x"2a190b",x"28170a",x"25150a",x"25160a",x"27160a",x"301c0c",x"361f0e",x"3c200e",x"221409",x"180f08",x"150e07",x"40230f",x"351d0d",x"361d0c",x"3f2310",x"3f230f",x"432711",x"381f0d",x"3f230f",x"25150a",x"25150a",x"352114",x"352114",x"382313",x"3b2414",x"402615",x"3c2312",x"331e0f",x"29170b",x"180f07",x"3d2310",x"4e3f34",x"4a2c17",x"3f2613",x"362012",x"3a2314",x"392111",x"28180b",x"483020",x"5c412d",x"593e2a",x"5b412d",x"5e432e",x"583d2a",x"5d422d",x"5a3f2b",x"5a3f2b",x"5f442f",x"5d412c",x"5d432e",x"61442f",x"614530",x"593e2b",x"5d412d",x"5a3f2b",x"5c402b",x"5c412d",x"614530",x"5d412c",x"573c28",x"593e29",x"533a26",x"47301f",x"5a3f2b",x"513825",x"533a28",x"4f3724",x"462e1e",x"4c3322",x"483020",x"543a28",x"533a27",x"4e3524",x"493221",x"493221",x"4b3322",x"48311f",x"453020",x"3a281a",x"18110a",x"1a130c",x"1a130c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4f463c",x"4f463c",x"382f27",x"4d2d17",x"4d2d17",x"2c170a",x"150e07",x"150e07",x"150e07",x"482812",x"382110",x"2e1a0c",x"311c0c",x"311b0c",x"301a0b",x"331c0c",x"3c220f",x"321c0c",x"3d230f",x"381f0e",x"191008",x"453123",x"4a3525",x"4c3625",x"453120",x"493322",x"473020",x"483120",x"493220",x"4c3422",x"4e3625",x"4b3322",x"493323",x"473120",x"4e3726",x"523a27",x"473221",x"503826",x"503725",x"4c3524",x"4a3422",x"513825",x"543c29",x"553c29",x"4e3624",x"523927",x"533a27",x"503725",x"553b28",x"624530",x"583d2a",x"523927",x"4f3724",x"493121",x"442e1e",x"3e271a",x"3d291a",x"2e1f13",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"55483d",x"55483d",x"584e44",x"584f44",x"4c301d",x"40230f",x"371e0d",x"402411",x"361e0d",x"331b0b",x"361c0c",x"3b200e",x"3e220f",x"341b0b",x"412511",x"4a2912",x"574d43",x"5a5046",x"594d42",x"675142",x"675142",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"1b1108",x"231409",x"150e07",x"150e07",x"28160a",x"150e07",x"271509",x"492915",x"2f2015",x"463c32",x"150e07",x"150e07",x"150e07",x"150e07",x"241409",x"150e07",x"150e07",x"150e07",x"150e07",x"322114",x"2b1b10",x"221810",x"221810",x"000000",x"523929",x"523929",x"331d0d",x"1c1108",x"211409",x"231409",x"1d1208",x"211409",x"150e07",x"241509",x"1e1208",x"251509",x"26150a",x"251509",x"261509",x"231409",x"241509",x"241409",x"221409",x"201309",x"1f1309",x"211409",x"231409",x"180f07",x"1d1108",x"201208",x"221409",x"180f07",x"191008",x"1b1108",x"211308",x"211309",x"221409",x"201208",x"1a1008",x"211309",x"251509",x"241509",x"26160a",x"211309",x"221409",x"221409",x"241509",x"241509",x"231409",x"201308",x"201308",x"251509",x"251509",x"1f1208",x"251509",x"1a1008",x"1d1108",x"1d1208",x"201309",x"1b1108",x"150e07",x"2e1a0b",x"150e07",x"7f5c3e",x"76563a",x"7b593c",x"825e41",x"7b593b",x"825f41",x"7e5c3e",x"7c593c",x"7f5c3e",x"79573a",x"7a583b",x"6e4f35",x"7a593c",x"7e5b3e",x"825f41",x"815e41",x"825f41",x"836041",x"815e41",x"815d3f",x"836042",x"805d3e",x"7d5b3d",x"846243",x"7a5b3e",x"816143",x"826143",x"826043",x"866345",x"7f5d3f",x"7d5d40",x"7b5a3d",x"77563a",x"745438",x"7a583c",x"7c5a3d",x"765639",x"7d5b3e",x"7c593c",x"815d3f",x"825e40",x"785639",x"7a583b",x"78573b",x"825f40",x"835f41",x"866243",x"866243",x"846042",x"856243",x"886444",x"7f5d3e",x"7f5d40",x"825e40",x"815e3f",x"5a4537",x"5a4537",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2913",x"4a2913",x"3b210f",x"2f1b0c",x"341d0d",x"251409",x"321d0d",x"341d0d",x"2e1a0a",x"311b0b",x"2d190b",x"2c180a",x"301a0a",x"2a1709",x"331c0b",x"341d0c",x"371e0d",x"2c180a",x"381f0d",x"341c0c",x"39200e",x"39200e",x"341c0c",x"39200d",x"371e0c",x"32190b",x"381e0c",x"371d0c",x"3c210e",x"3c210e",x"3c220f",x"3e230f",x"3f2310",x"3a200e",x"341c0c",x"381e0d",x"381f0e",x"361e0d",x"3a200e",x"361e0d",x"381f0e",x"3b210f",x"3c210f",x"381f0e",x"3e220f",x"3e2310",x"381f0e",x"361e0d",x"341d0d",x"3a210f",x"3c220f",x"351d0d",x"381f0e",x"361e0d",x"381f0d",x"331c0b",x"381f0d",x"341d0c",x"331c0c",x"3b200e",x"361d0d",x"341c0c",x"3a200d",x"3e220e",x"3f230f",x"3f2310",x"3e230f",x"402410",x"422611",x"432612",x"442712",x"412411",x"3e220f",x"391f0d",x"361c0c",x"331b0b",x"351c0c",x"331c0c",x"361e0d",x"341c0c",x"2c180b",x"2d180a",x"2d180a",x"2a160a",x"2e190a",x"251509",x"391f0e",x"351d0d",x"34281e",x"412410",x"3b210f",x"39200e",x"361e0d",x"412612",x"3e2411",x"361e0d",x"39200f",x"150e07",x"492813",x"150e07",x"221409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f2f2f",x"2f2f2f",x"323232",x"323232",x"343434",x"323232",x"313232",x"323232",x"2a2a2a",x"2d2d2d",x"323232",x"313131",x"323232",x"222222",x"343434",x"323232",x"292929",x"404040",x"343434",x"303030",x"2f2f2f",x"313131",x"2f2f2f",x"303030",x"2d2d2d",x"323232",x"303030",x"2b2726",x"2b2726",x"3e220f",x"221409",x"5f4b3e",x"150e07",x"482913",x"3b210e",x"381f0d",x"402310",x"422611",x"452813",x"391f0d",x"402410",x"2d190b",x"2d190b",x"362215",x"362215",x"382213",x"3b2314",x"402715",x"3b2312",x"331d0f",x"29170c",x"180f07",x"452812",x"493b30",x"4a2c17",x"3c2414",x"402615",x"442916",x"321d0f",x"311c0d",x"311c0d",x"5c412d",x"593e2a",x"5b412d",x"5e432e",x"583d2a",x"5d422d",x"5a3f2b",x"5a3f2b",x"5f442f",x"5d412c",x"5d432e",x"61442f",x"614530",x"593e2b",x"5d412d",x"5a3f2b",x"5c402b",x"5c412d",x"614530",x"5d412c",x"573c28",x"593e29",x"533a26",x"47301f",x"5a3f2b",x"513825",x"533a28",x"4f3724",x"462e1e",x"4c3322",x"483020",x"543a28",x"533a27",x"4e3524",x"493221",x"493221",x"4b3322",x"48311f",x"453020",x"3a281a",x"18110a",x"1a130c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"544a40",x"544a40",x"51483f",x"553928",x"553928",x"2d180a",x"150e07",x"150e07",x"150e07",x"452711",x"442813",x"3b2210",x"301c0c",x"361e0d",x"301a0b",x"361d0d",x"3a200e",x"381e0d",x"301b0c",x"361e0d",x"201309",x"654a32",x"634931",x"6d5037",x"654a32",x"6b4d35",x"6f5138",x"7a5a3e",x"7a593c",x"7a583c",x"836244",x"7b5b3f",x"7f5d41",x"825f41",x"816043",x"826042",x"876446",x"815e40",x"876445",x"7f5c3d",x"815e3f",x"8c6847",x"906b4a",x"8c6848",x"876244",x"8e6a4b",x"866244",x"886648",x"815d40",x"856444",x"815e42",x"815e41",x"866346",x"846345",x"805d42",x"73553a",x"5e442d",x"6e5138",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d332a",x"3d332a",x"594f45",x"584e43",x"6a5647",x"40230f",x"391f0d",x"3f2410",x"3d220f",x"361c0c",x"351d0b",x"3b200d",x"3a200e",x"30190a",x"3d220f",x"4b2b13",x"524940",x"413930",x"44372d",x"4e3526",x"4e3526",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"29170b",x"150e07",x"2f1b0c",x"492915",x"312318",x"463c33",x"150e07",x"150e07",x"150e07",x"150e07",x"261509",x"150e07",x"150e07",x"150e07",x"170f07",x"301f14",x"2a1b11",x"221810",x"221810",x"000000",x"503829",x"503829",x"361f0e",x"1f1208",x"221409",x"2b180b",x"221409",x"1d1108",x"150e07",x"211208",x"221309",x"251509",x"231409",x"1e1208",x"201208",x"221308",x"221308",x"211308",x"221409",x"241409",x"211309",x"1f1208",x"241409",x"201208",x"1e1208",x"211309",x"26160a",x"211409",x"1a1008",x"201309",x"1e1208",x"221409",x"1f1208",x"241509",x"201208",x"211308",x"28160a",x"25160a",x"29170a",x"29170a",x"28170a",x"231409",x"1f1309",x"251509",x"1e1208",x"231409",x"271609",x"211308",x"1e1208",x"1e1108",x"231409",x"24150a",x"28180b",x"201309",x"1e1208",x"170f07",x"170f07",x"341c0c",x"150e07",x"8a6645",x"7e5c3e",x"805e40",x"7d5c3f",x"725237",x"7e5b3d",x"7d5c3e",x"7d5c3e",x"846144",x"815e41",x"846142",x"7e5c3f",x"7e5c3f",x"846245",x"886446",x"815e41",x"7d5b3d",x"7d5c3f",x"7e5c3f",x"7e5b3d",x"7e5b3d",x"815e41",x"846243",x"7a593d",x"7c5a3c",x"705037",x"745338",x"7d5b3d",x"7c5a3c",x"7d5c3e",x"815f41",x"826041",x"79583c",x"7a593c",x"7f5d3f",x"836042",x"7c5a3c",x"7d5a3c",x"836142",x"856242",x"8c6747",x"826041",x"835f42",x"876344",x"876243",x"866446",x"866345",x"815e41",x"815d3f",x"825f41",x"846043",x"815d3f",x"815d3f",x"846143",x"896544",x"594133",x"594133",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"41240f",x"41240f",x"351e0d",x"311b0c",x"341d0d",x"341d0d",x"321c0c",x"321d0d",x"361e0d",x"150e07",x"281609",x"301a0b",x"371e0c",x"301b0b",x"341c0b",x"351d0b",x"391f0d",x"301b0c",x"39200e",x"371f0d",x"391f0d",x"3a200e",x"341d0c",x"351d0c",x"351c0c",x"371e0c",x"391f0d",x"3d210e",x"381f0d",x"3a210f",x"3f2310",x"3c230f",x"3b210f",x"3e2310",x"3e2310",x"3f240f",x"361f0d",x"3f2410",x"3a210f",x"3c220f",x"3b210f",x"3a210f",x"3b210f",x"381f0d",x"351c0c",x"351c0c",x"381f0d",x"341d0d",x"371f0e",x"341e0d",x"371e0d",x"331c0d",x"321c0c",x"351d0d",x"381e0d",x"371e0d",x"391f0e",x"361e0d",x"331c0c",x"301a0b",x"371e0d",x"381e0c",x"341c0c",x"3a1f0e",x"3d210f",x"3a200e",x"3e220f",x"3d210f",x"3a200e",x"391f0d",x"3a200d",x"3c210e",x"3a200e",x"3d210e",x"391f0d",x"3a200e",x"3e220f",x"3e220f",x"39200e",x"3c220f",x"3a200e",x"351d0d",x"39200e",x"3f2410",x"150e07",x"331d0d",x"402410",x"3a200e",x"342b23",x"412410",x"38200e",x"381f0e",x"381f0d",x"3f2310",x"3c2310",x"361e0d",x"381f0e",x"150e07",x"452511",x"150e07",x"150e07",x"000000",x"000000",x"8c7559",x"8c7559",x"160f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"312a25",x"312a25",x"323232",x"343434",x"343434",x"343434",x"2d2d2d",x"323232",x"353535",x"313131",x"303030",x"323232",x"323333",x"333333",x"2c2d2d",x"2f2f2f",x"313131",x"333333",x"2f2f2f",x"2f2f2f",x"323232",x"313131",x"2f2f2f",x"2f2f2f",x"292929",x"2a2a2a",x"282828",x"292929",x"292929",x"000000",x"543d2d",x"543d2d",x"150e07",x"3e220f",x"371e0d",x"3b200e",x"3d220f",x"412511",x"412511",x"3a200e",x"3f230f",x"2a180b",x"2a180b",x"362215",x"362215",x"392213",x"3d2413",x"412815",x"3b2211",x"331d0f",x"2b190c",x"190f08",x"3b200f",x"483b31",x"492b16",x"472a16",x"3c2513",x"3a2415",x"3c2312",x"27170b",x"27170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"5a5146",x"5a5146",x"584e44",x"52483e",x"52483e",x"3d210f",x"150e07",x"150e07",x"150e07",x"3e210f",x"3c2310",x"3e2410",x"331d0d",x"311b0c",x"2f1a0b",x"351e0d",x"39200e",x"321b0b",x"3f2410",x"331c0c",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"231608",x"251709",x"150e07",x"150e07",x"1a1107",x"1f1408",x"1e1308",x"211508",x"251709",x"231608",x"221608",x"1f1408",x"1b1108",x"1b1108",x"191007",x"191007",x"1f1408",x"1a1107",x"180f07",x"1c150c",x"23180d",x"1f160d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574d42",x"574d42",x"574d43",x"584d42",x"594132",x"40230f",x"3d220f",x"381f0e",x"3b210e",x"3a1f0d",x"371e0c",x"3c200e",x"3b200e",x"361c0b",x"3d220f",x"4c2b14",x"463d34",x"393028",x"3e2f25",x"4b3323",x"4b3323",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"190f07",x"150e07",x"150e07",x"2e190b",x"150e07",x"311c0d",x"472916",x"35271d",x"473e34",x"150e07",x"150e07",x"150e07",x"150e07",x"28170a",x"150e07",x"150e07",x"150e07",x"1a1008",x"332014",x"2f1d11",x"221810",x"221810",x"000000",x"4d382b",x"4d382b",x"301b0c",x"241509",x"28170b",x"231409",x"27170b",x"211409",x"150e07",x"25160a",x"27160a",x"25150a",x"25150a",x"27160a",x"241509",x"27160a",x"28170b",x"28170a",x"25150a",x"231409",x"241509",x"251509",x"241509",x"24150a",x"26160a",x"25160a",x"27160a",x"211309",x"241509",x"221309",x"1d1108",x"1f1208",x"170f07",x"190f07",x"1a0f07",x"1b0f07",x"231409",x"27160a",x"26160a",x"25150a",x"27160a",x"211309",x"1f1208",x"26160a",x"251509",x"251509",x"170f07",x"231409",x"251509",x"1f1208",x"1d1108",x"1f1309",x"211409",x"24150a",x"211409",x"231409",x"150e07",x"2b180a",x"150e07",x"8b6748",x"866345",x"8b6849",x"836144",x"795a3e",x"846245",x"78573b",x"765639",x"765639",x"805b3e",x"846041",x"856243",x"836244",x"866143",x"886647",x"846244",x"805f42",x"896647",x"7f5c40",x"7f5d40",x"7c5b3e",x"826143",x"7f5d3f",x"79583c",x"7e5d3f",x"79583b",x"79593c",x"8c6747",x"826143",x"886647",x"856243",x"846141",x"846244",x"876446",x"8b6748",x"7e5d41",x"846244",x"876446",x"78573b",x"735337",x"765639",x"7d5a3c",x"886545",x"856243",x"886647",x"866143",x"7a5a3f",x"846244",x"906b4b",x"896647",x"825e41",x"846143",x"896545",x"8a6748",x"846142",x"4f3c2f",x"4f3c2f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"432611",x"432611",x"39200e",x"311b0c",x"351e0d",x"331d0d",x"331d0d",x"39200f",x"3a200e",x"201309",x"341d0d",x"351d0d",x"381f0e",x"371e0d",x"381f0e",x"371f0e",x"2f190b",x"3c220f",x"3b200e",x"3a200e",x"402410",x"402410",x"3f2310",x"3b210e",x"3f230f",x"3c210e",x"3a200e",x"3b200d",x"3b200e",x"391f0d",x"381f0e",x"361e0d",x"361e0d",x"3d230f",x"432612",x"3c210f",x"3c210f",x"381f0e",x"331c0c",x"39200e",x"3a210e",x"3c220f",x"3a210f",x"3a210f",x"361e0d",x"361e0d",x"2f1a0b",x"341d0d",x"311b0c",x"331c0c",x"321c0c",x"301b0c",x"341d0d",x"331c0c",x"321a0b",x"321b0b",x"391f0d",x"391f0d",x"351c0c",x"311b0b",x"351d0c",x"3a200e",x"331c0c",x"412410",x"3f230f",x"3f2310",x"3a200e",x"3d220f",x"3c210e",x"361d0c",x"3e230f",x"3f2310",x"412511",x"402410",x"3b200e",x"3c210e",x"412410",x"3b210f",x"371f0e",x"39200e",x"39200e",x"3a210f",x"3c210f",x"3f2411",x"1c1108",x"301b0c",x"412310",x"381f0d",x"3d3027",x"462811",x"3b210f",x"3b200e",x"39200d",x"3f2411",x"361e0e",x"39200f",x"361e0d",x"150e07",x"42230f",x"150e07",x"150e07",x"000000",x"000000",x"8c7559",x"8c7559",x"160f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"303030",x"2e2e2e",x"2f2f2f",x"2f2f2f",x"282828",x"2f2f2f",x"2d2d2d",x"323232",x"313131",x"333333",x"2e2e2e",x"313131",x"343434",x"333333",x"333333",x"2e2e2e",x"313131",x"323232",x"333333",x"303030",x"323232",x"2c2c2c",x"2e2e2e",x"272727",x"2c2c2c",x"2c2c2c",x"000000",x"50392b",x"50392b",x"150e07",x"422511",x"381f0e",x"3b210e",x"3c220f",x"402410",x"422612",x"3c220f",x"3d230f",x"301c0c",x"301c0c",x"332013",x"332013",x"3c2514",x"3c2415",x"3f2513",x"3d2313",x"382011",x"2d1a0d",x"190f08",x"38200e",x"4b3b30",x"472916",x"422815",x"3f2514",x"452a17",x"331d0f",x"2d1a0d",x"2d1a0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"5c5247",x"5c5247",x"584e44",x"5a5046",x"5a5046",x"3d210f",x"150e07",x"150e07",x"412410",x"412410",x"3c2310",x"37200f",x"3b2210",x"2f1b0c",x"321c0c",x"351e0d",x"341d0d",x"331c0c",x"351e0d",x"361e0d",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"201508",x"291a09",x"241708",x"1d1208",x"221508",x"211508",x"201408",x"251708",x"291a09",x"2b1b09",x"281909",x"2d1c0a",x"2a1b09",x"231608",x"271909",x"221608",x"231608",x"211508",x"1c1208",x"1c1208",x"1c1208",x"1c1208",x"201408",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1a0b",x"2d1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574d42",x"574d42",x"534a40",x"4c4137",x"4a3223",x"3c210e",x"3b210f",x"402410",x"3a200e",x"3d220f",x"3c200d",x"3c200d",x"3c210e",x"321b0b",x"3a200e",x"452711",x"52483f",x"453c33",x"44362c",x"503729",x"503729",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"160f07",x"150e07",x"150e07",x"391f0d",x"150e07",x"2b180a",x"472a17",x"34261c",x"4c423a",x"150e07",x"150e07",x"150e07",x"150e07",x"29170b",x"150e07",x"150e07",x"150e07",x"150e07",x"321f12",x"281a10",x"231810",x"231810",x"000000",x"523b2d",x"523b2d",x"321c0c",x"231509",x"221409",x"201309",x"25160a",x"24150a",x"150e07",x"28170a",x"28170a",x"221409",x"26160a",x"27160a",x"2c190b",x"221409",x"26160a",x"25160a",x"26160a",x"251509",x"29170a",x"221409",x"221409",x"221409",x"221409",x"231409",x"26160a",x"251509",x"241509",x"27160a",x"26160a",x"26160a",x"27170a",x"25150a",x"24150a",x"25150a",x"241509",x"29170a",x"25150a",x"231409",x"241509",x"29180b",x"27160a",x"211309",x"201208",x"241509",x"25150a",x"221409",x"231409",x"25160a",x"25150a",x"201309",x"150e07",x"201309",x"201309",x"1e1208",x"1e1208",x"351c0c",x"150e07",x"8b6747",x"835f42",x"886546",x"866345",x"7e5d3f",x"715338",x"815f41",x"7c5a3b",x"775639",x"725234",x"775537",x"7f5c3d",x"846041",x"745437",x"8a6747",x"896647",x"846244",x"805e41",x"805e41",x"7e5c40",x"805d40",x"805e40",x"826043",x"846244",x"886446",x"826143",x"805f42",x"856142",x"876445",x"8a6749",x"836143",x"856244",x"856345",x"866243",x"8a6648",x"846244",x"825f41",x"805e40",x"886444",x"805c3e",x"7b593b",x"765536",x"7e5b3a",x"846041",x"815e3f",x"755438",x"886546",x"846244",x"866445",x"886546",x"896647",x"886344",x"8b6646",x"805d40",x"836143",x"473b31",x"473b31",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452611",x"452611",x"331c0c",x"2c180a",x"321b0b",x"311b0b",x"371e0d",x"37200e",x"3a210f",x"150e07",x"301c0d",x"361e0d",x"381f0d",x"331c0c",x"3e220f",x"3c220f",x"3f2310",x"412510",x"432511",x"472811",x"432510",x"432510",x"3f2310",x"412511",x"422511",x"3c210f",x"41240f",x"3f220e",x"432611",x"442712",x"412511",x"462812",x"432611",x"492a14",x"482a14",x"452712",x"3c220f",x"3b210e",x"3a210e",x"3d2310",x"412511",x"412511",x"3e230f",x"412410",x"432611",x"3a200e",x"39200e",x"381f0e",x"3b200e",x"39200e",x"381f0d",x"371e0d",x"371e0d",x"381f0d",x"3c210e",x"3e220f",x"391f0d",x"3b200d",x"391f0d",x"381e0d",x"361d0c",x"3b200d",x"351c0b",x"3b200d",x"3b200e",x"3b200d",x"3b200d",x"3a1f0d",x"3b200e",x"3d210e",x"3f230f",x"3d210e",x"3c1f0d",x"361d0c",x"381e0d",x"3a1f0d",x"3c210e",x"3f2310",x"381f0e",x"3e2310",x"3d2310",x"3f2310",x"3f2310",x"3e2310",x"150e07",x"2b180b",x"402410",x"3d220f",x"42372d",x"3d220f",x"3c220f",x"3b200e",x"331c0c",x"3f2411",x"39200e",x"3b210f",x"381f0e",x"150e07",x"42230f",x"150e07",x"150e07",x"000000",x"000000",x"91785b",x"91785b",x"160f07",x"191007",x"191007",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"313131",x"313131",x"333333",x"2f2f2f",x"313131",x"2b2b2b",x"2f2f2f",x"2d2d2d",x"313131",x"2e2e2e",x"2f2f2f",x"323232",x"343434",x"323232",x"2d2d2d",x"242424",x"333333",x"2d2d2d",x"333333",x"2d2d2d",x"303030",x"333333",x"2d2d2d",x"262626",x"2f2f2f",x"312e2c",x"312e2c",x"000000",x"533d2f",x"533d2f",x"150e07",x"442712",x"3b200e",x"311c0c",x"381f0d",x"3b210e",x"402612",x"351d0d",x"3b210f",x"301c0c",x"301c0c",x"311e11",x"311e11",x"3c2514",x"392212",x"3d2412",x"3a2111",x"371f0f",x"341d0e",x"191008",x"39200f",x"48392e",x"492b17",x"442917",x"452a16",x"492d18",x"3e2412",x"331e0e",x"331e0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584e44",x"000000",x"000000",x"000000",x"000000",x"000000",x"573219",x"573219",x"3c2310",x"341e0d",x"311d0d",x"321c0c",x"2f1a0b",x"361e0d",x"3a210f",x"341d0d",x"371f0e",x"371f0e",x"1d1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201408",x"221608",x"1c1208",x"231608",x"231608",x"211508",x"221508",x"291a09",x"271909",x"2d1c0a",x"2c1c09",x"291a09",x"2b1b09",x"301e0a",x"2d1d0a",x"2f1d0a",x"2d1c09",x"281909",x"261809",x"2a1a09",x"231608",x"201408",x"1f1408",x"1a1107",x"1c1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"28170b",x"28170b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584d43",x"584d43",x"473e35",x"42372d",x"513726",x"3c200e",x"3c210f",x"371e0d",x"361d0c",x"3e230f",x"3c210e",x"381e0c",x"3c210e",x"361d0c",x"3e220f",x"472812",x"53493f",x"4a4036",x"473a30",x"483426",x"483426",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"391e0d",x"150e07",x"150e07",x"4d2f1b",x"3b2b1f",x"463d34",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"150e07",x"150e07",x"150e07",x"170f07",x"2f1e13",x"2b1b10",x"24180f",x"24180f",x"000000",x"583f2e",x"583f2e",x"341d0d",x"23150a",x"211409",x"25160a",x"25160a",x"1d1208",x"150e07",x"231409",x"231409",x"25150a",x"2a180b",x"2d1a0b",x"2b190b",x"2b190b",x"25160a",x"26160a",x"27160a",x"221409",x"25150a",x"231509",x"241509",x"221409",x"25150a",x"231409",x"231409",x"27160a",x"241509",x"241509",x"2b180b",x"26160a",x"241509",x"221409",x"231409",x"150e07",x"201208",x"261509",x"1e1208",x"180f07",x"231409",x"241409",x"201309",x"26160a",x"2b190b",x"26160a",x"241509",x"251509",x"251509",x"28170a",x"2a180b",x"25150a",x"1d1108",x"23150a",x"211409",x"1b1008",x"1f1309",x"391e0d",x"150e07",x"876242",x"836041",x"846141",x"815e3f",x"7e5c3f",x"715238",x"7a573a",x"7b583a",x"7c593c",x"7e5c3e",x"775539",x"815f3f",x"856242",x"846244",x"826143",x"75563b",x"7d5b3e",x"805e3f",x"815f40",x"805d40",x"816042",x"846244",x"876545",x"825f42",x"7c5c3f",x"856244",x"825f41",x"7b593b",x"876343",x"856142",x"836041",x"7c5b3e",x"7d5b3d",x"876343",x"825f40",x"7d5b3d",x"825f41",x"7f5c3f",x"7b583b",x"7a573a",x"7d5a3c",x"825f41",x"866041",x"7c5b3d",x"836040",x"876446",x"866445",x"825f41",x"815e40",x"846142",x"876343",x"876343",x"896646",x"886546",x"8c6849",x"513e31",x"513e31",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"472812",x"472812",x"3c2311",x"331d0d",x"361f0e",x"38200e",x"371f0e",x"3d2311",x"301a0b",x"38200e",x"331e0e",x"28180b",x"2f1b0c",x"3f2410",x"39200e",x"1c1108",x"422510",x"2b180b",x"351d0d",x"4e2c14",x"40230e",x"492a13",x"482711",x"492913",x"412511",x"38200e",x"472812",x"2e1a0b",x"341c0c",x"3c200e",x"432510",x"34190a",x"2e1508",x"3f220e",x"40230f",x"422410",x"472711",x"432511",x"432510",x"462711",x"4b2a13",x"472711",x"452712",x"472812",x"4a2b15",x"4b2b14",x"4c2b15",x"4c2c15",x"4e2d16",x"4f2f16",x"4c2b14",x"4d2d15",x"4e2d15",x"4e2d15",x"4b2b15",x"502e16",x"4b2a14",x"4f2d15",x"502f16",x"4e2d15",x"42240f",x"472812",x"482810",x"46260f",x"3e210d",x"472710",x"4a2811",x"502d16",x"492913",x"3d2210",x"29180b",x"482a14",x"221409",x"341d0d",x"2d190b",x"4d2c15",x"1c1108",x"3a210f",x"3b200f",x"381f0e",x"39200e",x"3b210f",x"3b210f",x"3c210f",x"391f0e",x"24150a",x"381e0d",x"2f190b",x"453a31",x"422410",x"38200e",x"3b210e",x"311b0c",x"3e2411",x"371e0d",x"371f0e",x"361e0d",x"150e07",x"482811",x"150e07",x"150e07",x"000000",x"000000",x"887054",x"887054",x"160f07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"303030",x"2f2f2f",x"323232",x"2e2e2e",x"2d2d2d",x"323232",x"2d2d2d",x"2b2b2b",x"333333",x"2e2e2e",x"2c2c2c",x"333333",x"313131",x"2e2e2e",x"1c1c1c",x"202020",x"292929",x"212121",x"333333",x"2d2d2d",x"2f2f2f",x"303030",x"262626",x"2b2b2b",x"2a2a2a",x"282828",x"282828",x"000000",x"503c2f",x"503c2f",x"150e07",x"472912",x"3d2310",x"3f230f",x"3c210f",x"3a200e",x"412712",x"39200e",x"39200e",x"231509",x"231509",x"301d11",x"301d11",x"3b2514",x"362011",x"3e2413",x"3a2111",x"382010",x"2e1b0d",x"190f08",x"3b2210",x"4d3c2f",x"492b17",x"482c17",x"432816",x"492d18",x"382011",x"2b1a0d",x"2b1a0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472812",x"472812",x"331d0d",x"361e0d",x"311c0d",x"311b0c",x"2f1a0b",x"361f0d",x"3b2210",x"3f2511",x"38200f",x"371f0e",x"191008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"1d1308",x"181007",x"1e1308",x"1a1107",x"211508",x"241708",x"271909",x"251809",x"2c1c09",x"271909",x"251708",x"251709",x"271809",x"281909",x"2d1c09",x"2e1d0a",x"2f1d0a",x"321f0a",x"231608",x"2b1b09",x"2d1d0a",x"1f1408",x"191107",x"201508",x"1a1107",x"1b1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"554b40",x"554b40",x"473e35",x"40352c",x"4e3525",x"3b200e",x"3b210f",x"3a200e",x"361d0c",x"3e220f",x"3c210f",x"381f0d",x"341d0c",x"351d0c",x"3c210f",x"472812",x"51473d",x"483e34",x"44362c",x"463223",x"463223",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"160e07",x"150e07",x"150e07",x"2d190b",x"150e07",x"150e07",x"4c3222",x"392c22",x"493f36",x"150e07",x"150e07",x"150e07",x"150e07",x"25160a",x"150e07",x"150e07",x"150e07",x"180f07",x"2e1e12",x"2c1c11",x"1e1710",x"1e1710",x"000000",x"534034",x"534034",x"331d0d",x"23150a",x"26170a",x"201309",x"27170b",x"211309",x"150e07",x"28170a",x"29170a",x"28160a",x"221409",x"26160a",x"29170a",x"27170a",x"241509",x"241509",x"251509",x"26160a",x"29170b",x"221409",x"231409",x"221409",x"221409",x"1f1309",x"25160a",x"231409",x"241509",x"1f1208",x"211309",x"27160a",x"29180a",x"27160a",x"231409",x"241509",x"201309",x"1e1208",x"231409",x"1c1108",x"221409",x"251509",x"221409",x"211309",x"211308",x"211309",x"1e1208",x"211409",x"1f1309",x"251509",x"1e1208",x"211409",x"1d1208",x"201309",x"1d1208",x"211309",x"1d1208",x"381d0c",x"150e07",x"866041",x"846041",x"815f40",x"7a593b",x"775538",x"775638",x"755438",x"7b593c",x"745438",x"775639",x"7a593b",x"846041",x"825f42",x"7d5b3d",x"866443",x"866243",x"825f40",x"856344",x"866445",x"826041",x"7d5b3d",x"7d5b3e",x"7e5b3e",x"815d40",x"815f41",x"846042",x"815f41",x"7d5c3f",x"745439",x"795739",x"7b593c",x"7c5a3c",x"815c3f",x"835f40",x"836041",x"7b593b",x"765538",x"7b593a",x"755438",x"7d5a3d",x"7b593c",x"7b593a",x"7a583b",x"846041",x"7f5d3f",x"7f5c3e",x"866343",x"815e40",x"846041",x"896647",x"886546",x"846243",x"825f40",x"805e40",x"825f41",x"514135",x"514135",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482812",x"482812",x"341e0e",x"38200e",x"3a210f",x"3a200e",x"331c0c",x"311c0d",x"2d180a",x"402512",x"341e0e",x"2b1a0c",x"321c0d",x"4b2c14",x"150e07",x"150e07",x"150e07",x"150e07",x"452811",x"4b2912",x"4b2912",x"462711",x"442611",x"482811",x"3a200e",x"381e0d",x"3b200d",x"3e220f",x"3e220f",x"412511",x"3e2310",x"3a210f",x"402511",x"3f2411",x"3f2411",x"3c220f",x"371f0e",x"3c220f",x"3d230f",x"38200e",x"3a220f",x"39200f",x"382210",x"382210",x"3c2311",x"3a2210",x"351d0d",x"321c0c",x"321c0c",x"3c220f",x"3f2511",x"3d2411",x"402512",x"3f2411",x"3d2310",x"3f2410",x"412511",x"3e230f",x"3e2310",x"412511",x"402410",x"3b210f",x"3f2310",x"412410",x"3c210f",x"3b200e",x"3b210e",x"3c210e",x"391f0d",x"371f0d",x"381e0d",x"391f0d",x"3b200e",x"3a200e",x"1d1108",x"4f2d15",x"2c1a0c",x"3b2210",x"3f2310",x"432612",x"381f0e",x"3d2310",x"3a200e",x"3f2410",x"3f2411",x"26160a",x"3b200d",x"2f190b",x"4a3d32",x"3e210e",x"3c210f",x"381f0e",x"321b0b",x"38200e",x"351d0d",x"381f0e",x"341d0d",x"150e07",x"482913",x"150e07",x"150e07",x"333333",x"323232",x"2f2f2f",x"93795c",x"160f07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d4d4d",x"484848",x"363636",x"303030",x"303030",x"323232",x"323232",x"333333",x"303030",x"2f2f2f",x"303030",x"2e2e2e",x"3f3933",x"605950",x"48433f",x"2d2d2d",x"2f2f2f",x"323232",x"333333",x"303030",x"2a2a2a",x"5b534b",x"5e564e",x"5f574f",x"5f5850",x"5a524a",x"605850",x"5c544c",x"5d544c",x"5e564e",x"585049",x"393736",x"303030",x"303030",x"000000",x"513b2d",x"513b2d",x"150e07",x"4c2c15",x"412511",x"412411",x"432712",x"381f0d",x"422611",x"3b210f",x"3a200e",x"2d190b",x"2d190b",x"2f1d11",x"2f1d11",x"3a2313",x"351f11",x"3e2413",x"3a2111",x"382010",x"2e1a0d",x"180f08",x"402512",x"4c3e33",x"4b2d18",x"452a17",x"422816",x"432916",x"382011",x"331e0f",x"331e0f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2a14",x"4b2a14",x"37200f",x"361f0e",x"361f0e",x"321c0d",x"331c0c",x"3a210f",x"3a210f",x"3b2310",x"3f2310",x"3c220f",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f07",x"191007",x"1a1107",x"150e07",x"1b1108",x"2d1c09",x"291a09",x"2b1b09",x"271809",x"2b1b09",x"261809",x"281909",x"1f1408",x"281909",x"1f1408",x"291a09",x"201508",x"281909",x"2f1d0a",x"281909",x"201408",x"231608",x"291a09",x"201408",x"1b1208",x"201408",x"1e1308",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"52473c",x"52473c",x"433930",x"3c3026",x"4c3120",x"3a1f0d",x"3a200f",x"361e0c",x"361d0c",x"3b210e",x"3e230f",x"371f0d",x"321c0b",x"3a1f0d",x"412410",x"4a2912",x"544a40",x"4b4137",x"47382d",x"4c3526",x"4c3526",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402411",x"402411",x"231509",x"150e07",x"150e07",x"211309",x"150e07",x"150e07",x"543826",x"3b2c22",x"4a4138",x"150e07",x"150e07",x"150e07",x"150e07",x"241509",x"150e07",x"150e07",x"150e07",x"1c1108",x"2f1d12",x"2b1c10",x"251b13",x"251b13",x"000000",x"5d493b",x"5d493b",x"3a2110",x"241409",x"27170b",x"211409",x"211409",x"25160a",x"150e07",x"251509",x"241509",x"27160a",x"27160a",x"28170a",x"241409",x"231509",x"26160a",x"221409",x"25160a",x"221409",x"221409",x"231409",x"27160a",x"26160a",x"26160a",x"25150a",x"26160a",x"241509",x"1e1208",x"221409",x"1e1208",x"201308",x"28170a",x"251509",x"261609",x"29170a",x"27160a",x"26160a",x"25160a",x"26160a",x"27160a",x"211309",x"221409",x"231509",x"211409",x"25160a",x"23150a",x"27160a",x"221409",x"29180b",x"241509",x"1f1309",x"221409",x"201309",x"211409",x"1c1108",x"191008",x"321a0a",x"150e07",x"825f3f",x"826041",x"815f40",x"846040",x"845f40",x"7b593c",x"7f5c3e",x"7d5b3d",x"815f41",x"7d5a3b",x"715034",x"7b5939",x"7f5c3c",x"805e40",x"886546",x"825f41",x"7d5b3d",x"846041",x"896647",x"866345",x"816043",x"876345",x"7a573b",x"7a583b",x"79573a",x"7d5a3e",x"7c5a3b",x"846144",x"7d5b3f",x"866445",x"896547",x"866342",x"7e5c3d",x"886544",x"8a6545",x"825f41",x"7e5c3d",x"805d3e",x"805d3f",x"815d3f",x"836142",x"7d593b",x"6f4f32",x"7c5a3a",x"815d3d",x"7b5a3e",x"846345",x"826041",x"826040",x"846142",x"8c6849",x"836043",x"805e40",x"8c6949",x"7f5b3e",x"53463b",x"53463b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"3d2210",x"3d2210",x"38200f",x"351e0e",x"3c220f",x"3c210f",x"321b0c",x"39200e",x"2d1709",x"24160a",x"361f0f",x"2b190b",x"341e0e",x"482812",x"150e07",x"150e07",x"150e07",x"150e07",x"3e200d",x"3d200d",x"331b0b",x"3a1e0c",x"3a1f0d",x"2f190b",x"432510",x"3d200d",x"3e200d",x"43240f",x"472711",x"41240f",x"3f210e",x"3d200d",x"3e210f",x"442611",x"462711",x"452712",x"432611",x"462712",x"4a2b14",x"4a2b13",x"4d2d16",x"4c2f17",x"492c15",x"452913",x"3e2511",x"3e2410",x"412511",x"452713",x"472913",x"472d15",x"502e16",x"462813",x"502d15",x"4f2d15",x"462914",x"4a2b14",x"4f2e16",x"4a2d15",x"4d2d15",x"472812",x"4a2a13",x"492a14",x"4d2b14",x"4d2c14",x"442711",x"4d2c14",x"4b2a13",x"492912",x"4f2d15",x"4c2b14",x"462711",x"482812",x"462711",x"482811",x"221409",x"4d2b14",x"341f0e",x"4a2c15",x"3a210f",x"432713",x"371e0d",x"412511",x"361d0d",x"3e230f",x"150e07",x"2f1a0c",x"402410",x"2d190b",x"513f33",x"3d1f0d",x"3e2310",x"3f2310",x"311a0b",x"361f0e",x"341c0c",x"3e2411",x"301a0b",x"150e07",x"482913",x"150e07",x"150e07",x"333333",x"333333",x"2e2e2e",x"4f4f4f",x"160f07",x"180f07",x"180f07",x"484848",x"4b4b4b",x"4e4e4e",x"4d4d4d",x"333333",x"515151",x"484848",x"303030",x"303030",x"303030",x"323232",x"323232",x"303030",x"303030",x"2f2f2f",x"2e2e2e",x"393938",x"605a55",x"5b534a",x"514d48",x"5a5a5a",x"323232",x"323232",x"323232",x"323232",x"303030",x"585047",x"605951",x"676059",x"665f59",x"655e57",x"635b54",x"615951",x"5d564e",x"615950",x"5e564f",x"383736",x"313131",x"313131",x"000000",x"533d2e",x"533d2e",x"150e07",x"432611",x"412511",x"432611",x"3f2410",x"3d2310",x"422611",x"3c220f",x"371e0d",x"251509",x"251509",x"2f1d11",x"2f1d11",x"382213",x"382112",x"412614",x"3d2412",x"372010",x"29180c",x"180f08",x"3b2210",x"4b3c30",x"52321c",x"472a17",x"432816",x"442917",x"382010",x"2c1a0d",x"2c1a0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482812",x"482812",x"402612",x"3a220f",x"3b2210",x"3a200e",x"381f0e",x"341d0d",x"361f0e",x"3e2411",x"3c230f",x"3f230f",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"231608",x"301e0a",x"2b1b09",x"251709",x"291a09",x"261809",x"2e1d0a",x"2d1c09",x"1f1408",x"231608",x"221508",x"1b1108",x"221608",x"221608",x"2a1b09",x"2d1c09",x"261809",x"281909",x"291a09",x"1c1208",x"1a1107",x"201408",x"231608",x"1b1108",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"53483e",x"53483e",x"433a31",x"3c2e24",x"482d1c",x"371d0d",x"39200e",x"381f0d",x"381e0d",x"3c210e",x"3b200e",x"3b200e",x"3a1f0d",x"3a200e",x"402310",x"4a2912",x"554b41",x"4d4137",x"45362b",x"4e3524",x"4e3524",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b180a",x"2b180a",x"2e1a0b",x"150e07",x"150e07",x"2f1b0b",x"150e07",x"150e07",x"533725",x"3c2d22",x"4a4138",x"150e07",x"150e07",x"150e07",x"150e07",x"251509",x"150e07",x"150e07",x"150e07",x"1d1108",x"322114",x"312013",x"271c14",x"271c14",x"000000",x"5c4a3c",x"5c4a3c",x"392110",x"29180b",x"27170a",x"2a180b",x"2b190c",x"1c1108",x"150e07",x"251509",x"231409",x"251509",x"251509",x"27160a",x"241509",x"25150a",x"251509",x"231409",x"29180b",x"28170a",x"25150a",x"251509",x"25150a",x"27160a",x"25160a",x"25150a",x"241509",x"26160a",x"28170a",x"241509",x"231509",x"211409",x"221409",x"27160a",x"27170a",x"2b190b",x"2b190b",x"27170a",x"2b190c",x"26160a",x"26160a",x"1b1108",x"201309",x"1c1108",x"251509",x"221409",x"231509",x"231409",x"251509",x"211309",x"1f1208",x"201309",x"170f07",x"150e07",x"170f07",x"1f1208",x"1e1108",x"331a0b",x"150e07",x"7d5b3d",x"815c3e",x"7c5b3c",x"7d5a3d",x"7e5c3f",x"705036",x"7a583b",x"77553a",x"7a593b",x"7f5b3a",x"775738",x"775737",x"755436",x"7b593c",x"7b5a3d",x"745337",x"6f4e34",x"745438",x"765539",x"7d5c3d",x"7d5b3d",x"7c5b3e",x"78563a",x"7d5a3c",x"7b593c",x"705035",x"735337",x"765639",x"7d5b3d",x"77563a",x"755538",x"7d5a3d",x"79583b",x"7d5a3c",x"7d5b3d",x"7a583b",x"7b5a3d",x"785639",x"7e5b3e",x"76553a",x"7a593b",x"7e5a3a",x"7a5838",x"775536",x"795738",x"7a593c",x"7c5a3b",x"7b593b",x"755237",x"78573a",x"77563a",x"815e3f",x"815d3f",x"896545",x"805d3e",x"59493c",x"59493c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"311d0d",x"341e0e",x"2f1b0c",x"3c2511",x"38200e",x"3a210f",x"150e07",x"331f0f",x"371f0e",x"2a180a",x"301a0b",x"462710",x"150e07",x"150e07",x"150e07",x"150e07",x"482812",x"482711",x"3d210e",x"40230f",x"43230f",x"3b200e",x"492913",x"492912",x"472812",x"452611",x"442510",x"442611",x"452611",x"432410",x"452711",x"472812",x"462711",x"452712",x"432511",x"432511",x"412411",x"442711",x"462812",x"432611",x"432612",x"3f2410",x"3f2410",x"3e220f",x"402410",x"412410",x"3f2410",x"422711",x"422510",x"402310",x"422510",x"422511",x"432612",x"472913",x"462812",x"432712",x"452812",x"3f2410",x"422511",x"462813",x"472913",x"442712",x"462913",x"472913",x"452711",x"412410",x"402410",x"3f220f",x"3d220e",x"3d210f",x"452611",x"482811",x"512e15",x"553117",x"351f0f",x"4b2c16",x"3b210f",x"3f2512",x"39200d",x"3f2411",x"402511",x"150e07",x"341e0e",x"341d0d",x"472913",x"361e0d",x"4a3f35",x"3f200e",x"3e2410",x"3c210f",x"361e0d",x"2b190b",x"2f1b0c",x"3a210f",x"351d0d",x"150e07",x"492913",x"150e07",x"150e07",x"323232",x"323232",x"323232",x"3b3b3b",x"313131",x"363636",x"464646",x"484848",x"4b4b4b",x"4e4e4e",x"4d4d4d",x"333333",x"333333",x"303030",x"323232",x"323232",x"313131",x"323030",x"323030",x"323232",x"303030",x"2f2f2f",x"2e2e2e",x"393938",x"665f59",x"5a524b",x"4e4842",x"616161",x"333333",x"333333",x"313131",x"323232",x"303030",x"5b534c",x"635c54",x"615952",x"605850",x"5d554d",x"615951",x"5f574f",x"5b524a",x"5a524a",x"5a534b",x"333333",x"333333",x"333333",x"000000",x"523c2e",x"523c2e",x"150e07",x"462813",x"3e2310",x"3f2411",x"39200e",x"2b190b",x"3a2110",x"361e0e",x"341c0c",x"1d1108",x"1d1108",x"2f1d10",x"2f1d10",x"382112",x"382112",x"3f2613",x"3e2513",x"382010",x"301a0d",x"190f08",x"3f2410",x"4e3f33",x"50311a",x"452a17",x"3c2212",x"402614",x"3b2211",x"301d0e",x"301d0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"353535",x"323232",x"333333",x"323232",x"333333",x"000000",x"4a4a4a",x"4e4e4e",x"404040",x"474646",x"3c3c3c",x"000000",x"000000",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"494440",x"494440",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"47433e",x"48443f",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"63605d",x"64615e",x"000000",x"000000",x"472812",x"472812",x"341f0e",x"3b2210",x"3d2311",x"371f0e",x"3a210f",x"2d190b",x"361f0f",x"341e0e",x"361f0e",x"3a200e",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1108",x"2b1b09",x"2c1c09",x"1e1308",x"181007",x"281909",x"2d1d0a",x"34200a",x"291a09",x"211508",x"241708",x"241708",x"201508",x"211508",x"2a1a09",x"2d1d0a",x"2c1c09",x"281a09",x"301e0a",x"2c1c09",x"261809",x"181007",x"231608",x"261809",x"1a1107",x"150e07",x"160e07",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594e43",x"594e43",x"433a31",x"3d3229",x"513622",x"381d0d",x"371f0e",x"351d0c",x"381e0d",x"40240f",x"432611",x"3a1f0d",x"391f0d",x"3d220f",x"412410",x"4c2a13",x"51473d",x"4a4036",x"48392e",x"4f3626",x"4f3626",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"29170a",x"150e07",x"150e07",x"2b180b",x"150e07",x"150e07",x"563826",x"3c2e23",x"494036",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"150e07",x"382418",x"2f1e12",x"2b1f15",x"2b1f15",x"000000",x"5e4a3d",x"5e4a3d",x"37210f",x"25160a",x"221409",x"24150a",x"2a190b",x"1d1108",x"150e07",x"27160a",x"29170b",x"25150a",x"241509",x"27160a",x"27160a",x"231409",x"241509",x"231409",x"231409",x"26160a",x"29170b",x"241509",x"25150a",x"231509",x"27160a",x"211409",x"27170a",x"24150a",x"241509",x"24150a",x"2a180b",x"25160a",x"29180b",x"231409",x"231409",x"25150a",x"24150a",x"251509",x"28170a",x"241409",x"241509",x"27170a",x"28170a",x"170f07",x"231409",x"1e1208",x"1f1209",x"2b180b",x"231409",x"27160a",x"26160a",x"1f1208",x"201309",x"23150a",x"241509",x"201309",x"1f1208",x"331a0b",x"150e07",x"77563a",x"7a583b",x"7a583b",x"705036",x"76563a",x"6e4e34",x"533723",x"6d4d34",x"735437",x"715233",x"7b5838",x"7d5a3b",x"755438",x"755437",x"745337",x"7b593c",x"816041",x"7e5b3d",x"805e40",x"7d5b3e",x"7b583b",x"7f5c3d",x"765538",x"745337",x"77563a",x"725336",x"78573a",x"7f5b3e",x"7c5a3c",x"765539",x"76563a",x"78573b",x"78563a",x"7a593b",x"7b593c",x"735237",x"765639",x"715035",x"5d3e26",x"705035",x"78563a",x"6f5033",x"855e3d",x"7c583a",x"7b5a3b",x"79583a",x"7f5b3c",x"825f3f",x"856243",x"815e3f",x"826041",x"856142",x"825d3f",x"845f40",x"805d3f",x"544539",x"544539",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"412510",x"412510",x"351f0e",x"311c0c",x"361f0e",x"362210",x"3b210f",x"150e07",x"1d1007",x"35200f",x"341d0d",x"251509",x"311b0b",x"472710",x"150e07",x"150e07",x"150e07",x"150e07",x"361d0b",x"2c1407",x"2c1407",x"3b1f0c",x"381c0b",x"4a2b14",x"2e2e2e",x"492912",x"472812",x"452611",x"442510",x"442611",x"452611",x"2e2e2e",x"2b2b2b",x"323232",x"323232",x"452712",x"432511",x"323232",x"323232",x"363636",x"444444",x"5d5d5c",x"4f4f4f",x"3f2410",x"484847",x"4c4c4c",x"4a4a4a",x"383838",x"3a3a3a",x"313131",x"313131",x"313131",x"322c28",x"575757",x"636363",x"535353",x"515151",x"585858",x"4a4a4a",x"454545",x"5d5d5d",x"555555",x"5d5c5c",x"323232",x"333333",x"303131",x"452711",x"412410",x"402410",x"3f220f",x"3d220e",x"3d210f",x"452611",x"512e16",x"512e16",x"512e15",x"341e0e",x"452813",x"3b200e",x"3f2511",x"241509",x"412511",x"3d2310",x"26170b",x"331e0e",x"331c0c",x"4d2c15",x"371e0d",x"4b3f35",x"3c1f0d",x"3f2411",x"3c220f",x"3a200e",x"422611",x"150e07",x"331d0d",x"321c0c",x"150e07",x"4d2c15",x"150e07",x"150e07",x"323232",x"333333",x"303030",x"333333",x"333333",x"4d4d4d",x"353535",x"313131",x"303030",x"313131",x"323232",x"363636",x"313131",x"333333",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"303030",x"323232",x"2f2f2f",x"333333",x"4e4943",x"5d554d",x"494440",x"525252",x"2a2a2a",x"262626",x"2e2e2e",x"2f2f2f",x"242424",x"585048",x"5d554d",x"5e574f",x"5b534c",x"5e554d",x"5f574e",x"5c544c",x"5e564e",x"5f564e",x"5b534c",x"373634",x"292929",x"292929",x"000000",x"513b2c",x"513b2c",x"150e07",x"4a2b15",x"3d220f",x"361f0e",x"3b210f",x"3b2210",x"150e07",x"38200e",x"3b210e",x"2b180b",x"2b180b",x"2f1d10",x"2f1d10",x"382213",x"351f11",x"3d2513",x"3a2111",x"392010",x"301b0c",x"191008",x"3c220f",x"503f34",x"4f2f19",x"492b17",x"422714",x"422615",x"341f10",x"2c1a0c",x"2c1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"353535",x"353535",x"323232",x"333333",x"323232",x"333333",x"363636",x"4d4d4d",x"4e4e4e",x"404040",x"474646",x"3c3c3c",x"3d3d3d",x"2c2c2c",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"4d4945",x"494440",x"494440",x"353535",x"353535",x"000000",x"000000",x"000000",x"484440",x"47423e",x"48443f",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"615e5b",x"63605d",x"64615e",x"6b6866",x"000000",x"4a2b14",x"4a2b14",x"321d0d",x"37200f",x"3a2110",x"371f0e",x"3c2310",x"331d0d",x"3a210f",x"351e0e",x"3a210f",x"3c210f",x"1d1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"201408",x"241708",x"261809",x"1d1308",x"201408",x"301e0a",x"2d1d0a",x"271909",x"2a1a09",x"281909",x"261809",x"2a1a09",x"241708",x"241708",x"2c1c09",x"2e1d0a",x"2b1b09",x"241708",x"251809",x"2a1b09",x"271909",x"1c1208",x"1e1308",x"241708",x"1b1108",x"150e07",x"170f07",x"180f07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"544a40",x"544a40",x"463d34",x"3d3127",x"523521",x"432611",x"3a200e",x"361d0d",x"391f0d",x"40240f",x"402410",x"3a1f0d",x"331c0b",x"442611",x"412510",x"492812",x"554b41",x"443a31",x"43352b",x"4e3424",x"4e3424",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"251509",x"4b2c15",x"150e07",x"26160a",x"150e07",x"150e07",x"4e3526",x"3c2d23",x"4d433a",x"150e07",x"150e07",x"150e07",x"150e07",x"25150a",x"150e07",x"150e07",x"150e07",x"150e07",x"362519",x"312115",x"291f17",x"291f17",x"000000",x"5d4c3f",x"5d4c3f",x"392110",x"301c0d",x"25160a",x"221409",x"2b190c",x"201309",x"150e07",x"241509",x"231409",x"251509",x"221309",x"27160a",x"241509",x"29170a",x"241509",x"211308",x"1f1208",x"1f1208",x"241509",x"241509",x"25150a",x"231509",x"29180b",x"211409",x"28170a",x"28160a",x"1d1108",x"241509",x"26160a",x"241509",x"241409",x"231509",x"231409",x"201309",x"24150a",x"221409",x"29170a",x"261609",x"251509",x"241409",x"231409",x"211308",x"1e1108",x"1c1108",x"211309",x"231409",x"211309",x"241509",x"231409",x"201308",x"1f1208",x"211409",x"211409",x"201309",x"1d1108",x"351b0b",x"150e07",x"846041",x"7a583b",x"7b583b",x"7a593b",x"7a583b",x"79583a",x"735336",x"705034",x"6f4e33",x"79583b",x"7f5e3f",x"7d5b3e",x"7d5b3c",x"7a583b",x"825f41",x"886546",x"846345",x"815d3e",x"805d3d",x"7c5a3c",x"805c3e",x"7d5b3d",x"7f5c3d",x"7a583b",x"78573b",x"7c5a3d",x"77563a",x"7e5b3e",x"735238",x"7a593b",x"76553a",x"7a583c",x"7c5a3c",x"755539",x"7b593c",x"7c5a3c",x"78563a",x"7e5c3d",x"785638",x"725035",x"725035",x"815f3f",x"886544",x"856142",x"815c3e",x"866141",x"876443",x"8a6647",x"896647",x"7e5b3d",x"846040",x"825e40",x"805c3e",x"815e3f",x"866142",x"55473c",x"55473c",x"28170a",x"311b0b",x"000000",x"000000",x"40240f",x"4e2c14",x"5b4e43",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"422511",x"422511",x"3c2310",x"351e0e",x"25150a",x"1f1309",x"392411",x"150e07",x"27160a",x"2a180b",x"2d1a0b",x"241509",x"2c180a",x"43250f",x"371f0d",x"24150a",x"1e1309",x"1e1209",x"4a2a13",x"331d0d",x"432611",x"472711",x"341d0d",x"323232",x"424242",x"5c5c5c",x"363636",x"363636",x"323232",x"3b3b3b",x"686867",x"474747",x"2b2b2b",x"323232",x"343434",x"626262",x"626262",x"333333",x"323232",x"393939",x"5f5f5e",x"494949",x"4f4f4f",x"373737",x"353535",x"4c4c4c",x"565554",x"3f3f3f",x"313131",x"313131",x"313131",x"313131",x"393939",x"575757",x"636363",x"535353",x"515151",x"585858",x"4a4a4a",x"454545",x"5d5d5d",x"555555",x"393939",x"323232",x"333333",x"303131",x"303131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"522f15",x"522f15",x"502e15",x"2d1a0c",x"4b2c16",x"3c220f",x"321d0d",x"221409",x"3d2310",x"150e07",x"2a180b",x"29180b",x"2e1a0b",x"452813",x"3b210f",x"4b4035",x"3f220e",x"3a2210",x"39200f",x"3d2310",x"381f0d",x"150e07",x"311c0c",x"361e0d",x"150e07",x"492812",x"150e07",x"150e07",x"323232",x"333333",x"323232",x"313131",x"333333",x"323232",x"323232",x"333333",x"313131",x"333333",x"3c3c3c",x"343433",x"323232",x"333333",x"313131",x"333333",x"38210e",x"180f07",x"323232",x"333333",x"323232",x"454545",x"3e3e3d",x"3f3e3e",x"6e6964",x"5e564e",x"605c59",x"5f5f5f",x"313131",x"323232",x"323232",x"343434",x"323232",x"5e564f",x"6c6660",x"6e6761",x"6e6861",x"6c655e",x"6b655e",x"67615a",x"655e57",x"5e564e",x"59514a",x"353534",x"2e2e2e",x"2e2e2e",x"000000",x"543d2d",x"543d2d",x"150e07",x"442712",x"3d220f",x"39200e",x"3b2210",x"402511",x"150e07",x"331d0d",x"331c0d",x"28170a",x"28170a",x"2e1c10",x"2e1c10",x"362113",x"351f10",x"3c2313",x"382010",x"331d0e",x"2d190b",x"180f08",x"3f2411",x"533f32",x"52321a",x"472b17",x"472b17",x"452a17",x"3d2212",x"2b1a0c",x"2b1a0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"303030",x"343434",x"333333",x"323232",x"333232",x"383838",x"323232",x"333333",x"303030",x"424242",x"434343",x"3b3b3b",x"2c2c2c",x"343434",x"323232",x"333232",x"000000",x"45413e",x"474340",x"4d4945",x"494440",x"313232",x"313131",x"2f2f2f",x"000000",x"3f3c39",x"433f3b",x"484440",x"46423e",x"313131",x"313131",x"333333",x"000000",x"000000",x"44403d",x"504c49",x"605d5a",x"6b6866",x"6a6765",x"6a6765",x"462812",x"462812",x"3c2310",x"402511",x"3c2310",x"341d0d",x"38200f",x"36200e",x"361f0e",x"38200e",x"3b210f",x"39200e",x"1d1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"261809",x"271809",x"221508",x"261809",x"2b1b09",x"321f0a",x"2f1e0a",x"251809",x"2e1d0a",x"2c1c09",x"271909",x"291a09",x"201508",x"2a1a09",x"2a1a09",x"33200a",x"291a09",x"201408",x"211508",x"2a1b09",x"221508",x"1f1408",x"281a09",x"241708",x"1c1208",x"150e07",x"170f07",x"180f07",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574d43",x"574d43",x"4c4239",x"40352c",x"4e3322",x"442711",x"371f0e",x"381f0d",x"381f0d",x"3e230f",x"3e220f",x"361e0c",x"361c0b",x"402410",x"432611",x"482811",x"564c42",x"463b32",x"3f3126",x"4d3221",x"4d3221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"27170b",x"4c2b14",x"201309",x"191008",x"3f230f",x"150e07",x"573a28",x"3a2b20",x"4e443b",x"150e07",x"150e07",x"150e07",x"150e07",x"2b190c",x"150e07",x"150e07",x"150e07",x"1a1008",x"32231a",x"312116",x"2f251c",x"2f251c",x"000000",x"624f41",x"624f41",x"3a2210",x"26160a",x"211409",x"231409",x"27170a",x"1e1208",x"150e07",x"29180a",x"27160a",x"27160a",x"221409",x"29170a",x"29170a",x"29170a",x"27160a",x"211309",x"261509",x"201309",x"241509",x"26160a",x"251509",x"201309",x"231409",x"26160a",x"26160a",x"25160a",x"25160a",x"25150a",x"27170a",x"201309",x"28170a",x"26160a",x"261609",x"221409",x"1d1208",x"211309",x"231509",x"25160a",x"231509",x"1d1108",x"221409",x"241509",x"25160a",x"26160a",x"2b190b",x"201309",x"231409",x"241509",x"201309",x"241409",x"1e1208",x"201309",x"241509",x"201208",x"1f1309",x"361c0b",x"160f07",x"825e40",x"805c3e",x"7d5a3d",x"7e5b3e",x"7b583c",x"76563a",x"7c5a3b",x"7d5c3e",x"816040",x"77563a",x"7d5b3c",x"805c3e",x"7b593b",x"715034",x"765539",x"7d5c3e",x"7b593b",x"745437",x"64452c",x"77563a",x"7c5a3c",x"836041",x"7f5d3f",x"846244",x"7e5e41",x"815e40",x"815f41",x"816041",x"846242",x"815e40",x"805e40",x"805d3f",x"7a583b",x"7c593c",x"7f5b3e",x"7d5b3e",x"7b583b",x"7c5a3c",x"7e5b3c",x"826041",x"816040",x"7c593c",x"815e3e",x"805e3e",x"805d3d",x"795739",x"7d5a3c",x"836041",x"7e5b3d",x"7a593a",x"69462d",x"7f5c3e",x"815d40",x"846142",x"856243",x"56473b",x"1e1108",x"28170a",x"311b0b",x"170f07",x"40240f",x"40240f",x"4e2c14",x"5b4e43",x"5b4e43",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"38200f",x"2e1b0d",x"150e07",x"1c1108",x"372210",x"150e07",x"1c1108",x"150e07",x"2c190b",x"221409",x"2a170a",x"3e220e",x"323232",x"323232",x"393939",x"150e07",x"1d1108",x"2c1a0b",x"381f0e",x"381f0d",x"312e2c",x"313131",x"313131",x"5c5c5c",x"363636",x"313131",x"323232",x"3b3b3b",x"3b3b3b",x"565656",x"313131",x"343434",x"333333",x"616161",x"626262",x"333333",x"323232",x"3e3e3e",x"434242",x"494848",x"484848",x"323232",x"323232",x"323232",x"343434",x"323232",x"333333",x"313131",x"323232",x"303030",x"2f2f2f",x"323232",x"5a5a5a",x"363636",x"323232",x"323232",x"313131",x"333333",x"323232",x"323232",x"333333",x"333333",x"313131",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583419",x"583419",x"553319",x"382110",x"4b2d16",x"331c0c",x"442813",x"190f08",x"3f2411",x"3c210f",x"1a1008",x"150e07",x"2e1a0c",x"432511",x"3a200e",x"4e4238",x"3e210f",x"3c2310",x"38200e",x"3f2310",x"412511",x"442813",x"2f1c0c",x"3a210f",x"150e07",x"452610",x"150e07",x"150e07",x"000000",x"323232",x"333333",x"333333",x"323232",x"323232",x"323232",x"333333",x"323232",x"333333",x"3c3c3c",x"343433",x"323232",x"000000",x"452812",x"452812",x"38210e",x"180f07",x"150e07",x"323232",x"313131",x"313131",x"434343",x"585857",x"75706a",x"69645e",x"6a6561",x"5e5e5d",x"333333",x"333333",x"373737",x"4b4b4b",x"525252",x"6c655f",x"6b645e",x"6d6660",x"6d6760",x"6d6660",x"6c665f",x"645d56",x"68615a",x"655e56",x"5f5952",x"333333",x"323232",x"323232",x"000000",x"533d2d",x"533d2d",x"150e07",x"3d220f",x"371f0e",x"371f0d",x"3f2311",x"402512",x"3c230f",x"29180b",x"311c0c",x"25150a",x"25150a",x"2d1c0f",x"2d1c0f",x"352011",x"351f10",x"3a2111",x"392111",x"301b0d",x"29170b",x"180f07",x"3f2411",x"534134",x"4d2d18",x"432715",x"472c17",x"482b17",x"3e2513",x"382110",x"382110",x"373737",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"313131",x"313131",x"333333",x"333333",x"323232",x"313131",x"323232",x"333333",x"323232",x"363636",x"323232",x"313131",x"333333",x"303030",x"313131",x"383838",x"303030",x"2f2f2f",x"333232",x"313131",x"3c352f",x"3f3d3b",x"45413d",x"696664",x"414141",x"343434",x"2d2d2d",x"313131",x"383737",x"3a3937",x"433f3c",x"46423e",x"444241",x"323232",x"353535",x"333333",x"313131",x"3a3937",x"3e3b39",x"44403d",x"656260",x"424242",x"3e3e3e",x"000000",x"452812",x"452812",x"3d2310",x"3b220f",x"3d2411",x"381f0e",x"3a220f",x"3d2411",x"351f0e",x"3c220f",x"3e2310",x"3a210e",x"1e1208",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191007",x"251708",x"271809",x"271909",x"201508",x"2e1d0a",x"2f1d0a",x"281909",x"261809",x"2d1d0a",x"2b1b09",x"2d1c09",x"291a09",x"211508",x"301e0a",x"231608",x"211508",x"261809",x"2a1a09",x"271809",x"2d1c09",x"291a09",x"1e1308",x"1d1308",x"1c1208",x"191007",x"150e07",x"160e07",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"51483e",x"51483e",x"473e35",x"43372d",x"4f3525",x"442611",x"341c0c",x"3b200e",x"391f0d",x"412511",x"402410",x"422410",x"381d0c",x"3a1f0d",x"422511",x"462610",x"554b41",x"483c32",x"403228",x"493021",x"493021",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1108",x"1d1108",x"231409",x"482913",x"2a190b",x"150e07",x"492912",x"2c190b",x"543827",x"3d2c20",x"4b4239",x"150e07",x"150e07",x"150e07",x"150e07",x"29190b",x"150e07",x"150e07",x"150e07",x"1a1008",x"33251b",x"342419",x"342a21",x"342a21",x"000000",x"5b483a",x"5b483a",x"28160a",x"1e1208",x"241509",x"27160a",x"29170a",x"241509",x"241509",x"251509",x"221309",x"1f1108",x"201208",x"211308",x"231409",x"261609",x"251509",x"251509",x"281609",x"221309",x"201208",x"211309",x"221309",x"1d1108",x"1d1108",x"211308",x"251509",x"281609",x"281609",x"261509",x"231409",x"201309",x"201208",x"1f1208",x"1e1208",x"211409",x"28170a",x"201309",x"27160a",x"201309",x"1f1309",x"251509",x"211309",x"1f1208",x"221308",x"1f1208",x"201308",x"231409",x"231409",x"1f1309",x"1f1208",x"28170a",x"221409",x"28170a",x"261609",x"251509",x"261509",x"462610",x"181007",x"795739",x"775539",x"775639",x"735135",x"795739",x"7e5c3d",x"7e5b3e",x"7d5a3e",x"7c593b",x"705033",x"79573a",x"7c5a3d",x"765538",x"745336",x"795639",x"7a593b",x"7e5c3f",x"815f41",x"7f5e41",x"7b593b",x"79573a",x"7e5c3f",x"7c5c3e",x"7f5b3e",x"79583b",x"7b593b",x"775639",x"7b593b",x"7c5a3d",x"745438",x"765438",x"735236",x"765539",x"755438",x"7a583a",x"745236",x"795739",x"7e5c3d",x"7c5a3d",x"7b5a3d",x"7a583b",x"745335",x"7e5c3c",x"835f41",x"835f3f",x"7d5a3b",x"7e5a3c",x"815e3f",x"845f42",x"8d6948",x"886546",x"805d3e",x"805c3e",x"815e3f",x"856142",x"56483d",x"150e07",x"150e07",x"150e07",x"160e07",x"422611",x"422611",x"473e35",x"584c42",x"584c42",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"412410",x"412410",x"361f0f",x"361f0e",x"3d2511",x"321f0e",x"34200f",x"3c2512",x"2f1b0c",x"371f0e",x"231409",x"231409",x"28170a",x"41240f",x"313131",x"323232",x"323232",x"3c3c3c",x"4f4f4f",x"535353",x"5a5a5a",x"414141",x"323232",x"323232",x"333333",x"414141",x"333333",x"312f2d",x"333333",x"333333",x"3a3a3a",x"656462",x"3e3e3e",x"323232",x"5c5c5c",x"313131",x"5e5e5e",x"323232",x"333333",x"515151",x"646360",x"606060",x"454545",x"303030",x"333333",x"323232",x"585655",x"3c3c3c",x"333333",x"333333",x"323231",x"313131",x"323232",x"3f3f3f",x"5a5a59",x"5b5b5b",x"333333",x"323232",x"363636",x"333333",x"333333",x"333333",x"333333",x"32302f",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583419",x"583419",x"583419",x"311c0d",x"4d2e16",x"3e230f",x"472a14",x"2e1a0b",x"3a2110",x"371f0e",x"2d1a0c",x"3b2210",x"26160a",x"3b200e",x"381f0e",x"4f4339",x"40230f",x"3b220f",x"3c220f",x"3e2411",x"402511",x"402512",x"301b0c",x"3b210e",x"150e07",x"43240f",x"150e07",x"150e07",x"000000",x"474747",x"313131",x"353535",x"343434",x"343434",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"412610",x"412610",x"2a190b",x"170f07",x"150e07",x"150e07",x"150e07",x"2a180a",x"515151",x"626262",x"676665",x"61605e",x"676767",x"636262",x"393939",x"323232",x"515151",x"5b5b5b",x"595959",x"5e5d5d",x"636261",x"636261",x"656462",x"666564",x"61605f",x"605e5d",x"5c5a59",x"595856",x"575655",x"383838",x"313131",x"313131",x"000000",x"50392a",x"50392a",x"150e07",x"472812",x"351e0d",x"3a210f",x"3c210f",x"3e2310",x"402511",x"301c0c",x"381f0e",x"301c0d",x"301c0d",x"2b1b10",x"2b1b10",x"321e11",x"341f10",x"3a2212",x"382010",x"331d0e",x"29170a",x"180f07",x"3c2210",x"5e4738",x"492c17",x"4a2c18",x"402614",x"442815",x"402514",x"2b1a0c",x"333333",x"373737",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"3c3c3c",x"313131",x"323232",x"323232",x"323232",x"3b3937",x"383736",x"363635",x"373635",x"313131",x"333333",x"464646",x"323232",x"323232",x"313131",x"303030",x"323232",x"343434",x"343434",x"444444",x"5e5e5e",x"434242",x"3a3837",x"656362",x"373737",x"3e3e3e",x"333333",x"444444",x"414242",x"4d4d4d",x"3b3937",x"61605f",x"6b6866",x"323232",x"313131",x"474747",x"323232",x"484848",x"363534",x"3b3a38",x"666562",x"3e3e3e",x"3c3c3c",x"424242",x"000000",x"462913",x"462913",x"37200f",x"3c2310",x"3c2310",x"38200e",x"38200e",x"39210f",x"39210f",x"38200e",x"3a210f",x"3d2310",x"190f08",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1308",x"271909",x"241708",x"1f1408",x"1f1408",x"2b1b09",x"241708",x"241708",x"231608",x"291a09",x"291a09",x"2d1c0a",x"2f1e0a",x"241708",x"2f1e0a",x"2a1a09",x"241708",x"201408",x"2c1c09",x"2a1b09",x"271909",x"251809",x"1b1108",x"150e07",x"160e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"51473e",x"51473e",x"3f362d",x"33261d",x"4a2d1c",x"412511",x"39200e",x"3f2310",x"361d0d",x"432712",x"442611",x"402310",x"3a1f0c",x"361c0c",x"432711",x"462611",x"52483e",x"493d34",x"413429",x"493223",x"493223",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"241509",x"241509",x"150e07",x"150e07",x"2a190b",x"150e07",x"4d2d15",x"150e07",x"503727",x"3c2c20",x"4b4036",x"150e07",x"150e07",x"150e07",x"150e07",x"291a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"36271d",x"35261c",x"392e26",x"392e26",x"000000",x"584639",x"584639",x"361f0e",x"2f1b0c",x"2c1a0b",x"29180b",x"2b190b",x"2a180b",x"29170a",x"24150a",x"28170a",x"2a190b",x"29180b",x"2c1a0c",x"2d1a0c",x"27160a",x"24150a",x"28170a",x"25150a",x"251509",x"2a180a",x"251509",x"231509",x"231409",x"1f1208",x"221309",x"211309",x"271509",x"261509",x"26160a",x"26160a",x"221409",x"180f07",x"26160a",x"1e1209",x"28180b",x"28170b",x"2b190b",x"25160a",x"241509",x"26160a",x"231409",x"231409",x"231409",x"231409",x"1f1208",x"1d1208",x"251509",x"211409",x"27160a",x"24150a",x"150e07",x"24150a",x"221409",x"24150a",x"27170a",x"241509",x"4a2a13",x"170f07",x"845f40",x"835e3f",x"7c5a3d",x"755539",x"7e5c3e",x"7f5e3f",x"805e40",x"7b593c",x"7c5a3d",x"7d5b3c",x"78573a",x"7c5b3d",x"765639",x"755538",x"765438",x"715136",x"755437",x"77563a",x"7e5c3e",x"7a593b",x"79583c",x"6d4d33",x"5a3a20",x"765639",x"775538",x"765638",x"79573a",x"725236",x"7d5a3d",x"7b5a3c",x"7f5d3f",x"7c5b3c",x"765539",x"79573a",x"77563a",x"755539",x"7b5a3d",x"815f41",x"896544",x"7e5b3d",x"805e3f",x"7c5a3b",x"79583a",x"836041",x"815e3e",x"7e5b3d",x"7b593c",x"7a593b",x"7b593a",x"815d3f",x"836041",x"7f5b3e",x"7d5b3e",x"725136",x"613f25",x"57473c",x"150e07",x"150e07",x"150e07",x"150e07",x"452916",x"452916",x"423328",x"4a2a13",x"4a2a13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452611",x"452611",x"39200f",x"3f2511",x"3d2311",x"3f2713",x"3e2411",x"33200f",x"351d0d",x"351d0d",x"241509",x"28170a",x"361f0e",x"40230e",x"333333",x"323232",x"333333",x"353535",x"313131",x"313131",x"464646",x"5b5b5b",x"606060",x"5d5d5c",x"626262",x"434242",x"333333",x"323232",x"323232",x"333333",x"494949",x"5e5e5e",x"505050",x"313131",x"323232",x"333333",x"313131",x"323231",x"323232",x"646463",x"636261",x"606060",x"5f5f5f",x"464646",x"656464",x"5c5c5c",x"323232",x"5c5c5c",x"595959",x"5b5b5b",x"525251",x"474747",x"565656",x"5f5f5f",x"595959",x"545454",x"403e3e",x"323232",x"363636",x"333333",x"333333",x"333333",x"333333",x"32302f",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"573318",x"573318",x"593419",x"351e0e",x"4b2d16",x"3f2310",x"462813",x"3c210e",x"412511",x"402511",x"3a210f",x"341e0d",x"1d1108",x"3e220f",x"341c0c",x"56493e",x"40230f",x"3b2210",x"361e0d",x"22140a",x"3f2512",x"150e07",x"321c0d",x"381f0e",x"150e07",x"4d2a14",x"150e07",x"150e07",x"636261",x"636261",x"545454",x"595959",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"37200d",x"37200d",x"170f07",x"160e07",x"150e07",x"150e07",x"150e07",x"221409",x"221409",x"626262",x"676665",x"61605e",x"676767",x"636262",x"393939",x"323232",x"515151",x"5b5b5b",x"595959",x"5e5d5d",x"636261",x"636261",x"656462",x"666564",x"61605f",x"605e5d",x"5c5a59",x"595856",x"575655",x"383838",x"000000",x"000000",x"000000",x"4f3627",x"4f3627",x"150e07",x"452712",x"3b200e",x"3a2110",x"170f07",x"3d2310",x"150e07",x"2d1a0c",x"371f0e",x"23150a",x"23150a",x"2a1b10",x"2a1b10",x"321e11",x"341f0f",x"331e0f",x"351e0f",x"2d190d",x"2a170a",x"180f07",x"432712",x"514135",x"503019",x"412816",x"382212",x"412615",x"402514",x"362010",x"323232",x"454545",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"545454",x"4b4b4b",x"343434",x"323232",x"333333",x"333333",x"323232",x"3b3937",x"383736",x"3e3c39",x"333333",x"323232",x"303030",x"000000",x"000000",x"000000",x"303030",x"2e2e2e",x"303030",x"313131",x"434343",x"494949",x"5d5c5c",x"575656",x"464646",x"2b2b2b",x"353535",x"373737",x"464646",x"646464",x"5a5a5a",x"5a5a59",x"545454",x"464646",x"333333",x"323232",x"474747",x"545454",x"646464",x"504f4e",x"575656",x"515151",x"414141",x"343434",x"3e3e3e",x"000000",x"000000",x"452611",x"452611",x"37200f",x"3e2310",x"3d2411",x"351d0d",x"371f0e",x"402512",x"402511",x"3c220f",x"3f2411",x"3f2410",x"201309",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"181007",x"1f1408",x"1d1208",x"1e1308",x"1f1408",x"191107",x"201408",x"211508",x"201508",x"231608",x"2a1b09",x"2b1b09",x"261809",x"2d1c09",x"271909",x"241708",x"1e1308",x"231608",x"201408",x"2a1a09",x"2a1b09",x"241708",x"231608",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"554b41",x"554b41",x"3f342b",x"382c22",x"482d1b",x"41240f",x"3f2411",x"361d0d",x"341c0b",x"412611",x"432611",x"432611",x"3c210e",x"361c0c",x"432711",x"4a2912",x"51483e",x"42382e",x"3c2e24",x"462e20",x"462e20",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"251509",x"251509",x"150e07",x"150e07",x"000000",x"000000",x"3e2310",x"452812",x"4c3425",x"3e2d21",x"4b4239",x"150e07",x"150e07",x"150e07",x"150e07",x"28190c",x"150e07",x"150e07",x"150e07",x"150e07",x"37291f",x"35281e",x"362e26",x"362e26",x"000000",x"534337",x"534337",x"371f0e",x"28170a",x"241509",x"28160a",x"29170a",x"241509",x"231409",x"26160a",x"241509",x"1a1008",x"26160a",x"241509",x"251509",x"25150a",x"27160a",x"241509",x"231409",x"26160a",x"241509",x"221409",x"211309",x"201308",x"201309",x"1f1208",x"241509",x"241509",x"241509",x"221409",x"241509",x"170f07",x"201309",x"211309",x"26160a",x"201309",x"1c1108",x"25160a",x"25150a",x"1f1208",x"221409",x"28170a",x"1e1208",x"231409",x"211309",x"211309",x"201208",x"221409",x"231409",x"211309",x"211309",x"1f1208",x"221409",x"26160a",x"29170a",x"1a1008",x"1c1108",x"41230f",x"160e07",x"8b6645",x"886242",x"815e40",x"7d5b3c",x"7f5d3f",x"846244",x"856344",x"856344",x"836143",x"816042",x"896647",x"866445",x"805e40",x"78573b",x"7c5b3e",x"866345",x"826042",x"846244",x"815d40",x"826041",x"816041",x"846142",x"7d5b3e",x"7b5a3c",x"7a583a",x"7b593b",x"7c593b",x"856243",x"7f5c3e",x"815d3f",x"805d3e",x"7f5c3d",x"836040",x"7e5b3d",x"79593c",x"765538",x"7f5d3f",x"826143",x"826043",x"8c6848",x"8b6747",x"896747",x"8c6848",x"886544",x"846142",x"7a593c",x"815f41",x"856244",x"8a6646",x"896547",x"846142",x"896547",x"876444",x"886443",x"825f3f",x"5a4c41",x"432612",x"150e07",x"150e07",x"150e07",x"442815",x"442815",x"352a21",x"4f2d15",x"4f2d15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482913",x"482913",x"371f0e",x"402511",x"37200e",x"150e07",x"36200f",x"2b190b",x"301c0c",x"341e0d",x"211409",x"29170a",x"2a170a",x"482913",x"482913",x"343434",x"323232",x"353535",x"393939",x"393939",x"333333",x"313131",x"323232",x"343434",x"333333",x"323333",x"323232",x"323232",x"333333",x"323232",x"323232",x"323232",x"323232",x"3e3e3d",x"333333",x"333333",x"323232",x"5d5c5c",x"323231",x"000000",x"000000",x"323232",x"323232",x"333333",x"323232",x"4d4843",x"313131",x"313131",x"323232",x"333333",x"353535",x"333333",x"323232",x"313131",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a351a",x"5a351a",x"543017",x"331d0e",x"4d2e16",x"402310",x"402511",x"150e07",x"38200f",x"3c230f",x"38200e",x"381f0e",x"231409",x"3f2310",x"2e180a",x"4f4338",x"3f230f",x"3a210f",x"1f1208",x"150e07",x"3d2411",x"2b1a0c",x"180f07",x"2c180b",x"150e07",x"522f17",x"150e07",x"150e07",x"444444",x"5a5a5a",x"5d5d5d",x"626262",x"5d5d5d",x"5d5d5d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432711",x"432711",x"1f1308",x"1a1107",x"191007",x"150e07",x"150e07",x"271609",x"271609",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f392b",x"4f392b",x"150e07",x"422712",x"381f0d",x"25160a",x"150e07",x"311c0d",x"2d1a0c",x"150e07",x"38200e",x"311d0d",x"311d0d",x"2b1b10",x"2b1b10",x"311e11",x"352011",x"311d0f",x"361f0f",x"2c190c",x"27160a",x"180f07",x"3f2511",x"543e2f",x"4e2f1a",x"452b18",x"472a17",x"422815",x"432715",x"2a190c",x"333333",x"383838",x"444444",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d3d3d",x"474747",x"545454",x"313131",x"313131",x"333333",x"333333",x"000000",x"000000",x"000000",x"373635",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"303030",x"303030",x"303030",x"494949",x"4c4d4c",x"4e4e4f",x"4d4d4d",x"4b4b4b",x"414141",x"2b2b2b",x"000000",x"000000",x"5c5c5c",x"626363",x"5a5a5a",x"575757",x"4c4c4c",x"333333",x"000000",x"000000",x"646464",x"666665",x"5a5a59",x"5f5f5f",x"515151",x"4b4b4b",x"363636",x"000000",x"000000",x"000000",x"4b2b13",x"4b2b13",x"341e0e",x"39200f",x"38210f",x"3a200e",x"3c2310",x"412612",x"3c210f",x"3b2210",x"3f2411",x"3d2310",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"201408",x"1b1108",x"1b1108",x"191007",x"1d1308",x"1f1308",x"231608",x"1c1208",x"211508",x"2a1b09",x"2f1d0a",x"201408",x"271809",x"221608",x"241708",x"201508",x"231608",x"271809",x"231608",x"271909",x"1d1208",x"1d1308",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"50463c",x"50463c",x"423930",x"362a20",x"4c301e",x"41240e",x"3b210f",x"321b0b",x"261207",x"3e220f",x"3f2310",x"432611",x"3f230f",x"3e220f",x"3f230f",x"472710",x"534a3f",x"44392f",x"403126",x"4e3321",x"4e3321",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"28160a",x"1d1108",x"150e07",x"150e07",x"000000",x"000000",x"482913",x"482913",x"4d3526",x"3e2e22",x"463c32",x"150e07",x"150e07",x"150e07",x"150e07",x"24150a",x"150e07",x"150e07",x"150e07",x"1a1008",x"33251c",x"34261c",x"3a3128",x"3a3128",x"000000",x"554337",x"554337",x"321c0d",x"26160a",x"2c190b",x"241409",x"231409",x"251509",x"2c190b",x"2b180b",x"27160a",x"27170a",x"24150a",x"27160a",x"231409",x"29180b",x"26160a",x"28160a",x"29170a",x"27170a",x"251509",x"231409",x"201309",x"1f1209",x"201309",x"1f1309",x"25160a",x"211309",x"25160a",x"231509",x"25160a",x"221409",x"25150a",x"1f1209",x"26160a",x"201309",x"231409",x"1d1208",x"27170a",x"25160a",x"26160a",x"221409",x"1b1108",x"28170b",x"28170b",x"231509",x"241509",x"24150a",x"24150a",x"201309",x"201309",x"241509",x"241509",x"221409",x"25160a",x"25150a",x"2e1a0b",x"472812",x"160e07",x"7c5a3b",x"785538",x"7b5a3b",x"725235",x"7c593b",x"815e40",x"805e3e",x"826041",x"7c5b3e",x"815f40",x"79573a",x"846244",x"835f40",x"7f5d3f",x"7d5b3e",x"856143",x"846042",x"7e5c3e",x"856142",x"805f40",x"7d5b3e",x"7a593c",x"7b5a3d",x"7b5a3d",x"825e3d",x"7d5a3b",x"7b583a",x"7a593b",x"805d3f",x"7f5b3d",x"7d5b3c",x"765538",x"715236",x"745236",x"755538",x"725234",x"745438",x"805e3f",x"755539",x"866343",x"846243",x"846142",x"7e5b3d",x"826143",x"815e40",x"79593c",x"805d3f",x"815e40",x"846041",x"805d3f",x"886344",x"866343",x"836041",x"856141",x"876443",x"57493d",x"4b2b14",x"150e07",x"150e07",x"150e07",x"4a2c18",x"4a2c18",x"392c22",x"4e2d15",x"4e2d15",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2a13",x"4a2a13",x"3a210f",x"422712",x"402612",x"150e07",x"362210",x"150e07",x"27170a",x"351f0f",x"2b190b",x"26150a",x"2c180b",x"432511",x"432511",x"000000",x"323232",x"373737",x"3b3b3b",x"363636",x"323232",x"313131",x"323232",x"333333",x"323232",x"313131",x"343434",x"333333",x"2f2f2f",x"323232",x"323131",x"333333",x"454545",x"444444",x"32302f",x"333333",x"323232",x"4d4d4d",x"000000",x"000000",x"373737",x"373737",x"333333",x"333231",x"454545",x"4b4641",x"323232",x"323232",x"343434",x"333333",x"323232",x"3a3a3a",x"474747",x"4d4d4d",x"323130",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563218",x"563218",x"4c2b13",x"341e0e",x"4d2e16",x"3a200e",x"3b210f",x"150e07",x"3a210f",x"371f0e",x"341e0d",x"39210f",x"311d0d",x"3f2310",x"2f190b",x"54483d",x"402310",x"3c220f",x"3b210f",x"3f2411",x"2a190b",x"37200f",x"2c190b",x"2f1b0c",x"150e07",x"4b2a13",x"150e07",x"150e07",x"373737",x"373737",x"3f3f3f",x"3d3d3d",x"4a4a4a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2410",x"3e2410",x"1e1308",x"1c1208",x"191008",x"150e07",x"150e07",x"331c0c",x"331c0c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c382a",x"4c382a",x"150e07",x"4a2b15",x"321b0c",x"412511",x"3b2310",x"2b190c",x"301c0d",x"3d2310",x"341d0d",x"301c0d",x"301c0d",x"2a1b10",x"2a1b10",x"311e11",x"351f11",x"372111",x"331d0e",x"28180b",x"2f1a0b",x"180f08",x"3d2310",x"543f31",x"4d2f1a",x"472c18",x"432817",x"452915",x"3c2414",x"2b190c",x"313131",x"2c2c2c",x"323232",x"4a4a4a",x"4d4d4d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c5c5c",x"606060",x"3d3d3d",x"323232",x"353535",x"313131",x"313131",x"5f5f5f",x"5e5d5d",x"4b4b4b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e4e4f",x"4d4d4d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"626363",x"5a5a5a",x"595959",x"636363",x"636262",x"676767",x"505050",x"535353",x"454545",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2a12",x"4b2a12",x"3e2410",x"3c220f",x"3a2110",x"381f0e",x"381f0e",x"3e2411",x"3b220f",x"3d2310",x"402411",x"402511",x"201309",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1408",x"211508",x"191007",x"1c1208",x"1b1108",x"191007",x"1c1208",x"211508",x"1f1408",x"291a09",x"2b1b09",x"201508",x"221508",x"1e1308",x"1d1308",x"1c1208",x"1e1308",x"221608",x"231608",x"201508",x"221608",x"1e1308",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"17110a",x"17110a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d443b",x"4d443b",x"3d342b",x"352b22",x"482e1e",x"3c210d",x"39200e",x"361d0c",x"241106",x"442712",x"3c210e",x"3f230f",x"402410",x"3f230f",x"3c220f",x"442610",x"574e43",x"473e34",x"44362b",x"4e3424",x"4e3424",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"211309",x"211309",x"1e1108",x"1e1108",x"000000",x"000000",x"472913",x"472913",x"4c3425",x"3f2d20",x"4b4238",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"150e07",x"170f07",x"2b2018",x"332419",x"362c23",x"362c23",x"000000",x"534337",x"534337",x"341d0d",x"27160a",x"251509",x"251509",x"28160a",x"26160a",x"241509",x"241509",x"251509",x"1c1108",x"27160a",x"29170a",x"25160a",x"26160a",x"26160a",x"251509",x"221409",x"231409",x"241509",x"241509",x"241509",x"1f1208",x"1a1008",x"1f1309",x"170f07",x"1d1108",x"231409",x"1e1108",x"201308",x"1c1108",x"1f1208",x"241509",x"1c1108",x"231409",x"221409",x"27170a",x"211409",x"251509",x"221409",x"211309",x"26160a",x"29170a",x"27170a",x"231509",x"231509",x"231409",x"231409",x"150e07",x"28180b",x"23150a",x"231509",x"25160a",x"24150a",x"27170a",x"27170a",x"4b2b14",x"160f07",x"7b593a",x"7b593b",x"735335",x"6f5033",x"775739",x"725237",x"79573c",x"7b593d",x"775639",x"79573b",x"7a583c",x"755438",x"7a593d",x"7e5c3f",x"805f40",x"876446",x"836042",x"7e5c3e",x"79583a",x"735436",x"7b593c",x"755538",x"755539",x"7a593d",x"735336",x"815c3f",x"7c593c",x"79573a",x"79573a",x"765538",x"715135",x"745437",x"735436",x"745437",x"705033",x"725335",x"705135",x"725237",x"745439",x"7a583c",x"825f3f",x"7d5a3d",x"7e5b3d",x"7a583b",x"745439",x"7e5c3f",x"816041",x"846243",x"886343",x"815d3e",x"79583a",x"785739",x"825e3f",x"7c5a3c",x"805d3f",x"54463a",x"40220e",x"150e07",x"150e07",x"27160b",x"4c2e19",x"4c2e19",x"342a21",x"4d2c14",x"4d2c14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4b2b14",x"4b2b14",x"3d2310",x"3c2311",x"321e0e",x"29190c",x"35210f",x"150e07",x"241509",x"28180b",x"2f1b0c",x"28170a",x"2d1a0c",x"3f220e",x"3f220e",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"323232",x"333333",x"333333",x"323232",x"333333",x"333333",x"313232",x"333333",x"323232",x"323232",x"454545",x"505050",x"636363",x"525252",x"4f4f4f",x"666666",x"000000",x"000000",x"323232",x"323232",x"474747",x"616160",x"4e4e4e",x"545454",x"515151",x"515151",x"4b4b4b",x"494949",x"323232",x"626262",x"444444",x"313131",x"333333",x"343434",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"512f16",x"512f16",x"492812",x"2e1a0c",x"442712",x"3a200e",x"321c0d",x"2f1b0c",x"3f2411",x"3e2411",x"26170a",x"29180b",x"351f0e",x"422511",x"341c0c",x"4b3e33",x"40220f",x"361e0d",x"381f0e",x"38210f",x"2f1c0d",x"39210f",x"39200f",x"39210f",x"150e07",x"4c2a13",x"150e07",x"150e07",x"323232",x"323232",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"28190a",x"28190a",x"1c1208",x"160f07",x"150e07",x"150e07",x"150e07",x"351e0d",x"351e0d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3628",x"4d3628",x"150e07",x"452812",x"2e190a",x"3e2310",x"3b2210",x"25160a",x"2e1b0c",x"371f0e",x"351e0d",x"27170b",x"27170b",x"2a1a0f",x"2a1a0f",x"301e11",x"331f10",x"372111",x"331c0e",x"2f1b0d",x"2d1a0b",x"180f07",x"3b200f",x"513e30",x"4f311b",x"4b2f1a",x"432917",x"422817",x"3f2514",x"372010",x"323232",x"333333",x"343434",x"444444",x"4a4a4a",x"383838",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b4b4b",x"4d4d4d",x"5c5c5c",x"333333",x"323232",x"323232",x"323232",x"2f3030",x"5d5d5d",x"5f5f5f",x"616161",x"5f5f5f",x"525252",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e4e4e",x"555555",x"5d5d5d",x"636363",x"666666",x"565656",x"4f4f4e",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2b14",x"4c2b14",x"321c0d",x"3a200f",x"3b220f",x"371f0e",x"351e0d",x"321d0d",x"39210f",x"3d2310",x"3c220f",x"412611",x"1f1209",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"191007",x"191007",x"1d1208",x"160f07",x"181007",x"1d1308",x"1d1308",x"1d1308",x"191007",x"1a1107",x"281a09",x"241608",x"1d1308",x"1c1208",x"1e1308",x"201408",x"170f07",x"1b1108",x"1b1108",x"1e1308",x"1c1208",x"170f07",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"18110a",x"18110a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494037",x"494037",x"3d342c",x"3a2e25",x"472e1e",x"3f230e",x"321b0c",x"3b200e",x"241106",x"412511",x"3b200e",x"3e230f",x"3f230f",x"402410",x"3c210e",x"472711",x"554c42",x"483d33",x"45362a",x"513624",x"513624",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"27160a",x"27160a",x"29170a",x"29170a",x"000000",x"000000",x"492913",x"492913",x"4a3425",x"3e2d21",x"4a4037",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"150e07",x"332216",x"2f2116",x"352b23",x"352b23",x"000000",x"4b3e34",x"4b3e34",x"341d0d",x"2a180b",x"26160a",x"27160a",x"221409",x"221409",x"241509",x"211409",x"241509",x"27160a",x"251509",x"241509",x"241509",x"221409",x"231509",x"1e1208",x"231409",x"24150a",x"1e1208",x"211309",x"1d1208",x"221409",x"191008",x"150e07",x"1c1108",x"1f1309",x"1b1108",x"231409",x"27170b",x"25160a",x"201309",x"231509",x"1f1309",x"231409",x"201309",x"1f1209",x"150e07",x"28170b",x"29180b",x"28170b",x"28170b",x"26170a",x"27170a",x"2b190b",x"29180b",x"27160a",x"241409",x"241409",x"231409",x"28180b",x"28180b",x"2b190c",x"25150a",x"26160a",x"26160a",x"4e2d16",x"180f07",x"825f41",x"7e5c3f",x"7c5a3d",x"715136",x"735337",x"78563a",x"745337",x"7c5a3c",x"7c5a3c",x"79583d",x"7e5c3f",x"7b5a3d",x"7c5b3e",x"805e40",x"7d5c3e",x"7d5b3e",x"815e40",x"725136",x"704e34",x"775538",x"7d5b3c",x"7b5a3d",x"785639",x"7a583c",x"7b5a3d",x"7d5b3e",x"826042",x"805d3f",x"7d5c3e",x"7c5a3b",x"735334",x"7e5c3d",x"7d5b3e",x"79583c",x"735338",x"745438",x"715136",x"755439",x"6e5034",x"7e5c3e",x"805d3e",x"805d41",x"7d5b3e",x"7b5a3d",x"866343",x"846243",x"896544",x"846041",x"866143",x"7a583a",x"775337",x"7a583a",x"7e5c3e",x"7d5c3e",x"765538",x"4d3e33",x"4d2c14",x"150e07",x"150e07",x"29170b",x"4e2f1a",x"4e2f1a",x"322921",x"4a2913",x"4a2913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4e2d16",x"4e2d16",x"3b220f",x"3d2411",x"3b2310",x"2e1c0d",x"3b2512",x"150e07",x"1c1108",x"2f1c0d",x"39200f",x"311c0c",x"321c0c",x"462711",x"462711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"333333",x"333333",x"313232",x"333333",x"000000",x"000000",x"000000",x"636363",x"636363",x"525252",x"4f4f4f",x"666666",x"575757",x"595959",x"525252",x"323232",x"474747",x"595959",x"545454",x"4d4d4d",x"3a3a3a",x"333333",x"333333",x"343434",x"313131",x"605b56",x"3a3a3a",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"543017",x"543017",x"4a2912",x"341f0e",x"472913",x"432712",x"422612",x"301b0c",x"3f2511",x"29180b",x"2e1b0c",x"361f0e",x"3b2210",x"482913",x"371f0e",x"43372d",x"3e220f",x"361e0d",x"2f1b0c",x"3d2411",x"3d2311",x"150e07",x"321d0d",x"3a210f",x"150e07",x"4b2a13",x"150e07",x"150e07",x"333333",x"333333",x"323232",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"160f07",x"160f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"301b0b",x"301b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523828",x"523828",x"150e07",x"432711",x"29160a",x"341d0d",x"3a200f",x"3b210e",x"150e07",x"2f1b0c",x"341d0d",x"311c0d",x"311c0d",x"291a10",x"291a10",x"2f1d11",x"321d0f",x"372011",x"351e0f",x"2e1a0d",x"301c0c",x"180f07",x"3e2310",x"513d30",x"472c19",x"4a2e19",x"412716",x"412716",x"3e2515",x"2c1a0d",x"2c1a0d",x"323232",x"3d3d3d",x"323333",x"323232",x"313131",x"5d5d5d",x"646464",x"4e4e4e",x"3f3f3f",x"434343",x"505050",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"393939",x"535353",x"4b4b4b",x"333333",x"323232",x"323232",x"313131",x"313131",x"303030",x"333333",x"333333",x"5c5c5c",x"525252",x"333333",x"595959",x"555555",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"595959",x"484848",x"505050",x"545454",x"555555",x"5b5b5b",x"333333",x"323232",x"343434",x"534d46",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2b14",x"4b2b14",x"3a200e",x"381f0e",x"351e0d",x"351d0d",x"2e1a0b",x"301a0b",x"351f0e",x"3c210f",x"39200e",x"3e2411",x"1c1108",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1408",x"1f1408",x"1e1308",x"1d1308",x"1b1208",x"191007",x"181007",x"1d1308",x"1a1107",x"160e07",x"180f07",x"150e07",x"160f07",x"160f07",x"1a1107",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a4138",x"4a4138",x"3f352d",x"382c23",x"4d3220",x"3e230f",x"351d0c",x"351d0c",x"231107",x"3f2310",x"381e0d",x"402410",x"3f2410",x"442711",x"3f220f",x"482812",x"554c42",x"463d35",x"43342a",x"503523",x"503523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1208",x"1f1208",x"29170a",x"29170a",x"000000",x"000000",x"432712",x"432712",x"4d3526",x"3e2c1f",x"4d443b",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"150e07",x"150e07",x"150e07",x"1a1008",x"322115",x"2b2017",x"31281f",x"31281f",x"000000",x"54463c",x"54463c",x"3b2210",x"371f0e",x"331d0d",x"321d0d",x"2a180b",x"2f1a0b",x"2d190b",x"2f1b0c",x"2e1a0c",x"321c0d",x"201309",x"2e1a0b",x"26160a",x"2d190b",x"2e1a0b",x"2c180b",x"2b180b",x"2e1b0c",x"2e1a0c",x"2e1a0c",x"2a170a",x"27160a",x"28160a",x"201208",x"231409",x"301b0c",x"231509",x"2e1a0b",x"2d1a0c",x"2e1a0b",x"2c190b",x"2b190c",x"231509",x"2d1a0c",x"2c1a0b",x"321c0d",x"2a190b",x"2c1a0c",x"2c1a0c",x"2e1b0c",x"301c0d",x"311c0d",x"331e0e",x"37200f",x"2d1a0c",x"2e1b0d",x"2a180b",x"261509",x"2a170a",x"2d1a0c",x"2f1c0d",x"2c1a0b",x"211409",x"311c0d",x"2c190c",x"4a2a13",x"160e07",x"886243",x"886343",x"825e3f",x"7c593b",x"825e3f",x"805c3e",x"886342",x"7c5a3c",x"8c6745",x"856041",x"835e3f",x"7c5a3b",x"8b6443",x"8b6645",x"8c6645",x"825e3f",x"856040",x"825e3c",x"886342",x"876343",x"7f5b3e",x"856143",x"8a6645",x"876445",x"846142",x"805c3e",x"866142",x"866041",x"815d3e",x"815d3e",x"855f3f",x"815d3d",x"805c3e",x"7e5c3d",x"7f5b3d",x"7f5b3d",x"835e3f",x"7e5a3d",x"866243",x"846040",x"8b6645",x"846041",x"775639",x"775438",x"8a6443",x"8e6847",x"8a6444",x"815d3f",x"886343",x"8c6544",x"8e6745",x"8d6846",x"866142",x"866243",x"846142",x"493d32",x"522f16",x"150e07",x"150e07",x"211409",x"4c2e19",x"4c2e19",x"2c251e",x"4b2913",x"4b2913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"472914",x"472914",x"3b220f",x"3f2411",x"3a2110",x"301d0e",x"382511",x"150e07",x"241509",x"2b190b",x"311c0c",x"231509",x"2a180b",x"492913",x"492913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"656565",x"656565",x"454545",x"323232",x"333333",x"575757",x"595959",x"525252",x"404040",x"353535",x"4f4f4f",x"3f3f3f",x"383838",x"4d4d4d",x"565656",x"3d3d3d",x"333333",x"383838",x"333333",x"595959",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"502e16",x"502e16",x"4b2a14",x"2f1c0d",x"4a2b15",x"442813",x"3d2310",x"321c0c",x"412612",x"3c220f",x"301c0d",x"38200f",x"3a210f",x"482913",x"38200e",x"40342a",x"41230f",x"3f2410",x"3a200e",x"2e1a0c",x"381f0e",x"150e07",x"38200f",x"3d2310",x"150e07",x"4e2c15",x"150e07",x"150e07",x"323232",x"323232",x"333333",x"464646",x"464646",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2e1b0c",x"2e1b0c",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"201309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523a2a",x"523a2a",x"150e07",x"442611",x"281408",x"341d0d",x"26160a",x"3c210f",x"150e07",x"2c190b",x"37210f",x"2b1b0c",x"2b1b0c",x"28190f",x"28190f",x"2f1d11",x"301c0f",x"341e10",x"382010",x"2e190b",x"301c0c",x"180f07",x"3d220f",x"574132",x"472c1b",x"4b2f1b",x"482d1b",x"412816",x"402615",x"341f10",x"341f10",x"333333",x"434343",x"444545",x"333333",x"303030",x"3f3f3f",x"616161",x"4e4e4e",x"3f3f3f",x"434343",x"4f4f4f",x"323232",x"333333",x"434343",x"474747",x"4e4e4e",x"4c4c4c",x"5c5c5c",x"4b4b4b",x"484848",x"333333",x"333434",x"484848",x"323232",x"333231",x"323232",x"323232",x"696969",x"383838",x"323232",x"343434",x"333333",x"363636",x"5c5c5c",x"616161",x"595959",x"656565",x"606060",x"5d5d5d",x"000000",x"000000",x"000000",x"000000",x"555555",x"3f3f3f",x"363636",x"363636",x"3a3a3a",x"333333",x"595959",x"484949",x"575757",x"565656",x"363331",x"313131",x"323232",x"313131",x"323232",x"343434",x"323232",x"4c4742",x"43403d",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442711",x"442711",x"3c220f",x"361e0d",x"381f0e",x"2c180a",x"251308",x"2e1a0b",x"36200f",x"3d2310",x"3c210f",x"3c210f",x"1f1309",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1208",x"170f07",x"1b1108",x"1c1208",x"1d1308",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"453d34",x"453d34",x"3e332a",x"3c3027",x"513423",x"381e0d",x"31190b",x"3b210f",x"261308",x"3c210f",x"371e0d",x"3e230f",x"341c0c",x"422611",x"3d220f",x"482811",x"51473e",x"453b31",x"403229",x"503523",x"503523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1a1008",x"1a1008",x"201309",x"201309",x"000000",x"000000",x"432611",x"432611",x"3e2b21",x"3e2e23",x"4e443a",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"191008",x"332216",x"322317",x"312a23",x"312a23",x"000000",x"56463a",x"56463a",x"3d210e",x"3c200e",x"442611",x"40230f",x"3f210e",x"442510",x"462711",x"422510",x"432510",x"3e210e",x"3d210e",x"3f230f",x"422511",x"442611",x"422611",x"442711",x"452712",x"492a14",x"442712",x"4c2c15",x"4d2e16",x"472a14",x"422812",x"412511",x"3c230f",x"402511",x"432611",x"432611",x"442712",x"442a14",x"4d2d15",x"492a13",x"4c2c15",x"462812",x"462913",x"462914",x"4c2c14",x"4f2e16",x"4c2d15",x"482914",x"452711",x"472812",x"482913",x"4e2c15",x"4a2a14",x"492a14",x"4c2b15",x"4c2b14",x"4a2913",x"492913",x"4b2b13",x"4a2a13",x"452611",x"472711",x"432510",x"462711",x"482912",x"2d1a0b",x"2d190b",x"331d0c",x"39210f",x"36200e",x"351f0d",x"351f0d",x"39210e",x"37210d",x"2a190b",x"301c0b",x"39210e",x"3a220f",x"3a220e",x"3b230e",x"3c230f",x"402510",x"432810",x"331d0d",x"3c2310",x"38200e",x"321c0d",x"301a0b",x"341d0d",x"371f0e",x"2d190b",x"3b220f",x"321d0c",x"301b0b",x"301b0b",x"28160a",x"2f1b0b",x"2f190b",x"311a0b",x"311b0b",x"331c0c",x"361d0d",x"341d0c",x"361e0d",x"351d0c",x"321c0c",x"39200e",x"3c220f",x"3d230f",x"3f2510",x"432712",x"412612",x"412611",x"402411",x"3c210f",x"381f0e",x"3f2310",x"432813",x"432812",x"442712",x"503d30",x"462711",x"150e07",x"150e07",x"201409",x"4a2c18",x"4a2c18",x"35281e",x"4c2a13",x"4c2a13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482914",x"482914",x"37200f",x"3c2311",x"3b2311",x"3f2612",x"3a2411",x"321d0d",x"221409",x"2d190b",x"37200f",x"211309",x"28170a",x"442711",x"442711",x"000000",x"333333",x"323232",x"4b4b4b",x"4e4e4e",x"525252",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"423f3c",x"423f3c",x"494540",x"313131",x"313131",x"333333",x"323232",x"333333",x"333333",x"343434",x"323232",x"323232",x"333333",x"373634",x"393836",x"333333",x"313131",x"323232",x"323232",x"343434",x"343434",x"323232",x"3a3a3a",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"543218",x"543218",x"533117",x"36200f",x"4d2e16",x"422712",x"3a210f",x"301b0c",x"432712",x"39200e",x"2d1a0c",x"39200f",x"3a210f",x"472813",x"361e0e",x"48382c",x"3e220f",x"3a210f",x"381f0e",x"311c0d",x"412512",x"1b1108",x"3a2210",x"39200f",x"150e07",x"472711",x"150e07",x"150e07",x"414141",x"414141",x"494949",x"5d5d5d",x"5f5f5f",x"5f5f5f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"331d0d",x"331d0d",x"231608",x"160f07",x"150e07",x"150e07",x"160f07",x"1b1008",x"1b1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563e2d",x"563e2d",x"150e07",x"432612",x"2b1508",x"371f0e",x"29180b",x"38200e",x"150e07",x"341e0d",x"3a2110",x"26160a",x"26160a",x"27190f",x"27190f",x"2e1c11",x"311d0f",x"2c180c",x"382010",x"2e190b",x"2f1b0c",x"180f07",x"39200e",x"543e2f",x"4b2e1a",x"482d1a",x"482d1a",x"442b18",x"422816",x"2b1a0d",x"2b1a0d",x"000000",x"494949",x"303031",x"313131",x"323232",x"646464",x"625f5c",x"303030",x"323232",x"313131",x"333333",x"333333",x"343434",x"393939",x"474747",x"4e4e4e",x"4c4c4c",x"5b5b5b",x"4a4a4a",x"313131",x"303030",x"333333",x"5f5e5e",x"434343",x"323232",x"000000",x"000000",x"323232",x"323232",x"333333",x"333333",x"323232",x"313131",x"333333",x"5a5a5a",x"646464",x"606060",x"606060",x"5d5d5d",x"616060",x"5c5c5c",x"606060",x"535353",x"555555",x"484848",x"363636",x"363636",x"3a3a3a",x"333333",x"595959",x"5a5a5a",x"505050",x"323232",x"2f3030",x"343434",x"323232",x"323232",x"313131",x"333333",x"323232",x"373635",x"43403d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442611",x"442611",x"351d0d",x"381f0e",x"341d0d",x"2b170a",x"251308",x"311b0c",x"3c2311",x"361f0e",x"3f2311",x"3b200e",x"191008",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"191008",x"1a1008",x"190f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"161009",x"161009",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"473e35",x"473e35",x"433a31",x"42362d",x"513626",x"381e0d",x"361d0c",x"3a200e",x"271308",x"432612",x"3b200e",x"3d220f",x"341c0c",x"402410",x"381f0d",x"41230f",x"463e35",x"3e3229",x"413227",x"523625",x"523625",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1f1209",x"1f1209",x"170f07",x"170f07",x"000000",x"000000",x"3d220f",x"3d220f",x"3c291f",x"413024",x"4b4138",x"150e07",x"150e07",x"150e07",x"150e07",x"27180b",x"150e07",x"150e07",x"150e07",x"190f08",x"342215",x"302217",x"342c23",x"342c23",x"000000",x"000000",x"56463a",x"443429",x"462712",x"39200e",x"331d0c",x"3b210f",x"331c0c",x"321b0b",x"2e190a",x"2e190b",x"331c0c",x"311b0b",x"311c0c",x"2f1b0c",x"341d0d",x"301b0c",x"301b0b",x"2f1a0b",x"2e190b",x"2e190b",x"2c190b",x"2f1a0b",x"2d190b",x"2e1a0b",x"311c0c",x"2f1a0b",x"311c0c",x"2f1b0c",x"2d190b",x"29160a",x"301b0c",x"321d0d",x"2b180b",x"341d0d",x"2e1a0b",x"301b0c",x"2e1a0b",x"321c0d",x"331d0d",x"331c0d",x"331c0d",x"301b0c",x"2e1a0b",x"301c0c",x"301b0c",x"2e1a0c",x"301b0c",x"301c0c",x"2e1a0b",x"2f1b0c",x"2d190b",x"28160a",x"2e1a0b",x"2c190b",x"2a170a",x"2a170a",x"2b180b",x"2d190b",x"1a1008",x"2d190b",x"331d0c",x"39210f",x"36200e",x"351f0d",x"351f0d",x"39210e",x"37210d",x"2a190b",x"301c0b",x"39210e",x"3a220f",x"3a220e",x"3b230e",x"3c230f",x"402510",x"432810",x"331d0d",x"3c2310",x"38200e",x"321c0d",x"301a0b",x"341d0d",x"371f0e",x"2d190b",x"3b220f",x"321d0c",x"301b0b",x"301b0b",x"28160a",x"2f1b0b",x"2f190b",x"311a0b",x"311b0b",x"331c0c",x"361d0d",x"341d0c",x"361e0d",x"351d0c",x"321c0c",x"39200e",x"3c220f",x"3d230f",x"3f2510",x"432712",x"412612",x"412611",x"402411",x"3c210f",x"381f0e",x"3f2310",x"432813",x"432812",x"442712",x"351d0d",x"351d0d",x"150e07",x"150e07",x"160f07",x"2b1c11",x"2b1c11",x"36291f",x"311b0b",x"311b0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"432611",x"432611",x"38200f",x"341e0d",x"3b2310",x"3e2511",x"38200e",x"37210f",x"2a190b",x"2a180b",x"351e0d",x"231409",x"28170a",x"442611",x"442611",x"333232",x"333333",x"323232",x"4b4b4b",x"4e4e4e",x"565656",x"5e5e5e",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"333333",x"4f4f4f",x"000000",x"323232",x"333333",x"323232",x"2f2f2f",x"343434",x"3d3d3d",x"353535",x"333333",x"323232",x"333333",x"323232",x"323232",x"313131",x"323232",x"343434",x"3e3b39",x"585756",x"323232",x"333333",x"333333",x"333333",x"363636",x"3b3a3a",x"323232",x"3a3a3a",x"3e3e3e",x"3e3e3e",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"29170a",x"29170a",x"4e2c15",x"4e2c15",x"523017",x"382110",x"4d2e16",x"3b2210",x"3d2310",x"361e0d",x"402511",x"3e230f",x"2c190b",x"37200f",x"39210f",x"462812",x"361e0d",x"4a382d",x"412410",x"351d0d",x"2b180b",x"221409",x"3a2210",x"180f08",x"211409",x"37200f",x"150e07",x"482812",x"150e07",x"150e07",x"4d4d4d",x"4d4d4d",x"3b3b3b",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"3d230f",x"221608",x"170f07",x"160e07",x"150e07",x"1f1408",x"231608",x"231608",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"553c2c",x"553c2c",x"150e07",x"482a14",x"2c1609",x"2a180b",x"231509",x"371f0e",x"150e07",x"1c1108",x"351f0e",x"2e1b0c",x"2e1b0c",x"27190f",x"27190f",x"2d1c10",x"311d10",x"2d190c",x"351e0f",x"2a170a",x"301c0c",x"180f07",x"2f1a0b",x"4d3a2d",x"4a2c18",x"412817",x"432a19",x"432a18",x"412918",x"2b1a0d",x"2b1a0d",x"000000",x"000000",x"282828",x"282828",x"585858",x"595959",x"62605e",x"343434",x"333333",x"323232",x"313131",x"333333",x"343434",x"313131",x"333333",x"343434",x"3a3a3a",x"656565",x"333333",x"595959",x"434343",x"323232",x"333333",x"605f5f",x"000000",x"000000",x"323232",x"323232",x"323232",x"3d3d3d",x"444444",x"333333",x"323232",x"333333",x"454545",x"323232",x"323232",x"5b5650",x"5a5a5a",x"686868",x"5c5c5c",x"606060",x"535353",x"474747",x"4d4d4d",x"333333",x"303030",x"313131",x"323232",x"363534",x"333333",x"323232",x"333333",x"333333",x"393939",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472712",x"472712",x"3a200e",x"351d0d",x"301a0b",x"2c170a",x"271408",x"331d0d",x"331e0e",x"371f0e",x"38200e",x"381f0e",x"201309",x"150e07",x"150e07",x"170f07",x"1d140d",x"1b1108",x"1d1108",x"1e1208",x"1e1208",x"1c1108",x"190f07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"17110a",x"171009",x"171009",x"17110a",x"1a130c",x"19130c",x"19120c",x"171009",x"17100a",x"17100a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"494037",x"494037",x"41382f",x"41362d",x"503727",x"361c0b",x"331b0b",x"3f2310",x"2f180a",x"3f2410",x"3a200e",x"402410",x"3e220f",x"3d220f",x"381f0d",x"3e210d",x"4d443b",x"473b31",x"47392e",x"533827",x"533827",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"3d220f",x"3d220f",x"3c291f",x"3d2d21",x"4d443a",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"170f07",x"322216",x"302116",x"352c24",x"352c24",x"000000",x"000000",x"403228",x"403228",x"422510",x"381f0e",x"371f0d",x"371e0d",x"351d0d",x"2e1a0b",x"2c180a",x"2d180a",x"2e190b",x"331c0c",x"331c0c",x"331c0d",x"311c0c",x"311c0c",x"2e190b",x"301a0b",x"2d180a",x"281609",x"29170a",x"2c180b",x"2d190b",x"2a170a",x"2c180a",x"2c190b",x"2f1a0b",x"2f1a0b",x"2e1a0b",x"311c0c",x"2e1a0b",x"321c0c",x"351e0d",x"321c0c",x"2c190b",x"2f1a0b",x"2c190b",x"301b0c",x"321c0d",x"331d0d",x"301b0c",x"2f1b0c",x"2d1a0b",x"301c0d",x"2f1b0c",x"2a180b",x"2f1b0c",x"341e0e",x"301b0c",x"301c0d",x"361f0e",x"231509",x"2e1a0c",x"2d190b",x"29180a",x"2a180b",x"2e1a0b",x"26160a",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452711",x"452711",x"150e07",x"150e07",x"170f07",x"422716",x"422716",x"2f251d",x"40230f",x"40230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"452611",x"452611",x"38200f",x"38200f",x"2c1a0c",x"331e0d",x"361f0e",x"150e07",x"2a190b",x"37200f",x"361f0e",x"231409",x"2c180b",x"422410",x"323232",x"323232",x"4f4f4f",x"585858",x"5a5a5a",x"555555",x"5f5f5f",x"5d5d5d",x"5c5c5c",x"000000",x"323232",x"323232",x"333333",x"323232",x"333333",x"606060",x"333333",x"313131",x"323232",x"323232",x"5d5d5d",x"5f5f5f",x"606060",x"595959",x"595959",x"3f3f3f",x"4a4a4a",x"545454",x"323232",x"313131",x"313131",x"323232",x"323232",x"333333",x"393939",x"3d3d3d",x"474747",x"4d4d4d",x"5a5a5a",x"5b5b5b",x"313131",x"393939",x"4b4b4b",x"3b3b3b",x"424242",x"595959",x"606060",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"4c2c14",x"4c2c14",x"543118",x"341e0e",x"482b15",x"402511",x"3f2512",x"2c180a",x"402511",x"3a210f",x"2d1a0c",x"3a210f",x"381f0e",x"462812",x"331c0c",x"3d332a",x"422410",x"3b210f",x"371e0d",x"150e07",x"3e2512",x"150e07",x"39210f",x"23150a",x"150e07",x"4d2c14",x"150e07",x"150e07",x"000000",x"333333",x"333333",x"333333",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1c0b",x"2f1c0b",x"201508",x"1d1208",x"150e07",x"170f07",x"1e1308",x"2c1b0a",x"2c1b0a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"553d2c",x"553d2c",x"150e07",x"432511",x"361d0c",x"3e2411",x"150e07",x"371f0e",x"150e07",x"2f1b0c",x"180f07",x"27160a",x"27160a",x"27190f",x"27190f",x"29190e",x"2c1a0e",x"331d0f",x"321c0e",x"2a170a",x"28170a",x"170f07",x"371f0e",x"534031",x"472b18",x"442b19",x"3f2818",x"3e2717",x"452a18",x"392212",x"392212",x"000000",x"000000",x"323232",x"323232",x"4a4641",x"333333",x"666666",x"5c5c5c",x"505050",x"333333",x"333333",x"323232",x"323232",x"323232",x"343434",x"484848",x"4a4a4a",x"4e4d4c",x"696969",x"606060",x"4a4a4a",x"333333",x"333333",x"333333",x"000000",x"000000",x"333333",x"333333",x"323232",x"323232",x"555555",x"5f5f5f",x"333333",x"363636",x"414140",x"353535",x"3b3a3a",x"59524c",x"353535",x"3e3e3e",x"3a3a3a",x"333333",x"313131",x"323232",x"323232",x"323232",x"333333",x"333333",x"323232",x"4f4f4f",x"6c6c6c",x"393939",x"333333",x"3c3c3c",x"4b4b4b",x"313131",x"343434",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2913",x"4b2913",x"3d220f",x"2f190b",x"321c0c",x"2e190b",x"311b0c",x"351f0f",x"442813",x"361f0d",x"37200f",x"311b0c",x"1c1108",x"483421",x"150e07",x"171008",x"1d140d",x"1d120a",x"1d1208",x"1f1208",x"1e1208",x"1d1108",x"191008",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f08",x"17110a",x"19130c",x"17110a",x"19120b",x"19130c",x"1a130c",x"19130c",x"18110a",x"17110a",x"17110a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"483f36",x"483f36",x"40352b",x"40342a",x"4a3123",x"351c0d",x"341b0b",x"3e2310",x"331a0b",x"3e2310",x"3d220f",x"412511",x"3c220f",x"3f2310",x"391f0d",x"43240f",x"51473d",x"41372e",x"423428",x"503523",x"503523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"3f2310",x"3f2310",x"503525",x"443529",x"574d43",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"191008",x"312116",x"2e2017",x"3d3229",x"3d3229",x"000000",x"000000",x"4b3a2d",x"4b3a2d",x"452611",x"341c0c",x"321c0b",x"341d0c",x"361e0d",x"351d0d",x"2f1a0b",x"301a0b",x"301a0b",x"321b0b",x"351d0d",x"301b0c",x"321c0c",x"2f1a0b",x"301a0b",x"2e190a",x"2e190b",x"2a170a",x"28160a",x"2a170a",x"2f1b0b",x"301b0b",x"301b0b",x"2f1b0c",x"301b0c",x"2f1b0c",x"331c0c",x"321b0c",x"321c0d",x"2c190b",x"361f0e",x"361f0e",x"311c0d",x"341e0d",x"301b0c",x"27160a",x"2a180b",x"2c190b",x"29180b",x"2b180b",x"2a180b",x"2f1b0c",x"2d1a0b",x"2f1b0b",x"311c0d",x"2f1b0c",x"301b0c",x"2b190b",x"2f1a0b",x"2d190b",x"29170a",x"2c190b",x"2d1a0c",x"2a180b",x"27170a",x"2c190b",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2a12",x"4b2a12",x"150e07",x"150e07",x"1a1008",x"3d2514",x"3d2514",x"28211a",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2912",x"4a2912",x"3a210f",x"402512",x"2c190b",x"26170a",x"38200f",x"150e07",x"2e1a0c",x"36200f",x"361f0e",x"2c190b",x"26160a",x"3f230f",x"333232",x"424242",x"5c5c5c",x"373737",x"323232",x"383838",x"4e4e4e",x"5b5b5b",x"5b5b5b",x"3e3e3e",x"32302f",x"323232",x"323232",x"343434",x"5e5e5e",x"696764",x"323232",x"494949",x"555555",x"444444",x"414141",x"3f3f3f",x"363636",x"323232",x"323232",x"656565",x"545454",x"5a5a5a",x"333333",x"333333",x"333333",x"313131",x"545454",x"585858",x"474747",x"494a4a",x"494a4a",x"444444",x"494949",x"454545",x"484848",x"494949",x"494949",x"515151",x"606060",x"606060",x"606060",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"361f0e",x"361f0e",x"522f16",x"522f16",x"543118",x"351f0f",x"4c2d16",x"3f2411",x"412612",x"29170a",x"3d2310",x"150e07",x"311c0d",x"311c0c",x"38200f",x"422510",x"351d0d",x"45372c",x"422410",x"3c210f",x"381f0d",x"2d190b",x"361f0f",x"2e1a0c",x"3d2411",x"150e07",x"150e07",x"512f16",x"150e07",x"150e07",x"000000",x"343434",x"323232",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"351f0e",x"351f0e",x"1f1408",x"201408",x"150e07",x"160f07",x"201508",x"2c1a0a",x"2c1a0a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"553b2a",x"553b2a",x"150e07",x"3d210e",x"381f0d",x"402511",x"2c190b",x"371e0d",x"28170a",x"3b2210",x"150e07",x"2b190b",x"2b190b",x"26180f",x"26180f",x"27170d",x"2f1c0f",x"301c0e",x"2d1b0d",x"29170a",x"28170a",x"170f07",x"321c0d",x"554234",x"482c19",x"422919",x"402818",x"442a18",x"442a18",x"2b1a0d",x"2b1a0d",x"000000",x"000000",x"333333",x"333232",x"353433",x"323232",x"333333",x"333232",x"4a4a4a",x"525252",x"424242",x"363636",x"3c3c3c",x"323232",x"383838",x"464646",x"484848",x"5e5e5e",x"565656",x"333333",x"323232",x"4e4e4e",x"323232",x"333333",x"000000",x"000000",x"333333",x"333333",x"343434",x"353535",x"333333",x"323232",x"5c5c5c",x"363636",x"474747",x"353535",x"484541",x"534d48",x"333333",x"3d3d3d",x"3c3c3c",x"343434",x"333333",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"4f4f4f",x"6c6c6c",x"393939",x"353535",x"323131",x"323232",x"323232",x"313131",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452611",x"452611",x"3b200e",x"321a0b",x"301a0b",x"321c0c",x"3a200f",x"422612",x"402511",x"381f0e",x"3d2310",x"321c0d",x"1c1108",x"4c3624",x"463220",x"473320",x"442f1d",x"442f1d",x"432f1d",x"432f1e",x"45311f",x"483320",x"4c3522",x"4e3724",x"4f3824",x"4e3824",x"503823",x"513924",x"513a25",x"503a24",x"513924",x"513924",x"4f3824",x"4e3824",x"503924",x"503a24",x"503a25",x"543d27",x"513a25",x"533c27",x"543d27",x"543c27",x"533b26",x"503a25",x"4a331e",x"4b3520",x"483421",x"473320",x"45301e",x"583e28",x"583e28",x"17110a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463d34",x"463d34",x"3e362e",x"3f342a",x"492f1f",x"361d0b",x"331c0b",x"3b210f",x"351c0c",x"3b210f",x"3b200e",x"3e220f",x"3e2310",x"3e2310",x"381f0d",x"41230f",x"53493f",x"41372d",x"3e2f24",x"4a3120",x"4a3120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"402410",x"402410",x"4a3222",x"403024",x"564c42",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1b0c",x"150e07",x"150e07",x"150e07",x"170f07",x"322116",x"302117",x"3c3229",x"3c3229",x"000000",x"000000",x"524136",x"524136",x"3f210e",x"331c0c",x"341c0c",x"341d0c",x"321b0c",x"321c0c",x"341d0d",x"341d0c",x"331c0c",x"311b0c",x"301b0b",x"2d190a",x"2f190b",x"2c180a",x"2c170a",x"2c170a",x"2c180a",x"2c190b",x"301b0b",x"29170a",x"2e190b",x"2b170a",x"2b1709",x"271509",x"2a160a",x"2c180a",x"2e190b",x"2d190b",x"301b0c",x"331d0d",x"311c0c",x"311b0c",x"2e190b",x"28170a",x"311b0c",x"2d190b",x"29170a",x"2d190b",x"2b180b",x"2b180b",x"2c190b",x"311b0c",x"25150a",x"2e1a0c",x"2d190b",x"25160a",x"27160a",x"29170a",x"2a170a",x"27160a",x"2b180b",x"2b180b",x"29180a",x"29170a",x"2b180b",x"27170a",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"150e07",x"150e07",x"1b1108",x"422816",x"422816",x"2c251e",x"412410",x"412410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d2b14",x"4d2b14",x"3b220f",x"361e0d",x"341d0d",x"3b2210",x"2a180b",x"28170b",x"26160a",x"27170a",x"2a180b",x"29180b",x"2e1a0b",x"40230f",x"343434",x"606060",x"636363",x"333333",x"333333",x"3c3c3c",x"454545",x"454545",x"4d4d4d",x"3e3e3e",x"323232",x"323232",x"393939",x"3b3b3b",x"3a3a3a",x"3d3d3d",x"333333",x"404040",x"5a5a5a",x"4d4d4d",x"484848",x"3f3f3f",x"363636",x"323232",x"323232",x"323232",x"4f4f4f",x"616161",x"333333",x"323232",x"5b5b5b",x"565656",x"333333",x"414141",x"323232",x"343434",x"2c2d2d",x"454545",x"4c4c4c",x"414141",x"464646",x"424242",x"444444",x"4e4e4e",x"525252",x"5c5c5c",x"5c5c5c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1b130b",x"1b130b",x"150e07",x"150e07",x"502e16",x"502e16",x"523017",x"311d0e",x"4a2c16",x"3d2411",x"3f2512",x"29170a",x"37200f",x"2f1b0c",x"25150a",x"2f1a0c",x"311c0d",x"3d210e",x"351e0d",x"4a3c32",x"412411",x"311c0c",x"371f0d",x"3a210f",x"2f1c0d",x"321c0d",x"3e2411",x"22140a",x"150e07",x"553218",x"150e07",x"150e07",x"000000",x"000000",x"313131",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"231509",x"231509",x"150e07",x"150e07",x"181007",x"160f07",x"1d1208",x"2b1a0a",x"2b1a0a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"583e2d",x"583e2d",x"150e07",x"432711",x"331c0c",x"412611",x"3e2411",x"2a180b",x"311b0c",x"371f0e",x"27170a",x"2d1a0c",x"2d1a0c",x"24180f",x"24180f",x"26180e",x"2c1b0e",x"2e1c0d",x"2e1a0d",x"251509",x"1d1108",x"160e07",x"3c220f",x"4f3d30",x"472b19",x"3e2818",x"402818",x"432a18",x"452b19",x"382212",x"382212",x"000000",x"000000",x"000000",x"44403c",x"323232",x"333333",x"333333",x"323232",x"323232",x"4d4d4d",x"333333",x"323232",x"3d3d3d",x"585858",x"5e5d5d",x"646362",x"666666",x"444444",x"323232",x"323232",x"313131",x"323232",x"5a5a5a",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"303030",x"333333",x"333333",x"5e5e5e",x"4c4c4c",x"414141",x"000000",x"000000",x"534d48",x"333333",x"3d3d3d",x"3c3c3c",x"343434",x"333333",x"333333",x"323232",x"333333",x"000000",x"000000",x"000000",x"3c3c3c",x"4a4a4a",x"4f4f4f",x"414141",x"313131",x"323232",x"322f2e",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432510",x"432510",x"331c0d",x"321b0b",x"351d0d",x"2d190b",x"361f0e",x"412611",x"412511",x"39200e",x"3d2310",x"3c210f",x"1f1309",x"5e432d",x"1d140b",x"1d140b",x"1d140b",x"1e140b",x"22170c",x"271a0e",x"271a0d",x"271a0e",x"271b0d",x"261a0e",x"271b0e",x"281b0f",x"2c1d0f",x"2e1f0f",x"2f1f0f",x"2f1f10",x"2d1e0f",x"2b1d0f",x"2c1d0f",x"291b0e",x"281b0e",x"2a1c0f",x"2b1d0f",x"291c0f",x"2a1c0e",x"291b0e",x"2a1c0f",x"271a0d",x"25190c",x"281a0d",x"2b1d0e",x"20160d",x"20160c",x"20160c",x"1d140b",x"79593d",x"79593d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"453c33",x"453c33",x"3e342c",x"3d3229",x"4f3524",x"351a0b",x"361e0d",x"331d0d",x"341c0c",x"3a200e",x"391f0e",x"3c220f",x"402411",x"361d0d",x"3c210e",x"42240f",x"534a41",x"41362d",x"403127",x"4b3120",x"4b3120",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412411",x"412411",x"4a2e1c",x"342519",x"52483f",x"150e07",x"150e07",x"150e07",x"150e07",x"2e1b0d",x"150e07",x"150e07",x"150e07",x"1a1008",x"342115",x"302218",x"3b3129",x"3b3129",x"000000",x"000000",x"534135",x"534135",x"41240f",x"2f190a",x"301b0b",x"341c0c",x"2f1a0b",x"331c0c",x"301b0b",x"321c0c",x"2f1a0b",x"2e190b",x"301a0b",x"2f1a0b",x"301b0b",x"301a0b",x"2f1a0b",x"331c0c",x"321c0c",x"321c0c",x"29170a",x"2a170a",x"2b180a",x"2b180a",x"2e190a",x"2c180a",x"2c180a",x"2e190b",x"2f1a0c",x"321c0c",x"311c0c",x"301b0c",x"321d0d",x"321c0c",x"301b0b",x"301a0b",x"301b0c",x"2c190b",x"2d190b",x"2f1b0c",x"2d190b",x"301c0c",x"321d0d",x"2f1b0c",x"301c0d",x"311c0d",x"26160a",x"27160a",x"201309",x"231409",x"2c190b",x"2f1b0c",x"2c190b",x"29170a",x"221409",x"27160a",x"2d1a0b",x"2d1a0b",x"1d1108",x"1d1108",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"502d15",x"502d15",x"150e07",x"150e07",x"1f1309",x"462a17",x"462a17",x"2c241d",x"40230f",x"40230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"462511",x"462511",x"3b2210",x"3a2210",x"1f1209",x"36200f",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"231509",x"2b170a",x"40230f",x"363535",x"6d6a66",x"6b6866",x"313131",x"313131",x"4b4b4b",x"4b4b4b",x"434343",x"353535",x"323232",x"4a4a4a",x"373737",x"373737",x"3e3e3e",x"3d3d3d",x"434343",x"353535",x"4a4a4a",x"4e4e4e",x"595959",x"000000",x"000000",x"323232",x"333333",x"3f3f3f",x"313131",x"343434",x"464646",x"313131",x"4b4b4b",x"595959",x"323232",x"323232",x"323232",x"333333",x"323232",x"333333",x"313131",x"323232",x"3f3f3f",x"4b4b4b",x"484848",x"484848",x"4b4b4b",x"585858",x"5f5f5f",x"5c5c5c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"170f07",x"513017",x"513017",x"482812",x"331e0e",x"402612",x"3f2512",x"301c0d",x"321c0c",x"150e07",x"24150a",x"150e07",x"1a1008",x"2b190b",x"3a200e",x"3d2210",x"4e4237",x"432611",x"38200e",x"2d190b",x"3c2310",x"150e07",x"150e07",x"2c190c",x"371f0f",x"150e07",x"533117",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"381f0e",x"381f0e",x"150e07",x"160e07",x"150e07",x"180f07",x"201508",x"2d1a0b",x"2d1a0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5d4433",x"5d4433",x"150e07",x"432511",x"351d0d",x"361f0e",x"3e2511",x"150e07",x"201309",x"231409",x"38200f",x"221409",x"221409",x"25180f",x"25180f",x"25180d",x"2a1a0e",x"2b190c",x"2b190d",x"2d1a0b",x"201309",x"160e07",x"3d220f",x"503b2d",x"412919",x"432a19",x"3f2818",x"3e2618",x"3f2716",x"2b1a0e",x"2b1a0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"313131",x"626262",x"323231",x"323232",x"323232",x"333333",x"353433",x"3a3735",x"534d48",x"494746",x"353535",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"343434",x"313131",x"333333",x"414141",x"606060",x"484848",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e3e3e",x"4c4c4c",x"545454",x"616161",x"474747",x"313131",x"555555",x"323232",x"3a3a3a",x"333333",x"333333",x"322f2e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462711",x"462711",x"391f0d",x"351d0c",x"381f0e",x"331d0c",x"331d0d",x"3e220f",x"432712",x"3a200e",x"3f2410",x"3d2210",x"1c1108",x"59402a",x"1d140b",x"20160c",x"20160c",x"23180d",x"2a1d0f",x"2c1d10",x"291c0e",x"281b0e",x"2d1e10",x"2d1e10",x"2c1e11",x"2f2011",x"312212",x"332313",x"312112",x"312112",x"2e1f11",x"312113",x"302213",x"302012",x"2f2112",x"312113",x"312213",x"322314",x"312212",x"322313",x"322212",x"2e2011",x"2e1f11",x"2d1e0f",x"2c1d0f",x"25190e",x"24190e",x"251a0f",x"23180e",x"765639",x"765639",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"473e35",x"473e35",x"3a322a",x"362c24",x"4c3120",x"351c0b",x"361e0d",x"351e0d",x"391f0d",x"3b210f",x"3e2310",x"3e2310",x"39200f",x"391f0d",x"3b200e",x"3d210e",x"4e453b",x"41372d",x"403126",x"4b3221",x"4b3221",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f220f",x"3f220f",x"452815",x"312318",x"473e35",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1a0c",x"150e07",x"150e07",x"150e07",x"1a1008",x"312015",x"2d1f16",x"3f352c",x"3f352c",x"000000",x"000000",x"574132",x"574132",x"422410",x"321b0c",x"321b0b",x"311a0b",x"331c0c",x"311b0b",x"2e190b",x"361e0d",x"301a0b",x"311b0c",x"361e0d",x"311b0c",x"311b0b",x"331c0c",x"321c0c",x"321c0c",x"341d0d",x"321c0c",x"2d190b",x"2b180a",x"2d190b",x"2c180a",x"301a0b",x"2c190b",x"261609",x"27160a",x"301b0c",x"2e190b",x"2d190b",x"2c180a",x"2f1a0b",x"301c0c",x"331d0d",x"2e1a0b",x"2a170a",x"2a170a",x"2a170a",x"2c190b",x"2e1a0c",x"301b0c",x"2d1a0b",x"2d190b",x"311b0c",x"2e1a0b",x"2d190b",x"251509",x"2b180b",x"241509",x"2a180b",x"2f1a0c",x"2b180b",x"231409",x"2b190b",x"25160a",x"29180b",x"2b190b",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2a14",x"4b2a14",x"150e07",x"150e07",x"150e07",x"3c2514",x"3c2514",x"2d261f",x"3f230f",x"3f230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4e2d15",x"4e2d15",x"3c220f",x"3f2511",x"3e2512",x"402512",x"2e1b0c",x"2d1a0c",x"341d0d",x"311c0d",x"1f1309",x"2d1a0c",x"29170a",x"3d200d",x"363534",x"414141",x"5a5a5a",x"323232",x"333333",x"323232",x"434343",x"4b4b4b",x"333333",x"333333",x"323232",x"3c3c3c",x"3f3f3f",x"313131",x"535352",x"373737",x"343434",x"353535",x"454545",x"5f5e5e",x"5c5b5a",x"323232",x"31302f",x"333333",x"414141",x"333333",x"333333",x"373737",x"4d4d4d",x"505050",x"4e4e4e",x"5b5b5a",x"333333",x"000000",x"333333",x"333333",x"333333",x"313131",x"333333",x"323232",x"373737",x"3c3c3c",x"3e3e3e",x"4d4d4d",x"4c4c4c",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"1e1208",x"1e1208",x"472711",x"523017",x"26160a",x"402612",x"432713",x"422612",x"371f0e",x"2f1c0d",x"331d0e",x"341d0d",x"331c0d",x"24150a",x"3b200e",x"371f0e",x"4f4136",x"422410",x"402410",x"371f0e",x"27170b",x"3d2411",x"150e07",x"341d0d",x"3d2311",x"150e07",x"502e16",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f2410",x"3f2410",x"150e07",x"150e07",x"150e07",x"181007",x"1c1208",x"311d0b",x"311d0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"563c2b",x"563c2b",x"150e07",x"3f220f",x"381f0d",x"3a210f",x"2f1b0c",x"351d0d",x"150e07",x"341d0d",x"36200f",x"2e1a0b",x"2e1a0b",x"261910",x"261910",x"25160d",x"2a1a0e",x"28180c",x"27170b",x"2b190b",x"27160a",x"160e07",x"402410",x"4b382b",x"4a2e1b",x"442b19",x"3e2818",x"362216",x"402919",x"342011",x"342011",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"373737",x"626262",x"323232",x"333333",x"323232",x"323232",x"353333",x"3e3a39",x"4c4744",x"383838",x"4b4b4b",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"333333",x"333333",x"343434",x"343434",x"484848",x"333333",x"555555",x"545454",x"000000",x"000000",x"525252",x"454545",x"3b3b3b",x"333333",x"454545",x"494949",x"323232",x"545454",x"616161",x"4d4d4d",x"323232",x"323232",x"4e4e4e",x"454545",x"383838",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462812",x"462812",x"341d0c",x"331c0c",x"3d230f",x"321b0b",x"3c210f",x"2f190b",x"412511",x"3f2310",x"412512",x"402511",x"22150a",x"644a32",x"24190f",x"24190f",x"23180e",x"261a0e",x"2f2011",x"312112",x"352415",x"2b1d0f",x"2d1e0f",x"2e1f11",x"2e2012",x"2c1d10",x"312111",x"352313",x"332313",x"342312",x"302113",x"302113",x"2f2113",x"322313",x"302012",x"2f2011",x"372616",x"332414",x"342415",x"2f2011",x"2f1f11",x"302011",x"302011",x"302010",x"2e2011",x"291d11",x"261b10",x"24190f",x"23180e",x"5c432d",x"5c432d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463d34",x"463d34",x"383028",x"372d25",x"492f1e",x"371d0c",x"3a200e",x"371e0d",x"371e0d",x"371e0d",x"3d220f",x"341d0d",x"351d0d",x"3c210e",x"3c210f",x"3b1e0d",x"4a4138",x"40362e",x"44362b",x"4b3526",x"4b3526",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f220f",x"3f220f",x"412716",x"322116",x"473e36",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1b0c",x"150e07",x"150e07",x"150e07",x"190f07",x"322015",x"2b2017",x"42372e",x"42372e",x"000000",x"000000",x"4e3e33",x"4e3e33",x"3e220f",x"351d0d",x"38200e",x"361f0e",x"3a210f",x"371f0e",x"39200e",x"361f0e",x"361f0e",x"351d0d",x"2f1a0b",x"2a180a",x"321b0b",x"311b0b",x"2e190b",x"2f1a0b",x"2f190b",x"2d180a",x"2e190b",x"2b170a",x"28160a",x"2b180a",x"2c190a",x"2f1a0b",x"26160a",x"231409",x"29170a",x"2e190b",x"2e190b",x"311b0c",x"321d0d",x"311c0d",x"29170a",x"2c180a",x"2c180b",x"2e1a0b",x"2c180b",x"29170a",x"331d0d",x"311d0d",x"301c0d",x"311c0c",x"331d0d",x"2c190b",x"2c190b",x"2d1a0b",x"2c190b",x"311c0c",x"2d1a0b",x"2b180b",x"2e1a0c",x"2e1a0b",x"2a180b",x"2a180b",x"211409",x"27160a",x"190f08",x"190f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452510",x"452510",x"150e07",x"150e07",x"221409",x"432816",x"432816",x"382e26",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"522f16",x"522f16",x"39210f",x"3f2511",x"402512",x"38200f",x"38200f",x"39200e",x"2b190b",x"2d1a0c",x"150e07",x"201309",x"271609",x"3f220e",x"333232",x"454545",x"5e5e5e",x"3d3d3d",x"525252",x"333333",x"343434",x"313131",x"555555",x"525252",x"373737",x"373737",x"5b5b5b",x"515151",x"565656",x"333333",x"323232",x"373737",x"4e4e4e",x"64605d",x"64605d",x"333333",x"323232",x"585858",x"545454",x"363636",x"535353",x"515151",x"343434",x"515151",x"5f5f5f",x"616160",x"616160",x"000000",x"000000",x"000000",x"000000",x"000000",x"353535",x"323232",x"373737",x"3c3c3c",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"25160a",x"28170a",x"512f16",x"4d2c14",x"2d1a0c",x"3e2411",x"422712",x"432713",x"321c0d",x"3d2411",x"3a2110",x"2a170a",x"361e0d",x"150e07",x"3f2410",x"3c2310",x"54453a",x"462712",x"3f2411",x"3b220f",x"331e0e",x"432713",x"1c1108",x"361e0d",x"3e2411",x"150e07",x"4e2d15",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"3d230f",x"29170a",x"371f0e",x"351e0d",x"150e07",x"331d0c",x"422611",x"422611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533928",x"533928",x"150e07",x"3c200e",x"3a200e",x"3d230f",x"311c0c",x"361e0d",x"150e07",x"351e0e",x"3c2310",x"2d1a0c",x"2d1a0c",x"25180f",x"25180f",x"25160d",x"2a1a0f",x"28170c",x"25160b",x"27170a",x"241509",x"150e07",x"3f2410",x"4a372b",x"4a2e1b",x"422a1a",x"3f2819",x"3b2516",x"422a18",x"352011",x"352011",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"353333",x"3e3a39",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"393939",x"333333",x"313131",x"4e4e4e",x"414141",x"5f5f5f",x"4f4f4f",x"4d4d4d",x"525252",x"454545",x"3b3b3b",x"333333",x"333333",x"313131",x"303030",x"333333",x"3f3d3b",x"5f5f5f",x"313131",x"323232",x"2d2925",x"525252",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432511",x"432511",x"351c0c",x"321b0b",x"3b220f",x"321b0b",x"3a210f",x"371d0c",x"3c2210",x"3a210e",x"3e2410",x"3e2411",x"1b1108",x"6b5037",x"251a0f",x"25190f",x"251a0f",x"2d1f11",x"2b1d0f",x"372412",x"2c1e10",x"302113",x"312212",x"2f2011",x"332314",x"342314",x"352414",x"372516",x"2f1f12",x"312112",x"2d1f12",x"2d1f12",x"2e1f11",x"2e1f12",x"302112",x"322213",x"332314",x"322313",x"312113",x"332212",x"342313",x"332315",x"342314",x"312213",x"2f2114",x"2b1f13",x"281c11",x"25190f",x"22170e",x"644931",x"644931",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463d34",x"463d34",x"372f27",x"342b22",x"452a19",x"381e0c",x"3a200e",x"351c0c",x"3b210e",x"3c210f",x"361e0d",x"3a200e",x"3a210e",x"3e2310",x"3d220f",x"291307",x"54493f",x"4b4137",x"4a3d32",x"493326",x"493326",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"432816",x"352417",x"473d33",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1a0c",x"150e07",x"150e07",x"150e07",x"170f07",x"332216",x"362519",x"3f352c",x"3f352c",x"000000",x"000000",x"46372b",x"46372b",x"422511",x"301a0c",x"39210f",x"341e0d",x"361f0e",x"331c0c",x"150e07",x"3a200e",x"341c0c",x"361e0d",x"331d0d",x"321b0b",x"381f0e",x"3a210f",x"361e0d",x"341d0c",x"2f1a0b",x"321b0b",x"301a0b",x"2f1a0b",x"27160a",x"2e1a0b",x"311b0c",x"27160a",x"2b180b",x"27160a",x"2c180a",x"2d190a",x"2b180a",x"2a160a",x"271509",x"281609",x"28160a",x"2d190b",x"2f1a0b",x"301b0c",x"2e1a0b",x"2c180b",x"2b180b",x"2f1b0c",x"2f1a0b",x"2e1a0b",x"2e1b0c",x"27170a",x"27170a",x"2e1b0c",x"2a190b",x"2a180b",x"2d1a0b",x"2a170b",x"201208",x"231409",x"1d1108",x"221409",x"231409",x"241509",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341909",x"341909",x"150e07",x"150e07",x"1f1209",x"442916",x"442916",x"352d25",x"40230f",x"40230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4f2e15",x"4f2e15",x"3b2210",x"422612",x"3c2310",x"150e07",x"341e0d",x"150e07",x"2a180b",x"311b0c",x"1d1208",x"26170a",x"221309",x"3e220e",x"323232",x"333333",x"343434",x"5a5a5a",x"6a6a6a",x"5d5d5d",x"565656",x"444444",x"4b4b4b",x"555555",x"575757",x"5e5e5e",x"5a5a5a",x"535353",x"565656",x"313131",x"333333",x"3d3d3d",x"595959",x"5e5e5d",x"4c4c4c",x"373737",x"323232",x"313131",x"4f4f4f",x"555555",x"4c4c4c",x"5d5d5d",x"333333",x"393939",x"585858",x"656564",x"656564",x"3a3a3a",x"3b3b3b",x"323232",x"333333",x"363636",x"353535",x"323232",x"323232",x"3d3d3d",x"3b3b3b",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"1d1109",x"201308",x"472712",x"4e2d15",x"2d1a0d",x"3f2411",x"3f2512",x"3d2310",x"150e07",x"36200f",x"382110",x"2a180b",x"341d0c",x"150e07",x"412611",x"382210",x"544236",x"462611",x"381f0e",x"3b2210",x"3d2310",x"3f2411",x"150e07",x"381f0e",x"452814",x"150e07",x"4b2c15",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d230f",x"29170a",x"1e1308",x"221508",x"150e07",x"331d0c",x"422611",x"422611",x"000000",x"000000",x"000000",x"343434",x"343434",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503726",x"503726",x"150e07",x"3d210e",x"3a200e",x"3b200e",x"3f2410",x"351d0d",x"150e07",x"38200f",x"3b220f",x"231409",x"231409",x"26190f",x"26190f",x"24160d",x"2a1a0e",x"2c1a0e",x"29180c",x"2b190b",x"27160a",x"150e07",x"3e2310",x"4c382c",x"4b2f1d",x"402919",x"3e2718",x"392416",x"3e2818",x"28190d",x"28190d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"393939",x"5c5c5c",x"323232",x"323232",x"333333",x"323232",x"606060",x"4f4f4f",x"4a4a4a",x"3e3e3e",x"313131",x"353535",x"313131",x"323232",x"333333",x"323232",x"343434",x"5c5a59",x"5d5c5c",x"353535",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2d15",x"4f2d15",x"361e0d",x"39200e",x"3e230f",x"341c0c",x"3c210f",x"351e0d",x"442712",x"3c220f",x"422612",x"422612",x"1e1208",x"6c4f36",x"25190f",x"21170d",x"261a0f",x"2c1e0f",x"2d1e0f",x"2b1d0f",x"2e1f11",x"2d1f11",x"322312",x"312212",x"322112",x"332212",x"342212",x"352412",x"2f1f11",x"302012",x"2a1d10",x"2b1d11",x"2f2113",x"2c1e10",x"2e1f11",x"312112",x"302113",x"2e1f11",x"2c1e11",x"302112",x"322112",x"322212",x"312112",x"312111",x"2c1f11",x"271c11",x"271b10",x"261b0f",x"21160d",x"493422",x"493422",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"443a31",x"443a31",x"322a22",x"352a22",x"492d1d",x"321b0b",x"381f0e",x"331c0c",x"3b210e",x"381f0e",x"3b210f",x"3b210f",x"3d2310",x"3a210e",x"3c210e",x"271106",x"584e43",x"4b4036",x"483b32",x"493326",x"493326",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200e",x"38200e",x"412616",x"342216",x"483f36",x"150e07",x"150e07",x"150e07",x"150e07",x"2a190b",x"150e07",x"150e07",x"150e07",x"170f07",x"312015",x"34251b",x"42372e",x"42372e",x"000000",x"000000",x"47362a",x"47362a",x"4b2b14",x"351d0d",x"351e0e",x"331d0d",x"331d0d",x"39210f",x"150e07",x"2f1a0b",x"3a200d",x"381f0d",x"331c0c",x"321c0c",x"351d0d",x"3a210f",x"361f0e",x"361f0d",x"341d0d",x"331c0c",x"321c0c",x"2d190b",x"29170a",x"2c180b",x"2f1a0b",x"2c180b",x"2a170a",x"2f1a0b",x"301b0b",x"2f1a0b",x"2d190b",x"2d190b",x"2b180b",x"2c190b",x"2b170a",x"2f1a0b",x"2d1a0b",x"2e1a0c",x"2b180a",x"2a170a",x"2d1a0b",x"311c0d",x"2e1b0c",x"2b180b",x"2c190b",x"331d0d",x"341e0d",x"2b180b",x"2c190b",x"2d190b",x"2f1b0c",x"251509",x"1f1208",x"1f1108",x"1c1008",x"1e1209",x"211309",x"231409",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"34190a",x"34190a",x"150e07",x"150e07",x"1b1108",x"472b18",x"472b18",x"342c25",x"41230f",x"41230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"3d2410",x"2c190b",x"38200e",x"150e07",x"38200e",x"150e07",x"311c0c",x"150e07",x"341e0e",x"321d0d",x"2c180b",x"452611",x"535353",x"535353",x"545454",x"575757",x"515151",x"464646",x"353535",x"313131",x"444444",x"494949",x"575757",x"666565",x"545454",x"545454",x"3c3c3c",x"383838",x"323232",x"383838",x"3e3e3e",x"595959",x"4c4c4c",x"414141",x"3c3c3c",x"373737",x"333333",x"333333",x"3f3f3f",x"565656",x"323232",x"393939",x"464646",x"333333",x"363636",x"3a3a3a",x"3b3b3b",x"323232",x"333333",x"4f4f4f",x"434343",x"343434",x"353535",x"3d3d3d",x"3b3b3b",x"323232",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"2b180b",x"432510",x"4c2d15",x"341f0e",x"3f2411",x"321d0e",x"3c2210",x"150e07",x"361f0e",x"38200f",x"2e1b0c",x"150e07",x"301c0c",x"452712",x"361f0f",x"4c3b2f",x"432510",x"3a200f",x"371f0e",x"3b2210",x"432813",x"150e07",x"38200e",x"412612",x"150e07",x"4f2d16",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"281809",x"261809",x"1e1308",x"221508",x"241708",x"201508",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"343434",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513827",x"513827",x"150e07",x"3a1f0d",x"39200e",x"3c2310",x"3a210f",x"361d0d",x"150e07",x"311b0c",x"39210f",x"2d1a0c",x"2d1a0c",x"25180e",x"25180e",x"26170d",x"2a1a0e",x"2a180c",x"27180c",x"29170b",x"2a180b",x"150e07",x"3e2410",x"4b382d",x"472d1b",x"432a19",x"3e2818",x"3f2617",x"3f2719",x"321e10",x"321e10",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"4d4d4d",x"595959",x"3f3d3b",x"555555",x"4b4b4b",x"383838",x"303030",x"333333",x"333333",x"32302f",x"323232",x"323232",x"353535",x"383432",x"51504f",x"4a4a4a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2b14",x"4c2b14",x"412511",x"3a200e",x"3d220f",x"341c0c",x"3f2310",x"3f2410",x"402511",x"3d220f",x"3f2411",x"432713",x"1d1208",x"6a4d35",x"261a0f",x"23180e",x"271b0e",x"2b1e10",x"2d1e0f",x"2c1e0f",x"2d1e10",x"302011",x"2e1f11",x"352312",x"2c1d0f",x"2e1f0f",x"2b1c0f",x"2c1e10",x"2f2112",x"302213",x"2d1f12",x"2d1f12",x"312215",x"312112",x"2e2013",x"2e2012",x"2f2012",x"302113",x"302113",x"312113",x"332213",x"312212",x"312111",x"2f1f11",x"2b1d0f",x"261a0f",x"23180e",x"23180e",x"21170d",x"59412b",x"59412b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"463d35",x"463d35",x"3b322a",x"362c25",x"472e20",x"381e0d",x"3a200e",x"331c0c",x"381f0e",x"361e0d",x"402511",x"3f2410",x"3f2410",x"3f2410",x"3d220f",x"2a1206",x"544a40",x"4a4036",x"473a30",x"4f382a",x"4f382a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452712",x"452712",x"442918",x"37271b",x"453c34",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1b0c",x"150e07",x"150e07",x"150e07",x"191008",x"2f1f15",x"35261c",x"453a31",x"453a31",x"000000",x"000000",x"4f3e32",x"4f3e32",x"472712",x"331d0d",x"38200f",x"331d0d",x"38200f",x"37200f",x"150e07",x"351d0b",x"371e0d",x"331c0c",x"351d0c",x"351d0d",x"371e0d",x"371f0e",x"351e0d",x"371f0e",x"361e0e",x"361f0e",x"341d0d",x"351e0d",x"311b0c",x"331c0c",x"2d190b",x"331c0c",x"2e1a0b",x"2c180a",x"301a0b",x"2c180a",x"2b180a",x"2b180a",x"2a170a",x"2c180a",x"2a180a",x"28160a",x"2d190b",x"241509",x"2a170a",x"2b180b",x"29180b",x"2f1b0c",x"301c0d",x"311d0d",x"2f1c0d",x"2d1a0c",x"2f1b0c",x"2b190b",x"2a180b",x"301b0c",x"2a180b",x"251509",x"201108",x"1d1108",x"1c1108",x"221409",x"29180b",x"1f1208",x"160f07",x"160f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462711",x"462711",x"150e07",x"150e07",x"201309",x"4b2e19",x"4b2e19",x"3d2f25",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4b2913",x"4b2913",x"3e230f",x"3c220f",x"331d0d",x"2f1b0c",x"39200e",x"150e07",x"1d1208",x"2e1a0b",x"3b2210",x"2c1a0b",x"2c180b",x"4b2a13",x"4e4e4e",x"616161",x"4d4d4d",x"323232",x"3e3e3e",x"4d4d4d",x"393939",x"303030",x"323232",x"3c3c3c",x"5b5b5b",x"666565",x"545454",x"555555",x"4e4e4e",x"343434",x"5e5e5e",x"464646",x"5c5c5c",x"5d5d5d",x"414141",x"383838",x"4a4a4a",x"505050",x"5e5e5e",x"525252",x"323232",x"313131",x"323232",x"545454",x"4b4b4b",x"3b3b3b",x"333333",x"4b4b4b",x"696969",x"686868",x"535353",x"525252",x"545454",x"525252",x"3d3d3d",x"5b5b5b",x"5e5e5e",x"454545",x"333333",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"361e0d",x"462610",x"502e15",x"2b190b",x"442713",x"402512",x"351e0e",x"2d1a0b",x"361e0d",x"2a180b",x"2e1b0d",x"2e190b",x"351d0c",x"472813",x"361f0e",x"4c3b2f",x"432510",x"3e2310",x"331c0c",x"341e0e",x"3f2511",x"150e07",x"371f0e",x"402512",x"150e07",x"502f16",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2f1c09",x"2f1c09",x"201508",x"241708",x"211508",x"211508",x"000000",x"000000",x"000000",x"000000",x"000000",x"343434",x"323232",x"333333",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503829",x"503829",x"150e07",x"3f230f",x"3a200e",x"3f2511",x"2d1a0c",x"341d0c",x"150e07",x"2b180a",x"341d0d",x"2a180b",x"2a180b",x"24170d",x"24170d",x"27190e",x"2a190e",x"29180c",x"2a180c",x"28170a",x"1c1108",x"150e07",x"3c2210",x"513b2e",x"492e1c",x"3e2719",x"3b2618",x"3b2517",x"432a18",x"26170c",x"26170c",x"40220f",x"4d2c15",x"462812",x"42230f",x"452712",x"4b2a14",x"4b2b15",x"482913",x"452611",x"432511",x"4a2a14",x"4d2d15",x"482913",x"482913",x"472812",x"472913",x"452712",x"422410",x"432510",x"452711",x"452711",x"432510",x"412410",x"472711",x"3f220f",x"412310",x"412410",x"422410",x"3e220f",x"432511",x"422511",x"402410",x"3f230f",x"3b210f",x"412411",x"565656",x"616161",x"312e2d",x"545454",x"4a4a4a",x"383838",x"323232",x"323232",x"333333",x"462711",x"432511",x"422611",x"452711",x"442611",x"492812",x"432611",x"452611",x"452711",x"462812",x"472913",x"492a14",x"4a2a14",x"492a13",x"432611",x"442611",x"422510",x"3f230f",x"41230f",x"412410",x"3f230f",x"432611",x"3e230f",x"402411",x"3f2310",x"432612",x"4b2a13",x"4b2a13",x"3c210f",x"3d220f",x"3d220f",x"331c0c",x"3f2410",x"402411",x"3e2310",x"3d2310",x"432511",x"432612",x"1d1208",x"61462e",x"23180e",x"20160d",x"281b0d",x"2e1f10",x"281a0d",x"2a1c0e",x"2d1f10",x"302011",x"312112",x"342312",x"312212",x"302011",x"302113",x"2f2112",x"322315",x"2f2114",x"302113",x"2b1f12",x"2f2113",x"2f2012",x"2e2012",x"2c1e11",x"302011",x"302111",x"2d1f10",x"302111",x"342312",x"322212",x"322212",x"312212",x"332312",x"261a0e",x"23180e",x"20160d",x"20160c",x"4c3724",x"4c3724",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"413931",x"413931",x"382f27",x"332b23",x"462f21",x"361d0c",x"351e0d",x"311b0c",x"3b220f",x"3a1f0d",x"462914",x"3e2410",x"412511",x"412511",x"3d220f",x"3c1f0d",x"564c42",x"494036",x"45382d",x"513726",x"513726",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432611",x"432611",x"432818",x"38291f",x"453c34",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"170f07",x"2e1f15",x"36271c",x"433a31",x"433a31",x"000000",x"000000",x"44352a",x"44352a",x"472812",x"38200f",x"351e0e",x"361f0e",x"351e0e",x"351e0d",x"150e07",x"321c0b",x"341c0c",x"301b0b",x"361e0c",x"311c0c",x"361e0e",x"341d0d",x"321c0c",x"341d0c",x"331c0c",x"341d0c",x"301b0c",x"2e190b",x"311b0c",x"2e190b",x"2d190b",x"2e190b",x"301b0b",x"2e1a0b",x"2e190b",x"2d190b",x"301a0b",x"2b170a",x"271509",x"281609",x"2a170a",x"29170a",x"29160a",x"281609",x"261509",x"28160a",x"2a170a",x"2b180b",x"26160a",x"271609",x"29170a",x"271609",x"251509",x"231409",x"251409",x"1a1007",x"211208",x"221409",x"1f1108",x"1f1208",x"180f07",x"180f07",x"25160a",x"221409",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"442611",x"442611",x"150e07",x"150e07",x"25160a",x"3b2414",x"3b2414",x"322b24",x"412410",x"412410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482812",x"482812",x"3f2310",x"3c230f",x"38200e",x"2f1b0c",x"3a210f",x"150e07",x"2e1a0c",x"311b0c",x"3a210f",x"29180b",x"2d190b",x"4d2b14",x"4f4f4f",x"505050",x"323232",x"333333",x"413f3c",x"4c4c4c",x"454545",x"333333",x"333333",x"3c3c3c",x"343434",x"666666",x"343434",x"4e4e4e",x"505050",x"323232",x"555555",x"5a5a5a",x"3e3e3e",x"333333",x"393939",x"383838",x"363636",x"373737",x"393939",x"353535",x"676767",x"313131",x"333333",x"585858",x"595959",x"686868",x"646464",x"5b5b5b",x"5c5c5c",x"636363",x"636363",x"565656",x"4e4f4f",x"515151",x"4c4c4c",x"4a4a4a",x"4e4e4e",x"505050",x"575655",x"393939",x"3f3f3f",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"351d0d",x"4f2d15",x"311c0c",x"422611",x"3f2411",x"39200f",x"311c0d",x"371f0e",x"341e0d",x"2e1a0c",x"311b0c",x"2f1a0b",x"472913",x"39210f",x"4a3729",x"452611",x"3f2310",x"351e0d",x"311d0d",x"38200e",x"150e07",x"301c0c",x"38200f",x"150e07",x"4b2b14",x"150e07",x"150e07",x"000000",x"000000",x"655445",x"54463a",x"483c30",x"544132",x"493e34",x"584e44",x"584e43",x"655346",x"574d43",x"584e43",x"5e5146",x"5e5146",x"000000",x"2d1a09",x"261809",x"261809",x"271909",x"2a1a0a",x"261809",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"513d2f",x"513d2f",x"150e07",x"3f230f",x"371e0d",x"3c2310",x"211409",x"301a0b",x"150e07",x"241509",x"331d0d",x"25160a",x"25160a",x"24170d",x"24170d",x"28190e",x"2b1a0f",x"29190c",x"2b190c",x"2a170a",x"1d1108",x"150e07",x"3a210f",x"4e3b2e",x"4a2d1a",x"3d2618",x"3f2918",x"3d2718",x"3f2717",x"362111",x"43250f",x"40220f",x"4d2c15",x"462812",x"42230f",x"452712",x"4b2a14",x"4b2b15",x"482913",x"452611",x"432511",x"4a2a14",x"4d2d15",x"482913",x"482913",x"472812",x"472913",x"452712",x"422410",x"432510",x"452711",x"452711",x"432510",x"412410",x"472711",x"3f220f",x"412310",x"412410",x"422410",x"3e220f",x"432511",x"422511",x"402410",x"3f230f",x"3b210f",x"412411",x"422611",x"3e2310",x"442712",x"3f2310",x"442712",x"472813",x"462813",x"442711",x"442711",x"462711",x"432511",x"422611",x"452711",x"442611",x"492812",x"432611",x"452611",x"452711",x"462812",x"472913",x"492a14",x"4a2a14",x"492a13",x"432611",x"442611",x"422510",x"3f230f",x"41230f",x"412410",x"3f230f",x"432611",x"3e230f",x"402411",x"3f2310",x"432612",x"422512",x"492813",x"3a200e",x"3a200e",x"3a200e",x"381f0d",x"39200e",x"3f2411",x"3b220f",x"3e2310",x"3c220f",x"412511",x"1e1208",x"6b4f36",x"22180d",x"22170d",x"2a1d0f",x"2f2011",x"2f1f0f",x"2d2011",x"291c0f",x"332313",x"332312",x"362514",x"332212",x"2f2012",x"302011",x"2f2011",x"2f2012",x"2e2013",x"2f2012",x"2c1e11",x"2c1f11",x"2b1d11",x"312213",x"322314",x"332314",x"322214",x"312113",x"312212",x"312111",x"362515",x"312112",x"322111",x"2e1f10",x"271a0f",x"22170d",x"22170d",x"22180e",x"4b3724",x"4b3724",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d362d",x"3d362d",x"352d26",x"342c24",x"452d1e",x"371d0c",x"361e0d",x"301a0b",x"371e0d",x"371e0d",x"3a1f0e",x"432712",x"3f2310",x"3c220f",x"3e220f",x"3c200d",x"554b41",x"473d33",x"41352b",x"513523",x"513523",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422510",x"422510",x"432a1c",x"38291f",x"483e35",x"150e07",x"150e07",x"150e07",x"150e07",x"2c190b",x"150e07",x"150e07",x"150e07",x"150e07",x"332115",x"33251a",x"443a31",x"443a31",x"000000",x"000000",x"4d392b",x"4d392b",x"4a2912",x"3e2411",x"351e0d",x"341d0d",x"37200e",x"38200e",x"150e07",x"311b0b",x"311b0b",x"321b0b",x"2d190a",x"321c0c",x"351d0d",x"331c0c",x"311c0c",x"301b0b",x"341d0d",x"361e0d",x"341d0c",x"321c0c",x"2e1a0b",x"2c190a",x"311b0c",x"2f1a0b",x"2f1a0b",x"301a0b",x"2f1a0b",x"2d190b",x"311c0c",x"301b0c",x"331d0d",x"331d0e",x"341e0e",x"2e1a0c",x"2f1b0c",x"2f1b0c",x"28170a",x"2f1b0c",x"2e1a0c",x"301b0c",x"2a180b",x"2c190b",x"29170a",x"29170a",x"28160a",x"271609",x"261509",x"211308",x"261509",x"251509",x"1e1108",x"201208",x"201208",x"221509",x"24150a",x"1f1209",x"190f08",x"190f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2d15",x"4c2d15",x"150e07",x"150e07",x"1f1309",x"432714",x"432714",x"3a2e25",x"3e2310",x"3e2310",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"432510",x"432510",x"3a210f",x"371f0e",x"3c2310",x"27170b",x"3d2310",x"150e07",x"27160a",x"351e0d",x"38200f",x"2d1a0b",x"311a0b",x"502d15",x"5e5e5e",x"2f2f2f",x"3a3a3a",x"4e4d4c",x"4e4d4c",x"595959",x"4c4c4c",x"4e4e4e",x"626262",x"616161",x"464646",x"4f4f4f",x"464646",x"434343",x"454545",x"505050",x"545454",x"393939",x"363636",x"323232",x"333333",x"000000",x"000000",x"3b3b3b",x"333333",x"393938",x"4c4c4c",x"494949",x"2f3030",x"515151",x"525252",x"343434",x"323232",x"323232",x"353535",x"313132",x"313131",x"4f4f4f",x"616161",x"5b5b5b",x"515151",x"505050",x"565656",x"4e4e4d",x"3c3c3c",x"535353",x"4d4d4d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"331c0b",x"4d2d15",x"311c0d",x"412411",x"3f2411",x"3c230f",x"2c1a0c",x"38200e",x"2f1b0c",x"2c1a0c",x"311b0c",x"301a0b",x"432712",x"3b210f",x"4c382a",x"412410",x"39200f",x"3a210f",x"1b1108",x"331c0d",x"150e07",x"2e1a0c",x"2f1b0c",x"150e07",x"4b2a13",x"150e07",x"150e07",x"000000",x"655445",x"655445",x"54463a",x"483c30",x"544132",x"493e34",x"584e44",x"584e43",x"655346",x"574d43",x"584e43",x"5e5146",x"5e5146",x"000000",x"271909",x"2a1b09",x"2b1b09",x"271909",x"38220d",x"38220d",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"333333",x"323232",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"574335",x"574335",x"150e07",x"3d210f",x"341d0c",x"402511",x"150e07",x"301a0b",x"150e07",x"2f1a0b",x"28170b",x"2f1c0d",x"2f1c0d",x"25180e",x"25180e",x"29190e",x"2c1a0e",x"2d1b0d",x"2d190d",x"28170a",x"201208",x"160e07",x"3b200e",x"533e31",x"4a2e1b",x"442a19",x"412919",x"402717",x"3e2616",x"2a190d",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1b120a",x"1f160f",x"221911",x"241b13",x"221810",x"21170f",x"23170f",x"3f2410",x"3f2410",x"361e0d",x"3e230f",x"321b0c",x"39200e",x"3d2310",x"3e2310",x"381f0e",x"361f0d",x"432712",x"1a1008",x"674b33",x"21160d",x"21170d",x"271a0d",x"291c0e",x"2d1d0e",x"2b1d0f",x"342212",x"322110",x"322211",x"352413",x"332314",x"2d1e10",x"332313",x"322213",x"2c1f12",x"312214",x"2e2011",x"2a1d10",x"2f2013",x"2c1e11",x"2d1f11",x"2f2011",x"2d1f11",x"2e1f10",x"2a1c0f",x"2a1c0f",x"2c1e0f",x"2e1e0f",x"2f1f0e",x"2e1f0e",x"2c1d0e",x"271a0d",x"25190e",x"21170d",x"20160d",x"4c3724",x"4c3724",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"423a31",x"423a31",x"373028",x"332b23",x"473022",x"371e0c",x"321b0b",x"331c0c",x"412511",x"351c0c",x"3d2210",x"472a14",x"412511",x"402410",x"402410",x"3e210e",x"564c41",x"50473e",x"493b31",x"563926",x"563926",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422510",x"422510",x"503323",x"3c2c20",x"484037",x"150e07",x"150e07",x"150e07",x"150e07",x"28170b",x"150e07",x"150e07",x"150e07",x"1a1008",x"2f1f15",x"35251a",x"41362d",x"41362d",x"000000",x"000000",x"49372b",x"49372b",x"482812",x"3c2311",x"341d0d",x"331d0d",x"341d0d",x"371f0e",x"150e07",x"351d0c",x"321c0b",x"311c0b",x"311c0c",x"361f0e",x"331c0c",x"371f0d",x"351d0d",x"331d0d",x"371e0d",x"341d0d",x"371f0e",x"321c0c",x"2e1a0b",x"2d190b",x"351d0d",x"301b0b",x"321c0c",x"29160a",x"301b0c",x"311c0c",x"301b0c",x"331c0c",x"2e1a0b",x"2e1a0b",x"2f1a0b",x"301b0c",x"2d190b",x"2c190b",x"2b180b",x"2c190b",x"2f1a0b",x"2d190b",x"2d190b",x"321d0d",x"2e1b0c",x"2e1b0c",x"301b0c",x"2a180b",x"27160a",x"251509",x"2e1a0c",x"251509",x"1d1008",x"1d1108",x"241409",x"221409",x"27170a",x"221409",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2e16",x"4f2e16",x"150e07",x"150e07",x"1c1108",x"442916",x"442916",x"332b23",x"3f230f",x"3f230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"462611",x"462611",x"3d2410",x"3a210f",x"351e0e",x"402512",x"3e2411",x"361e0d",x"1a1108",x"2b190b",x"371f0d",x"2b180b",x"2d180a",x"522f15",x"5f5f5e",x"2c2c2d",x"343434",x"575656",x"575656",x"4e4e4e",x"464646",x"323232",x"303030",x"353535",x"4b4b4b",x"484848",x"3e3e3e",x"333333",x"303030",x"383838",x"414141",x"535353",x"323232",x"323232",x"323232",x"5b5b5b",x"4e4e4e",x"3b3b3b",x"333333",x"363534",x"4e4e4e",x"555555",x"424242",x"535353",x"373737",x"323232",x"323232",x"323232",x"353535",x"313131",x"333333",x"3c3c3c",x"494949",x"424242",x"413f3e",x"4b4b4b",x"484848",x"3b3b3b",x"3b3b3b",x"4d4d4d",x"575757",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"361d0d",x"4c2a14",x"36200f",x"3f2310",x"381f0e",x"361f0e",x"3b2210",x"422612",x"39200f",x"150e07",x"2b180b",x"311b0c",x"432611",x"371f0e",x"4f3d31",x"3e220f",x"311c0d",x"38200e",x"150e07",x"341d0d",x"150e07",x"301a0c",x"1b1108",x"150e07",x"452611",x"150e07",x"150e07",x"000000",x"5a4d41",x"5a4d41",x"5e5145",x"5a4d40",x"6a5342",x"584d43",x"584e44",x"584e43",x"635245",x"584e43",x"54493f",x"5b4e43",x"5b4e43",x"000000",x"281909",x"281909",x"281909",x"2a1a09",x"2f1d0a",x"3a230d",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"404040",x"474747",x"474747",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f3b2e",x"4f3b2e",x"150e07",x"412410",x"2e1a0b",x"3e2310",x"150e07",x"321b0c",x"150e07",x"38200e",x"1b1108",x"24150a",x"24150a",x"27170d",x"27170d",x"2a1a0e",x"2f1d0f",x"2f1c0d",x"2e1a0d",x"2a180b",x"241409",x"170f07",x"351d0c",x"503d30",x"492d1a",x"412918",x"412817",x"3f2717",x"382315",x"2a190d",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"1a1109",x"1f160f",x"241b13",x"251c14",x"271d15",x"251c14",x"251c14",x"231911",x"4d2b13",x"3d220f",x"3b210e",x"3c220f",x"351e0c",x"3b200e",x"3f2411",x"3d220f",x"381f0d",x"3c210f",x"442712",x"211409",x"674b32",x"20160c",x"23180d",x"271a0d",x"2c1d10",x"2d1e10",x"302011",x"332313",x"342311",x"2f2111",x"302011",x"2f2011",x"2d1e10",x"2d1e10",x"2d1f11",x"2c1d10",x"2f1f11",x"2e1e11",x"281b0e",x"2b1d10",x"2b1d10",x"2e1f11",x"291c10",x"2b1d10",x"2c1d10",x"2d1e11",x"291c0f",x"2b1d0f",x"2d1e0f",x"2e1f0f",x"2d1d0e",x"291c0f",x"281b0e",x"25190c",x"23180d",x"1e150c",x"4b3624",x"4b3624",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"433a31",x"433a31",x"3a322a",x"3b322a",x"4a3324",x"3e230f",x"321b0b",x"351d0c",x"3e2310",x"391f0e",x"432612",x"422612",x"3b210f",x"3e2410",x"3e230f",x"40230e",x"594f45",x"584d43",x"584b40",x"594335",x"594335",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"432712",x"432712",x"493023",x"3c2c20",x"4a4137",x"150e07",x"150e07",x"150e07",x"150e07",x"2b190b",x"150e07",x"150e07",x"150e07",x"190f07",x"2b1d13",x"2f2017",x"393028",x"393028",x"000000",x"000000",x"4a372a",x"4a372a",x"4b2c15",x"2f1c0d",x"341d0d",x"361f0e",x"301a0b",x"311b0c",x"150e07",x"311b0c",x"321c0c",x"321c0c",x"2d190b",x"371f0e",x"351d0c",x"351d0d",x"331c0c",x"321c0c",x"321c0c",x"311c0c",x"311c0c",x"311b0c",x"311c0c",x"2c190b",x"331c0c",x"331d0d",x"361e0d",x"351e0d",x"2f1a0b",x"2b180a",x"2a180b",x"2f1a0b",x"301b0c",x"2a180a",x"311b0c",x"301b0c",x"2f1a0b",x"28160a",x"2b180a",x"2d190b",x"2a170a",x"251509",x"261509",x"271609",x"2b180a",x"28160a",x"29170a",x"2c190b",x"29170a",x"2b180b",x"2a180a",x"1f1208",x"1e1108",x"1f1108",x"201308",x"241509",x"25160a",x"191008",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2d16",x"4f2d16",x"150e07",x"150e07",x"1f1209",x"4a2c17",x"4a2c17",x"362c23",x"432611",x"432611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482811",x"482811",x"3d2310",x"3c2311",x"150e07",x"3d2310",x"2c1a0b",x"331d0d",x"150e07",x"150e07",x"351e0d",x"2f1a0b",x"2f190b",x"512e16",x"5a5a5a",x"545454",x"323232",x"333333",x"595959",x"515151",x"353535",x"383838",x"383838",x"4e4e4e",x"4e4e4e",x"383838",x"383838",x"414141",x"545454",x"323232",x"393938",x"515151",x"555555",x"313131",x"323232",x"616161",x"5b5b5b",x"434343",x"313131",x"333333",x"454545",x"4c4c4c",x"333333",x"535353",x"3c3c3c",x"333130",x"333130",x"000000",x"000000",x"000000",x"000000",x"3c3c3c",x"474747",x"414141",x"413f3e",x"4b4b4b",x"484848",x"3a3a3a",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3a1f0d",x"492812",x"37200f",x"422511",x"3e2511",x"150e07",x"412612",x"361f0f",x"2d1a0b",x"150e07",x"150e07",x"2e1a0b",x"402410",x"361e0d",x"4b392c",x"41240f",x"301b0c",x"371f0e",x"3a2210",x"321c0c",x"3c2310",x"371f0e",x"1b1108",x"150e07",x"4a2913",x"150e07",x"150e07",x"000000",x"675445",x"675445",x"5c5044",x"5d5044",x"6a5545",x"54493f",x"594f45",x"5a4f45",x"5d5146",x"594f46",x"554a40",x"544a3f",x"544a3f",x"000000",x"261809",x"261809",x"2b1b09",x"281909",x"39220d",x"39220d",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"3e3e3e",x"3e3e3e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3a2d",x"4d3a2d",x"150e07",x"412410",x"341d0d",x"412612",x"3f2411",x"311b0c",x"381f0e",x"39200f",x"150e07",x"2e1b0c",x"191007",x"181007",x"28180d",x"2c1b0e",x"331f10",x"311c0e",x"311c0e",x"2b180a",x"28160a",x"180f07",x"3d220f",x"4c3729",x"492c1a",x"462b19",x"3f2717",x"3e2516",x"3f2615",x"311d0f",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"191109",x"1c140c",x"201710",x"261c14",x"2a2017",x"291e16",x"291f17",x"291f17",x"281e16",x"482811",x"3b210e",x"3f2310",x"3f2410",x"371e0d",x"3e2310",x"3f2411",x"3f2411",x"341c0c",x"3e220f",x"3f2411",x"1c1108",x"654931",x"23180e",x"261a0d",x"281b0e",x"2d1e0e",x"2b1c0e",x"281c0f",x"2a1c0e",x"2f1f11",x"2f2011",x"2d1e11",x"291c0f",x"2b1c0f",x"2e1f10",x"2d1e11",x"291b0e",x"2c1e10",x"2a1d0f",x"322112",x"2e2012",x"2b1d0f",x"2f2011",x"2e1f12",x"261a0f",x"2d1f12",x"271a0e",x"271b0f",x"271a0d",x"2b1d0f",x"2b1c0d",x"25190c",x"25190c",x"261a0d",x"26190d",x"24180b",x"1f160d",x"412e1d",x"412e1d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584e43",x"584e43",x"50463d",x"423930",x"493224",x"40230f",x"2e1a0b",x"331c0c",x"3e2310",x"391f0d",x"402511",x"462914",x"402410",x"3f2410",x"402410",x"42240f",x"574d43",x"5e544b",x"584d43",x"594537",x"594537",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422511",x"422511",x"4e3221",x"3b2c21",x"4e453c",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"150e07",x"170f07",x"2b1d12",x"2e2017",x"342b23",x"342b23",x"000000",x"000000",x"4d3a2c",x"4d3a2c",x"4d2d16",x"38200f",x"311c0d",x"3b2210",x"301a0b",x"2f1a0b",x"150e07",x"301a0b",x"2d180a",x"2e190a",x"321c0c",x"351d0d",x"331c0c",x"341c0c",x"361e0d",x"361e0d",x"321c0c",x"331d0d",x"2f1a0b",x"331c0c",x"331d0d",x"331c0c",x"3a210f",x"311c0c",x"2d190b",x"2d190b",x"2d1a0b",x"351e0d",x"321d0d",x"2e190b",x"2e190b",x"2c180a",x"2a170a",x"261509",x"281609",x"2d190b",x"2c180b",x"2f1a0b",x"29170a",x"251509",x"27160a",x"2c180b",x"27160a",x"251509",x"261609",x"27160a",x"241409",x"231409",x"27160a",x"28160a",x"1d1108",x"1e1108",x"241509",x"27160a",x"25160a",x"221409",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2e17",x"4f2e17",x"150e07",x"150e07",x"1a1008",x"492c17",x"492c17",x"352e26",x"412410",x"412410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4e2c14",x"4e2c14",x"3f2511",x"3a2210",x"3e2310",x"402612",x"150e07",x"26160a",x"3c2310",x"150e07",x"331c0c",x"2d1a0b",x"2d180a",x"4d2c14",x"565656",x"525252",x"686868",x"383838",x"404040",x"373737",x"4e4e4e",x"6a6a6a",x"5d5d5d",x"4b4b4b",x"434343",x"414141",x"393939",x"464646",x"434343",x"4a4a4a",x"5a5a5a",x"606060",x"484848",x"323232",x"323232",x"626161",x"626161",x"5a5a59",x"525252",x"585858",x"393939",x"313131",x"414141",x"646363",x"4d4d4d",x"353535",x"353535",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"434343",x"454545",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"341c0c",x"472812",x"2c1a0c",x"412511",x"3d2411",x"39200e",x"3e2411",x"150e07",x"25160a",x"38200f",x"150e07",x"2c190b",x"412511",x"361e0e",x"4d3c30",x"3f230f",x"2c190b",x"351e0d",x"2c1a0c",x"331c0c",x"150e07",x"351d0d",x"201309",x"150e07",x"522f17",x"150e07",x"150e07",x"000000",x"605043",x"605043",x"5c5044",x"5d5145",x"605144",x"443022",x"392f26",x"41372d",x"615244",x"4b4137",x"4c3e33",x"483121",x"483121",x"000000",x"281909",x"281909",x"301e0a",x"2a1b09",x"36200b",x"36200b",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"434343",x"434343",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523d30",x"523d30",x"150e07",x"3f230f",x"331c0c",x"402612",x"331e0e",x"311b0b",x"150e07",x"371f0e",x"221409",x"2d1b0c",x"1b1108",x"191107",x"28180d",x"2d1b0f",x"341f11",x"331d0e",x"321c0e",x"2e190b",x"2a180a",x"180f07",x"381f0e",x"4c3a2e",x"4e301c",x"432a18",x"422917",x"422817",x"3e2514",x"25160b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"180f07",x"170f07",x"170f07",x"170f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"160f07",x"160f07",x"160f07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"171009",x"19120b",x"1d1610",x"1e1711",x"201912",x"211a14",x"211a14",x"1f1811",x"1f1812",x"4b2b13",x"3d220f",x"3e220f",x"3d220f",x"3b200e",x"3e2310",x"412410",x"3f2411",x"361d0c",x"3f2410",x"412511",x"211409",x"664b33",x"21160d",x"22170d",x"261a0e",x"291c0e",x"2a1c0e",x"251a0f",x"2d2011",x"2a1d10",x"2c1e10",x"261a0f",x"291c10",x"2b1e10",x"302113",x"291c0f",x"291c10",x"261a0f",x"2c1d0f",x"2b1c0f",x"291b0e",x"2c1d0f",x"2c1d0f",x"271b0f",x"261a10",x"271b0f",x"281b0f",x"261a0f",x"2a1c0f",x"2d1e0f",x"271b0e",x"281b0e",x"24180d",x"281b0e",x"281a0c",x"24170b",x"20170d",x"453321",x"453321",x"000000",x"4a4a4a",x"444444",x"646464",x"656565",x"323232",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"584e43",x"584e43",x"584d43",x"544a40",x"533a2a",x"3e230f",x"341d0d",x"341c0c",x"381f0e",x"381e0d",x"3f2410",x"3f2411",x"3f2310",x"3f2310",x"391f0d",x"3f220e",x"574d42",x"574d43",x"574c42",x"452712",x"452712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452812",x"452812",x"523624",x"3c2c20",x"4f453c",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"150e07",x"150e07",x"150e07",x"150e07",x"271910",x"302016",x"342b23",x"342b23",x"000000",x"000000",x"4b372a",x"4b372a",x"4e2e16",x"3c2311",x"341d0d",x"392110",x"38200f",x"2e190b",x"150e07",x"3a200e",x"38200e",x"371f0d",x"341d0c",x"2f1a0b",x"351d0d",x"361e0d",x"341d0d",x"351d0d",x"351e0d",x"311c0c",x"311c0c",x"341d0d",x"341d0d",x"341d0d",x"2e1a0b",x"29180a",x"231409",x"321c0c",x"2f1b0c",x"2a180b",x"2c190b",x"321d0d",x"2f1b0c",x"341d0d",x"301c0c",x"2e1a0b",x"29170a",x"271509",x"29170a",x"2d190b",x"2d1a0b",x"28160a",x"29170a",x"2a180a",x"231409",x"231409",x"1f1208",x"261509",x"231308",x"261409",x"271509",x"29170a",x"1f1208",x"221409",x"221409",x"231409",x"29180b",x"25160a",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"533018",x"533018",x"150e07",x"150e07",x"1c1108",x"4c2f19",x"4c2f19",x"44362c",x"432611",x"432611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"532f16",x"532f16",x"3d2410",x"38200f",x"3e2411",x"3d2310",x"321c0c",x"2e1a0b",x"3a2210",x"1e1209",x"341d0d",x"2d190b",x"2d180a",x"4e2c15",x"4e2c15",x"383838",x"404040",x"484848",x"4c4c4c",x"595959",x"4d4d4d",x"3e3e3e",x"3b3b3b",x"464646",x"454545",x"3d3d3d",x"393939",x"3d3d3d",x"000000",x"656565",x"5f5f5f",x"5c5c5c",x"505050",x"4a4a4a",x"363636",x"393939",x"4c4c4c",x"444444",x"494949",x"323232",x"333333",x"3b3b3b",x"4b4b4b",x"515151",x"3f3f3f",x"484848",x"353535",x"000000",x"000000",x"000000",x"000000",x"474747",x"444444",x"434343",x"454545",x"3a3735",x"444444",x"373737",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"422410",x"492812",x"29180b",x"442713",x"392110",x"361e0d",x"3b2210",x"331d0d",x"341e0e",x"37200f",x"150e07",x"311b0c",x"432712",x"361e0e",x"4c3e33",x"452711",x"321c0d",x"321c0d",x"180f07",x"371f0e",x"150e07",x"301b0c",x"2e190b",x"150e07",x"512f17",x"150e07",x"150e07",x"000000",x"000000",x"605043",x"5c5044",x"78624b",x"ac8e6c",x"b0916f",x"967d5e",x"947a5d",x"8c7358",x"957b5c",x"4c3e33",x"483121",x"483121",x"000000",x"2f1c0a",x"2f1c0a",x"2d1c0a",x"281a09",x"361f0b",x"361f0b",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"313131",x"414141",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"90765a",x"90765a",x"726352",x"564b40",x"523c2f",x"150e07",x"3f2310",x"331c0c",x"3e2411",x"1c1108",x"311b0b",x"150e07",x"38200f",x"2f1b0c",x"24150a",x"1d1308",x"1c1208",x"29190e",x"2e1c0f",x"331d0f",x"341d0e",x"321c0e",x"311b0c",x"2f1a0c",x"170f07",x"3c220f",x"4d3a2d",x"4b2e1a",x"452b18",x"382314",x"412816",x"3d2515",x"2b180c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"170f07",x"170f07",x"170f07",x"180f07",x"191008",x"191008",x"191008",x"191008",x"191008",x"191008",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"1c150e",x"1d160f",x"1f1912",x"1f1811",x"1e1811",x"1d160f",x"1c160f",x"4d2b13",x"3c210f",x"3e220f",x"3e2310",x"3a200e",x"402511",x"3a200e",x"412612",x"331c0c",x"3d2310",x"3e230f",x"1f1309",x"694c33",x"251a0f",x"22170d",x"25190d",x"281c0f",x"291c0f",x"271b0f",x"291c0f",x"281c10",x"2a1d11",x"261b0f",x"271b0f",x"291c0f",x"2a1e11",x"271b10",x"24190f",x"271a0f",x"271a0e",x"281a0e",x"2a1c0e",x"271a0d",x"2a1c0e",x"271a0e",x"251a0f",x"20160c",x"281b0f",x"2a1d0f",x"2b1d0f",x"2a1c0f",x"271a0d",x"25190e",x"261a0d",x"261a0d",x"25190c",x"281b0e",x"20170e",x"4d3826",x"4d3826",x"000000",x"4a4a4a",x"444444",x"646464",x"5b5b5b",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594f45",x"594f45",x"584e43",x"554b40",x"564134",x"371e0d",x"381f0e",x"381f0d",x"38200e",x"371e0d",x"3a200e",x"422612",x"412511",x"3a210f",x"381f0d",x"3a1f0d",x"28170a",x"574d43",x"574c42",x"452712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"412511",x"412511",x"533725",x"3c2c20",x"4e443a",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"150e07",x"150e07",x"150e07",x"170f07",x"2d1d11",x"2d1f15",x"352b23",x"352b23",x"000000",x"000000",x"503b2c",x"503b2c",x"533218",x"3b2210",x"38200e",x"3d2411",x"351e0e",x"2c180a",x"150e07",x"2f1a0b",x"301a0b",x"2d190b",x"311b0b",x"341d0d",x"371f0e",x"361f0e",x"37200e",x"371f0e",x"351e0d",x"37200e",x"39200e",x"341d0d",x"341d0d",x"301c0d",x"2b180a",x"2c190b",x"29170b",x"2c190b",x"2f1a0c",x"331c0d",x"321c0d",x"311c0c",x"321c0d",x"311c0d",x"341e0e",x"2f1b0c",x"2e1a0c",x"321c0c",x"2e1a0b",x"2a170a",x"2d180a",x"2b180b",x"2b180b",x"27160a",x"2a180b",x"2c190b",x"2a180a",x"29180b",x"2b180b",x"2f1a0b",x"211308",x"241509",x"1e1108",x"211309",x"25150a",x"150e07",x"25160a",x"221409",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2c15",x"4d2c15",x"150e07",x"150e07",x"1d1109",x"4e311d",x"4e311d",x"43362c",x"462711",x"462711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"563218",x"563218",x"3e2310",x"3a2210",x"2f1a0c",x"150e07",x"341d0d",x"150e07",x"150e07",x"321d0e",x"361e0d",x"2c190b",x"2f190b",x"4d2b14",x"3c3c3c",x"363636",x"323232",x"3f3f3f",x"363636",x"313131",x"3b3b3b",x"434343",x"3c3c3c",x"3e3e3e",x"3f3f3f",x"3a3a3a",x"333333",x"323232",x"363636",x"000000",x"606060",x"565656",x"353535",x"323232",x"373737",x"494949",x"363636",x"373737",x"424242",x"3a3a3a",x"323232",x"383838",x"454545",x"454545",x"333333",x"3d3d3d",x"616060",x"464646",x"000000",x"000000",x"3d3d3d",x"4f4f4f",x"454444",x"505050",x"575757",x"3b3b3b",x"373737",x"373636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"4c2b14",x"4c2b14",x"4d2c15",x"2f1b0d",x"3c220f",x"412612",x"361e0e",x"150e07",x"351e0d",x"150e07",x"150e07",x"2e1a0c",x"341d0d",x"452712",x"361e0d",x"503f32",x"462812",x"3a210f",x"331d0d",x"201309",x"361f0e",x"150e07",x"2e1a0c",x"351e0e",x"150e07",x"512f16",x"150e07",x"150e07",x"333333",x"3f3f3f",x"444444",x"866c54",x"78624b",x"ac8e6c",x"b0916f",x"967d5e",x"947a5d",x"8c7358",x"957b5c",x"957b5c",x"000000",x"484848",x"333333",x"323232",x"333333",x"333333",x"353433",x"3f3c39",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"323232",x"333333",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"90765a",x"90765a",x"726352",x"564b40",x"4e382a",x"150e07",x"432510",x"321b0b",x"2f1b0c",x"2e1b0c",x"341d0c",x"150e07",x"2a180b",x"361f0e",x"2e1a0c",x"191007",x"181007",x"2a1a0e",x"2f1c0f",x"341d0f",x"331d0e",x"301b0d",x"2c190b",x"2d190b",x"170f07",x"39200e",x"4e3c31",x"51321c",x"3d2314",x"3f2615",x"452b18",x"3f2715",x"25160b",x"180f07",x"201309",x"241509",x"1b1108",x"1f1309",x"211409",x"1f1309",x"211409",x"1d1208",x"211409",x"1c1108",x"231409",x"231409",x"1f1208",x"1e1208",x"201309",x"1a1008",x"241509",x"261609",x"231409",x"211409",x"251509",x"251509",x"211309",x"231409",x"211409",x"26160a",x"211409",x"211409",x"201409",x"211409",x"1d1208",x"201309",x"1d1208",x"1d1108",x"241509",x"231409",x"1d1108",x"1c1108",x"1c1108",x"1f1208",x"1c1108",x"221409",x"241509",x"26160a",x"1c1108",x"211309",x"251509",x"201309",x"221409",x"27160a",x"231409",x"190f08",x"241509",x"29180a",x"26160a",x"27170a",x"25160a",x"28170a",x"26160a",x"27160a",x"27160a",x"29170b",x"231509",x"1f1208",x"1f140a",x"291a10",x"2b1d11",x"2c1d11",x"291c12",x"2a1b10",x"22160d",x"4f2d15",x"361e0d",x"3c220f",x"39200f",x"381f0d",x"3d2310",x"3b200e",x"442712",x"361e0d",x"3c220f",x"3d220f",x"1c1108",x"6b4f36",x"231a10",x"21160d",x"22170d",x"271a0d",x"24190d",x"23180d",x"23180e",x"24190e",x"251a0e",x"24180d",x"23180e",x"291d10",x"2d1f11",x"281b0e",x"261a0f",x"23180d",x"23180d",x"2a1c0e",x"281b0e",x"2c1e0f",x"291b0e",x"291b0d",x"291c0e",x"281c0f",x"281b0e",x"261a0e",x"281a0d",x"2a1c0f",x"27190d",x"261a0d",x"271a0d",x"21170c",x"271b0e",x"291b0e",x"23190f",x"4c3725",x"4c3725",x"333333",x"333333",x"333333",x"333333",x"303030",x"353535",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594f45",x"594f45",x"594f45",x"584e44",x"482f1f",x"391f0d",x"381f0d",x"3a200e",x"3f2411",x"3c220f",x"391f0e",x"402511",x"38200e",x"402510",x"3a200d",x"3b200d",x"2c180a",x"2c180a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"533825",x"392a1f",x"554b41",x"150e07",x"150e07",x"150e07",x"150e07",x"29180b",x"150e07",x"150e07",x"150e07",x"190f08",x"2f1c11",x"2d1f15",x"352c24",x"352c24",x"000000",x"000000",x"503a2a",x"503a2a",x"4c2c15",x"3d2411",x"341e0e",x"3d2411",x"341e0e",x"2d190b",x"150e07",x"3a210f",x"39200f",x"39200e",x"38200e",x"3a200f",x"341d0d",x"2f1a0b",x"321c0c",x"341d0d",x"331c0c",x"311b0b",x"2b180b",x"2f1a0b",x"311c0c",x"311b0c",x"311b0c",x"27160a",x"351d0d",x"301b0c",x"331d0d",x"341d0d",x"2c180b",x"2a180a",x"321c0c",x"331d0d",x"29180b",x"361f0e",x"331d0d",x"321d0d",x"2a180b",x"321d0d",x"311c0d",x"2c190b",x"2d190b",x"2b180b",x"2a180a",x"2a170a",x"29170a",x"231409",x"211309",x"2f1b0b",x"2b180a",x"27160a",x"211208",x"26160a",x"211309",x"221409",x"24150a",x"201309",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2f17",x"4b2f17",x"150e07",x"150e07",x"201309",x"53331c",x"53331c",x"403329",x"452611",x"452611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"532f16",x"532f16",x"3d220f",x"3f2511",x"39200e",x"201309",x"39200e",x"150e07",x"26160a",x"351f0f",x"371f0d",x"2d1a0b",x"321b0c",x"4b2a12",x"474747",x"424242",x"4b4b4b",x"5d5d5d",x"4b4b4b",x"3e3e3e",x"575757",x"484848",x"474747",x"535353",x"646464",x"4f4f4f",x"323232",x"363636",x"363636",x"3a3a3a",x"373737",x"383838",x"323232",x"5b5b5b",x"5f5f5e",x"3e3e3e",x"474747",x"3c3c3c",x"3b3b3b",x"5e5e5e",x"515151",x"3d3d3d",x"484848",x"4d4d4d",x"444444",x"343434",x"616060",x"424242",x"3d3d3d",x"303030",x"3c3c3c",x"4d4d4d",x"5a5a5a",x"3e3e3e",x"363636",x"565656",x"5b5b5b",x"353535",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482813",x"482813",x"472813",x"301c0d",x"412511",x"402512",x"39200f",x"29180b",x"3c2311",x"1d1208",x"1c1108",x"38200f",x"331c0c",x"492a14",x"351d0c",x"504236",x"4a2b14",x"3c220f",x"351e0e",x"3d2411",x"38210f",x"150e07",x"201309",x"3d2411",x"150e07",x"502f16",x"150e07",x"323232",x"333333",x"3d3d3d",x"444444",x"181007",x"170f07",x"170f07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"545453",x"484848",x"333333",x"323232",x"333333",x"333333",x"353433",x"3f3c39",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"947b5e",x"947b5e",x"917d65",x"584d42",x"573f30",x"150e07",x"40230f",x"30190a",x"361e0e",x"412512",x"3a200e",x"150e07",x"2d190b",x"3c2310",x"2d1a0c",x"303030",x"323232",x"2a1a0f",x"2f1c0d",x"341d0f",x"321c0e",x"301c0d",x"311b0c",x"27160a",x"170f07",x"371e0d",x"49382c",x"4f321c",x"3f2717",x"3c2515",x"412815",x"3f2614",x"2a190c",x"1d1208",x"3d220e",x"1a130c",x"1a130c",x"17110a",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"180f07",x"180f07",x"191008",x"191008",x"1a1008",x"1a1008",x"191008",x"191008",x"191007",x"190f07",x"190f07",x"1a1007",x"191007",x"1a1008",x"191008",x"191008",x"190f08",x"1a110a",x"191109",x"18100a",x"18110a",x"412410",x"351d0c",x"422510",x"402411",x"3e2310",x"3f2411",x"381f0d",x"3f2511",x"381e0d",x"3d220f",x"39200e",x"3d220f",x"422511",x"211409",x"6b4e35",x"23180f",x"1e140b",x"1e150b",x"21170d",x"21160d",x"24190e",x"22170d",x"22170d",x"20160c",x"23180d",x"23180d",x"24190e",x"2a1c0f",x"291b0d",x"271b0d",x"261a0d",x"26190d",x"271a0e",x"291c0e",x"291b0e",x"261a0d",x"281b0e",x"281c0e",x"261a0e",x"271b0e",x"23170d",x"281b0d",x"281b0e",x"2a1c0d",x"22170b",x"281b0d",x"271a0c",x"281a0e",x"281a0e",x"20170d",x"513c27",x"513c27",x"000000",x"323232",x"323232",x"3f3f3f",x"424242",x"333333",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"594f45",x"594f45",x"584e44",x"4f301c",x"3d210e",x"361e0d",x"3b200f",x"3d2310",x"351e0d",x"3e2310",x"432713",x"3f2410",x"402511",x"381e0d",x"3c200d",x"2b180b",x"2b180b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"513523",x"37291f",x"544a40",x"150e07",x"150e07",x"150e07",x"150e07",x"201309",x"150e07",x"150e07",x"150e07",x"191008",x"2d1c11",x"332317",x"3a322a",x"3a322a",x"000000",x"000000",x"44362b",x"44362b",x"452711",x"3d2411",x"39210f",x"38210f",x"38200e",x"311c0c",x"150e07",x"3a210f",x"3b2210",x"3c2310",x"3b2210",x"3d2410",x"3d2310",x"3d2411",x"3e2511",x"3b2310",x"3a2210",x"3b2210",x"37200f",x"361f0e",x"331c0c",x"37200f",x"2c1a0b",x"331e0e",x"321c0d",x"341d0d",x"2b190b",x"2a180b",x"2f1a0b",x"351f0e",x"38210f",x"361f0f",x"331d0d",x"321d0d",x"321d0d",x"351e0e",x"341e0e",x"361f0e",x"2d1a0b",x"2d1a0b",x"29170a",x"251509",x"231409",x"1d1108",x"28170a",x"241509",x"2d190b",x"27160a",x"27160a",x"26160a",x"1c1008",x"211309",x"1d1108",x"241509",x"1d1108",x"211409",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"502f17",x"502f17",x"150e07",x"150e07",x"1f1209",x"4c2e19",x"4c2e19",x"42352b",x"452711",x"452711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"502e15",x"502e15",x"3d230f",x"402511",x"39200f",x"3f2310",x"412611",x"3a200f",x"150e07",x"3b2210",x"3b210e",x"311c0d",x"381f0e",x"472711",x"616161",x"5e5e5e",x"4a4a4a",x"454545",x"494949",x"494949",x"484848",x"4d4d4d",x"565656",x"585858",x"505050",x"545454",x"5a5a5a",x"676767",x"5d5d5d",x"373737",x"323232",x"474747",x"606060",x"313131",x"323232",x"323232",x"353535",x"373737",x"373737",x"323232",x"3d3d3d",x"5c5c5c",x"323232",x"595959",x"434343",x"454545",x"5f5f5f",x"323232",x"3d3d3d",x"4b4b4b",x"373737",x"5a5a5a",x"4e4e4e",x"313131",x"333333",x"323232",x"515151",x"313131",x"313131",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2a14",x"4a2a14",x"442511",x"2b190c",x"402410",x"432713",x"3a210f",x"3c2310",x"412511",x"402512",x"150e07",x"351f0f",x"381f0e",x"472913",x"341d0c",x"53463c",x"492b14",x"39210f",x"23150a",x"442813",x"3f2511",x"3b2210",x"150e07",x"331e0e",x"150e07",x"4c2a13",x"150e07",x"323232",x"323232",x"333333",x"333333",x"4f4f4f",x"1a1107",x"1b1208",x"1a1007",x"6f5a43",x"4d3e2e",x"554433",x"876f55",x"3c3c3b",x"646464",x"363636",x"323232",x"323232",x"313131",x"323232",x"343333",x"45413e",x"333333",x"313131",x"303030",x"323232",x"313131",x"313232",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"8f7659",x"8f7659",x"816d58",x"574c40",x"5c4638",x"150e07",x"432511",x"31190b",x"211409",x"412511",x"381f0e",x"3e2310",x"150e07",x"2f1b0c",x"26170a",x"606060",x"484848",x"29190c",x"2d1b0d",x"341d0f",x"311d0e",x"301c0d",x"301b0c",x"29170a",x"180f07",x"341d0c",x"45362a",x"472c19",x"482d18",x"3a2312",x"462b17",x"3e2412",x"311c0d",x"311c0d",x"19120b",x"19120b",x"171009",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f07",x"190f07",x"191008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"180f07",x"180f07",x"170f07",x"170f07",x"160e07",x"160e07",x"150e07",x"150e07",x"452510",x"452510",x"3a200e",x"3a210f",x"412511",x"381f0d",x"3f2410",x"3a1f0d",x"3c210f",x"3b210e",x"402410",x"402511",x"1a1108",x"6a4e35",x"20160c",x"1d140b",x"1f150b",x"1e140b",x"20160c",x"21170d",x"21160d",x"21170d",x"251a0f",x"24190f",x"23180d",x"24190e",x"2a1c0f",x"24190e",x"261a0d",x"261a0e",x"261a0d",x"291b0e",x"24190e",x"21170d",x"1f150b",x"23170d",x"22170d",x"21170d",x"21170d",x"21160d",x"20160c",x"2b1c0e",x"281b0d",x"2b1d0e",x"2a1c0e",x"2c1d0e",x"271a0c",x"22170b",x"1f150c",x"352619",x"352619",x"4b4b4b",x"5d5d5d",x"323232",x"3f3f3f",x"424242",x"323232",x"313130",x"383838",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2f1c",x"4d2f1c",x"3d200e",x"381f0d",x"391f0e",x"3d220f",x"331c0c",x"402512",x"3e2511",x"432712",x"422611",x"3a200e",x"3e230f",x"2d190b",x"2d190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e220f",x"3e220f",x"553823",x"35281e",x"53483f",x"150e07",x"150e07",x"150e07",x"150e07",x"27170a",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1c11",x"2d2016",x"3f372f",x"3f372f",x"000000",x"000000",x"45372c",x"45372c",x"4e2e17",x"402612",x"39210f",x"371f0e",x"361e0d",x"311c0c",x"150e07",x"371f0e",x"381f0e",x"39200f",x"3f2511",x"38200f",x"3d2311",x"39210f",x"39200f",x"3b2210",x"392110",x"38200f",x"37200f",x"37200f",x"2f1b0c",x"351e0d",x"2d190b",x"2d190b",x"301b0c",x"2d190b",x"2a180b",x"301c0c",x"301b0c",x"2f1a0b",x"301b0c",x"2f1b0b",x"2d1a0b",x"2d1a0b",x"2d1a0b",x"311c0c",x"301b0b",x"28170a",x"29170a",x"241408",x"241308",x"261509",x"27160a",x"27160a",x"28170a",x"271609",x"2a170a",x"271609",x"29170a",x"211309",x"1e1108",x"201308",x"221409",x"24150a",x"26160a",x"1f1309",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2a14",x"4a2a14",x"150e07",x"150e07",x"211409",x"53311a",x"53311a",x"3b3128",x"412410",x"412410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"533016",x"533016",x"3f2411",x"3f2411",x"3a210f",x"3c220f",x"3c220f",x"3c210f",x"150e07",x"3a2210",x"39200e",x"321c0d",x"38200f",x"482811",x"5d5d5c",x"4b4b4b",x"4e4e4e",x"565656",x"595959",x"575757",x"565656",x"3f3f3f",x"323232",x"323232",x"333333",x"353535",x"323232",x"323232",x"5c5c5c",x"4a4a4a",x"323232",x"434342",x"484848",x"323232",x"333333",x"414141",x"424242",x"000000",x"333333",x"494848",x"383838",x"515151",x"565656",x"505050",x"484848",x"4b4b4b",x"515151",x"515151",x"686868",x"616161",x"494949",x"525252",x"555555",x"434343",x"343332",x"3f3f3f",x"494846",x"636363",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"323232",x"323232",x"000000",x"000000",x"4a2a13",x"4a2a13",x"442510",x"2f1b0d",x"3f2310",x"3f2411",x"371f0e",x"412511",x"442813",x"422612",x"150e07",x"361f0f",x"361e0d",x"482913",x"39200f",x"544538",x"4d2c15",x"37200f",x"422612",x"432813",x"3c2411",x"3a2210",x"3c210f",x"241509",x"150e07",x"492912",x"150e07",x"323232",x"323232",x"333333",x"333333",x"333333",x"303030",x"333333",x"323232",x"444444",x"474747",x"494745",x"444444",x"333333",x"343434",x"323130",x"323333",x"333333",x"323232",x"646464",x"5c5c5c",x"5c5c5c",x"323232",x"333333",x"5c5c5c",x"595959",x"343434",x"323232",x"404040",x"414141",x"3e220f",x"3c210e",x"422510",x"422510",x"40230f",x"402310",x"3c200e",x"3a1f0d",x"391e0d",x"3c200d",x"3c200e",x"371c0c",x"3a1f0d",x"422511",x"452712",x"452813",x"3f2411",x"331d0d",x"3f2410",x"251509",x"665547",x"150e07",x"412410",x"311b0b",x"3e2310",x"3f2411",x"3a200e",x"3d230f",x"371f0e",x"180f07",x"2d1a0c",x"323232",x"323232",x"28180c",x"2d1b0d",x"351e0f",x"311c0d",x"2e190b",x"301b0b",x"2c190b",x"180f07",x"381f0e",x"4d3a2d",x"492b17",x"442917",x"3d2514",x"462915",x"3e2412",x"27170b",x"27170b",x"171009",x"171009",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"170f07",x"170f07",x"180f07",x"180f07",x"190f07",x"191008",x"191008",x"191008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"191008",x"180f08",x"180f07",x"160f07",x"160e07",x"160e07",x"150e07",x"150e07",x"4f2d14",x"4f2d14",x"3a200e",x"3d220f",x"3f2411",x"39200e",x"432611",x"3f220f",x"3d210e",x"3c210f",x"3e220f",x"452712",x"221409",x"674c33",x"1d140b",x"20160c",x"1d140b",x"1c130a",x"1e140b",x"1f150c",x"20150c",x"20150c",x"1f150b",x"22170d",x"1f150b",x"22170d",x"23180d",x"22170d",x"23180e",x"23180d",x"21170d",x"22170d",x"22170d",x"23180d",x"20150b",x"1e140b",x"1e140b",x"1f150b",x"1f150c",x"1f150b",x"1e140b",x"24180b",x"23170b",x"2e1e0d",x"281b0d",x"24170b",x"21160b",x"1d140b",x"1f160d",x"261b11",x"261b11",x"4b4b4b",x"5d5d5d",x"404040",x"4a4a4a",x"3c3c3c",x"3c3c3c",x"313130",x"343434",x"343434",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"503321",x"503321",x"3a1f0d",x"3a200e",x"341c0c",x"3a200e",x"371e0d",x"3e2310",x"3f2411",x"432712",x"412512",x"3c210f",x"452611",x"29170a",x"29170a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"422510",x"422510",x"4f3322",x"33251c",x"51473d",x"150e07",x"150e07",x"150e07",x"150e07",x"231509",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1d13",x"302319",x"423931",x"423931",x"000000",x"000000",x"49382b",x"49382b",x"4f2f17",x"3d2411",x"3a210f",x"38200e",x"341d0c",x"331d0d",x"150e07",x"3e2410",x"3b220f",x"39200f",x"3a210f",x"3e2410",x"3d2411",x"3d2411",x"3c2310",x"3e2511",x"3a2211",x"3c2311",x"3a2210",x"3a2210",x"37200f",x"361f0f",x"371f0e",x"37200f",x"2e1b0c",x"331d0d",x"311c0d",x"311c0c",x"2f1b0c",x"341d0d",x"301b0c",x"311b0c",x"331c0d",x"2e190b",x"2d190b",x"341d0d",x"2e1a0c",x"2a180b",x"301c0c",x"29180b",x"2f1b0c",x"2c190b",x"2b190b",x"2b180b",x"2c180b",x"2a180b",x"2d190b",x"241509",x"29170a",x"27160a",x"1f1208",x"241509",x"201308",x"241509",x"29180b",x"27170a",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e2411",x"3e2411",x"150e07",x"150e07",x"201309",x"54331b",x"54331b",x"3c2f25",x"422510",x"422510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"522f16",x"522f16",x"3e2411",x"412511",x"381f0e",x"3f2411",x"3b220f",x"3b200e",x"150e07",x"331c0c",x"3a200e",x"341d0d",x"3b210f",x"4f2d15",x"4f2d15",x"464646",x"414141",x"464646",x"414141",x"383737",x"323232",x"313131",x"323232",x"323232",x"333333",x"333333",x"323232",x"343434",x"332f2c",x"535353",x"565656",x"555555",x"323232",x"333333",x"333333",x"414141",x"444444",x"393939",x"535353",x"4f4f4f",x"545454",x"3d3d3d",x"313131",x"3a3a3a",x"3e3e3e",x"3e3e3e",x"4a4a4a",x"4e4e4e",x"373737",x"323232",x"353231",x"3a3a3a",x"434343",x"383838",x"323232",x"43403e",x"534f4c",x"686868",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"323232",x"323232",x"000000",x"4a2a13",x"4a2a13",x"472712",x"2f1c0d",x"412410",x"442813",x"361e0d",x"3f2411",x"402411",x"3a210f",x"150e07",x"341e0e",x"331c0d",x"462812",x"3b2210",x"5d4e42",x"482913",x"331e0e",x"3b2210",x"422713",x"3a2311",x"3a2210",x"341d0d",x"1a1008",x"150e07",x"422410",x"422511",x"301a0b",x"3f220f",x"391f0e",x"333333",x"333333",x"3f3f3f",x"454545",x"454545",x"383838",x"343434",x"313131",x"313131",x"343434",x"323232",x"333333",x"3f230f",x"333333",x"333333",x"333333",x"313131",x"313131",x"333333",x"333333",x"3d3b39",x"3c3a38",x"323232",x"2f2f2f",x"323232",x"3b200e",x"3e220f",x"3c210e",x"422510",x"422510",x"40230f",x"402310",x"3c200e",x"3a1f0d",x"391e0d",x"3c200d",x"3c200e",x"371c0c",x"3a1f0d",x"422511",x"452712",x"452813",x"3f2411",x"361f0e",x"3f2410",x"432712",x"261609",x"150e07",x"3e230f",x"361e0d",x"3b220f",x"39200e",x"361e0d",x"381f0e",x"371e0d",x"1a1008",x"211409",x"333333",x"323232",x"28170c",x"2e1b0d",x"331d0e",x"341d0e",x"321c0d",x"2f1b0c",x"2c190b",x"180f07",x"3d210f",x"513e31",x"4a2d18",x"402715",x"3f2614",x"412714",x"3e2413",x"2f1b0c",x"2f1b0c",x"422612",x"452713",x"472812",x"412410",x"3f220f",x"3d220f",x"412410",x"3d220f",x"3f230f",x"422511",x"40240f",x"3f230f",x"432511",x"452712",x"472812",x"462812",x"442712",x"452712",x"472913",x"492a13",x"482913",x"452712",x"452611",x"442611",x"452712",x"442611",x"432510",x"452711",x"422510",x"442711",x"442712",x"452812",x"472913",x"462712",x"402410",x"3e230f",x"3e220f",x"3c210f",x"3b200e",x"442610",x"3f220f",x"41240f",x"3e220e",x"3c210e",x"3f230f",x"3e210e",x"422410",x"432510",x"40240f",x"3a200d",x"3e210e",x"42240f",x"3c210e",x"41240f",x"3c210e",x"3d210e",x"3c200d",x"3e220e",x"3f220e",x"3f220e",x"432510",x"442510",x"422510",x"422510",x"432611",x"422511",x"412511",x"442611",x"482a14",x"150e07",x"492912",x"492912",x"402410",x"3a200e",x"3e2310",x"3f2410",x"412510",x"3c210f",x"381f0d",x"381f0d",x"3f2410",x"452813",x"1d1208",x"6a4c34",x"523c27",x"4b3623",x"4e3824",x"503a26",x"503a26",x"523b27",x"553e2a",x"503925",x"4a3421",x"4b3422",x"473321",x"493421",x"4a3421",x"4d3724",x"513a26",x"4f3825",x"493421",x"543c28",x"4d3724",x"4a3521",x"4b3520",x"4a3420",x"4a3520",x"483420",x"483320",x"4a3421",x"4a3422",x"463220",x"513924",x"4f3823",x"4f3823",x"4e3823",x"4c3724",x"4a3421",x"483321",x"422f1e",x"422f1e",x"323232",x"333333",x"313131",x"333333",x"313131",x"313131",x"323232",x"333333",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"462c1c",x"462c1c",x"3a200d",x"361d0c",x"351c0c",x"361d0d",x"381f0e",x"3c220f",x"3e2410",x"3f2310",x"462813",x"3b210e",x"432510",x"27160a",x"27160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"402410",x"402410",x"4e3220",x"36281e",x"544a3f",x"150e07",x"150e07",x"150e07",x"150e07",x"221409",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2016",x"36281d",x"463b32",x"463b32",x"000000",x"000000",x"483628",x"483628",x"513017",x"3e2411",x"371f0e",x"351d0d",x"2f1a0b",x"38200e",x"150e07",x"321c0c",x"2f1a0b",x"321c0c",x"331c0d",x"331c0c",x"371f0e",x"361e0d",x"351e0d",x"311c0c",x"341d0d",x"361e0d",x"341d0d",x"341d0d",x"361f0e",x"38200e",x"331d0d",x"361f0e",x"311d0d",x"311c0d",x"2f1a0c",x"331d0d",x"311b0c",x"351e0d",x"301b0c",x"341d0d",x"301b0c",x"2d190b",x"301b0c",x"321c0d",x"311c0c",x"2e1b0c",x"2c190b",x"301c0d",x"2f1c0c",x"2e1a0c",x"2c1a0b",x"2b190b",x"2d1a0b",x"27160a",x"29180a",x"2c190b",x"211309",x"27160a",x"231409",x"251509",x"1b1008",x"211409",x"27160a",x"24150a",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482914",x"482914",x"150e07",x"150e07",x"1e1209",x"51321a",x"51321a",x"332b23",x"422411",x"422411",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"553116",x"553116",x"402511",x"432712",x"3a210f",x"3e2310",x"3c220f",x"402511",x"2f1b0d",x"38200e",x"412511",x"2f1b0c",x"3c210f",x"4c2a13",x"4c2a13",x"000000",x"404040",x"464646",x"414141",x"383737",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"5f5e5d",x"5f5e5d",x"616161",x"555555",x"2f2f2f",x"474747",x"474747",x"323232",x"494949",x"4c4c4c",x"393939",x"353535",x"6d6a68",x"616060",x"515151",x"444444",x"323232",x"323232",x"4e4e4e",x"525252",x"4e4e4e",x"4b4b4b",x"505050",x"4d4d4d",x"3a3a3a",x"393939",x"343433",x"3f3f3f",x"393939",x"3d3d3d",x"666666",x"343333",x"383838",x"363636",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"303030",x"373737",x"373737",x"000000",x"492a14",x"492a14",x"472913",x"2b190c",x"3f230f",x"432713",x"361e0e",x"412511",x"3e2310",x"432713",x"2c1a0c",x"39210f",x"371f0e",x"4d2c14",x"3e2311",x"54473c",x"452711",x"3e2310",x"2c190b",x"381f0e",x"381f0e",x"381f0e",x"150e07",x"2b180b",x"381f0e",x"3d210e",x"3a210e",x"422510",x"3f240f",x"614f40",x"695647",x"422510",x"371e0c",x"381f0e",x"3c210e",x"3b210e",x"351d0d",x"3c220f",x"422410",x"472712",x"402310",x"432611",x"422510",x"462812",x"492913",x"482812",x"442610",x"452611",x"452611",x"442611",x"452712",x"4c2c15",x"432611",x"3e220f",x"452711",x"3a1f0d",x"3b200d",x"3d200e",x"412310",x"3f230f",x"422510",x"42230e",x"452610",x"442510",x"3e210e",x"40230f",x"422410",x"41240f",x"422510",x"40230f",x"432510",x"452812",x"462813",x"452712",x"432510",x"412411",x"3f2310",x"442712",x"422511",x"412511",x"27170a",x"3b210e",x"3a200e",x"3a200e",x"150e07",x"311b0c",x"2d190b",x"2d190b",x"8d7458",x"27170b",x"2d1a0d",x"331d0e",x"331c0c",x"341e0e",x"2f1a0b",x"28170a",x"180f07",x"3d230f",x"534133",x"4e2f19",x"3c2413",x"382211",x"3f2514",x"3e2311",x"27160b",x"27160b",x"17110a",x"171009",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f08",x"180f07",x"170f07",x"170f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"19120b",x"1c150e",x"1c150e",x"1a120b",x"1a120b",x"4c2b14",x"4c2b14",x"3d220f",x"3f2410",x"422511",x"3e230f",x"412511",x"3d220f",x"3c200e",x"3e220f",x"402310",x"442712",x"201309",x"6a4c34",x"523c27",x"4b3623",x"4e3824",x"503a26",x"503a26",x"523b27",x"553e2a",x"503925",x"4a3421",x"4b3422",x"473321",x"493421",x"4a3421",x"4d3724",x"513a26",x"4f3825",x"493421",x"543c28",x"4d3724",x"4a3521",x"4b3520",x"4a3420",x"4a3520",x"483420",x"483320",x"4a3421",x"4a3422",x"463220",x"513924",x"4f3823",x"4f3823",x"4e3823",x"4c3724",x"4a3421",x"483321",x"422f1e",x"333333",x"333333",x"333333",x"323232",x"333333",x"333333",x"333333",x"323232",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d3324",x"4d3324",x"3e220f",x"331b0b",x"371e0c",x"321b0b",x"381f0e",x"351d0d",x"3e2310",x"402411",x"422612",x"39200e",x"42240f",x"2d190b",x"2d190b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3f230f",x"3f230f",x"4d3222",x"36281e",x"564d43",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1108",x"150e07",x"150e07",x"150e07",x"1c1108",x"342418",x"37291f",x"443b32",x"443b32",x"000000",x"000000",x"4a392d",x"4a392d",x"4e2d16",x"3b2310",x"351e0d",x"371e0d",x"321b0c",x"351d0d",x"150e07",x"301b0c",x"351d0d",x"381f0e",x"361f0d",x"321c0c",x"331c0c",x"311b0c",x"341d0d",x"351e0d",x"351d0d",x"351d0d",x"331c0d",x"351e0d",x"331c0d",x"321d0d",x"321c0c",x"301b0c",x"2d190b",x"2a180a",x"2f1a0b",x"331d0d",x"2d190b",x"331c0c",x"311c0c",x"331d0c",x"321c0d",x"2e1a0b",x"2c190b",x"251509",x"2b180a",x"2d190b",x"2c180b",x"2b180b",x"2a180b",x"311c0c",x"2b180b",x"26160a",x"29180a",x"25150a",x"29180b",x"2a180b",x"26160a",x"221309",x"231409",x"241509",x"191008",x"1b1008",x"231409",x"241509",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"452812",x"452812",x"150e07",x"150e07",x"211409",x"5c381e",x"5c381e",x"43342b",x"3f2310",x"3f2310",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"543116",x"543116",x"422612",x"412511",x"3c230f",x"2f1b0c",x"402410",x"150e07",x"341d0d",x"3a210f",x"3f230f",x"2f1a0b",x"3f230f",x"512d15",x"512d15",x"000000",x"363636",x"3e3e3e",x"444444",x"464645",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"605f5f",x"5c5a59",x"4e4e4e",x"323232",x"484848",x"515151",x"595959",x"585858",x"525252",x"303131",x"313131",x"6d6b6a",x"676767",x"525252",x"595959",x"323232",x"313131",x"515151",x"4d4d4d",x"4f4f4f",x"525252",x"4a4a4a",x"505050",x"5f5f5f",x"686868",x"606060",x"626261",x"696969",x"676767",x"363636",x"3a3a3a",x"343333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"312f2f",x"454545",x"454545",x"000000",x"482912",x"482912",x"4e2d16",x"361f0f",x"412411",x"442813",x"39200f",x"392110",x"3b200e",x"150e07",x"3e2511",x"38200f",x"3a220f",x"482913",x"38200e",x"4c3d33",x"40230f",x"361d0d",x"381e0d",x"371e0d",x"2e190b",x"311b0b",x"150e07",x"2a170a",x"311a0b",x"341c0c",x"351d0c",x"361d0c",x"331a0b",x"5f5144",x"5c4d41",x"2e1709",x"2b1508",x"2f190a",x"361d0c",x"381f0d",x"361e0d",x"351e0d",x"3a200e",x"381f0d",x"3b200e",x"3e230f",x"3b200e",x"3a200e",x"3c210f",x"3a200e",x"3b200e",x"39200e",x"3d210f",x"3b210e",x"371e0d",x"361d0c",x"381e0c",x"3a1f0d",x"3c210e",x"371e0d",x"3e220f",x"3a200e",x"3b210f",x"3c210f",x"3c210f",x"3d210e",x"3b200d",x"3a200e",x"381e0c",x"351c0c",x"3b200d",x"3d210e",x"3c210e",x"3d210f",x"3c210e",x"3a200e",x"381f0d",x"351c0c",x"261207",x"251106",x"251207",x"291408",x"2e1709",x"2a1508",x"30190b",x"30190b",x"341c0c",x"381f0d",x"150e07",x"321c0c",x"2d190b",x"90775a",x"8d7458",x"27170b",x"2f1b0d",x"311b0c",x"331c0c",x"331d0d",x"2e1a0b",x"2a180a",x"180f07",x"412611",x"4f3f33",x"503019",x"402614",x"382211",x"3f2513",x"3e2311",x"28160b",x"28160b",x"17110a",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"180f07",x"180f07",x"170f07",x"170f07",x"170f07",x"160f07",x"170f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"19130c",x"1b140d",x"1c150e",x"1b150d",x"1c150e",x"1c150e",x"452712",x"452712",x"3c210e",x"3e2310",x"3f2410",x"3f2410",x"3f230f",x"3a200e",x"3e230f",x"3c210f",x"3e2310",x"452712",x"201309",x"201309",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"333333",x"333333",x"323232",x"323232",x"333333",x"333333",x"333333",x"32302f",x"323232",x"323232",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"523a2a",x"523a2a",x"40230f",x"351d0c",x"331d0c",x"321c0c",x"341d0d",x"39200e",x"412511",x"422611",x"422611",x"3b210f",x"432510",x"25160a",x"25160a",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3b210f",x"3b210f",x"513321",x"34271e",x"574e44",x"150e07",x"150e07",x"150e07",x"150e07",x"231409",x"150e07",x"150e07",x"150e07",x"170f07",x"33241a",x"35271e",x"433930",x"433930",x"000000",x"000000",x"42352a",x"42352a",x"4f2e16",x"3a2210",x"341e0d",x"321c0c",x"311c0c",x"311b0c",x"150e07",x"361f0e",x"361f0e",x"381f0e",x"341d0d",x"331d0d",x"331d0d",x"341d0d",x"321c0c",x"2f1a0b",x"2e190b",x"2e1a0b",x"301b0c",x"321c0c",x"301a0b",x"2e1a0b",x"2c180b",x"2b180a",x"2c180a",x"281509",x"29160a",x"2c180a",x"271609",x"2b180a",x"2b180a",x"281609",x"261509",x"221308",x"211208",x"1f1108",x"251409",x"281609",x"2c190b",x"27160a",x"2a180a",x"28160a",x"231409",x"241509",x"231409",x"201309",x"27160a",x"28170a",x"251509",x"261509",x"221309",x"29170a",x"211409",x"1c1108",x"28170b",x"201309",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2c14",x"4c2c14",x"150e07",x"150e07",x"1c1108",x"52311a",x"52311a",x"3d3128",x"452712",x"452712",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"532f16",x"532f16",x"432712",x"3f2410",x"3e2310",x"3e2310",x"39200e",x"3a210f",x"412511",x"39200d",x"3d220e",x"301b0b",x"351d0b",x"4d2a12",x"4d2a12",x"484848",x"363636",x"3e3e3e",x"444444",x"464645",x"525252",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5c5a59",x"484848",x"393939",x"343434",x"555555",x"4b4b4b",x"3c3c3c",x"363636",x"333333",x"333333",x"363636",x"363636",x"676767",x"4c4c4c",x"434343",x"363636",x"000000",x"000000",x"313131",x"4a4a4a",x"484848",x"4a4a4a",x"434343",x"404040",x"474747",x"555555",x"535353",x"454343",x"333434",x"323232",x"313131",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"3e3e3e",x"3e3e3e",x"000000",x"4b2a13",x"4b2a13",x"4f2d15",x"341f0e",x"462914",x"4a2c15",x"3d2210",x"452813",x"3b2210",x"371f0e",x"3a2210",x"3b2210",x"3f2511",x"492913",x"361f0e",x"543c2c",x"482913",x"39200f",x"3c220f",x"371f0e",x"351d0d",x"341d0d",x"311c0c",x"2b190b",x"371f0e",x"3b210f",x"3b200e",x"3c210f",x"422611",x"432611",x"412511",x"402411",x"412511",x"3d2310",x"402411",x"3c210f",x"3e220f",x"3e230f",x"422612",x"452813",x"432612",x"432611",x"442813",x"3c210f",x"402310",x"3e230f",x"3f2410",x"3a200e",x"3a200e",x"3b200e",x"3c210f",x"3d220f",x"32190a",x"3b200e",x"422410",x"3a200d",x"3a1f0d",x"391f0d",x"381e0d",x"3b200e",x"402410",x"412511",x"3e220f",x"3f2410",x"381e0d",x"391f0d",x"391f0d",x"3b200d",x"381e0d",x"391f0d",x"3a200e",x"391f0d",x"3f230f",x"3c210f",x"371e0d",x"361d0c",x"3f2310",x"3c220f",x"391f0d",x"361e0d",x"381f0e",x"321c0c",x"351d0d",x"341d0c",x"2e190b",x"251509",x"1e1208",x"170f07",x"1a1107",x"26160a",x"2e1a0b",x"311b0c",x"321b0c",x"311b0c",x"2d190b",x"27160a",x"180f08",x"3b2310",x"45382d",x"4c2d17",x"462b17",x"3e2513",x"3f2412",x"3f2411",x"422512",x"422512",x"19120c",x"171009",x"171009",x"17110a",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160e07",x"160f07",x"170f07",x"170f07",x"180f07",x"180f07",x"180f07",x"190f08",x"190f08",x"190f08",x"190f08",x"170f07",x"170f07",x"180f07",x"170f07",x"160f07",x"160e07",x"160e07",x"160e07",x"160e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"171009",x"1a130c",x"1c150e",x"1e1710",x"1d170f",x"1d160e",x"1d160e",x"402410",x"402410",x"3e220f",x"422511",x"422611",x"3f2410",x"3f230f",x"3c210e",x"412511",x"3d220f",x"402410",x"412510",x"1e1208",x"2b180b",x"26150a",x"221309",x"28170a",x"29170a",x"251509",x"27160a",x"231409",x"29170a",x"28160a",x"28170a",x"29170a",x"231409",x"28170a",x"25150a",x"2c190b",x"2b180a",x"28170a",x"2a170a",x"23150a",x"28170a",x"2c190b",x"2b190b",x"2c190b",x"2a180b",x"2a180a",x"23140a",x"27160a",x"27170a",x"29180b",x"25150a",x"27160a",x"231409",x"231409",x"241509",x"241509",x"211409",x"2c190b",x"27160a",x"28160a",x"221409",x"26160a",x"29170b",x"26160a",x"2d190b",x"2b190b",x"27160a",x"231409",x"28160b",x"2b190b",x"29180b",x"29170a",x"2b180b",x"29180b",x"2d190c",x"2a180b",x"2f1a0c",x"2a180a",x"27160a",x"28180b",x"271a0f",x"2d1c10",x"2c1c11",x"523c2d",x"412410",x"381e0d",x"381f0d",x"371e0d",x"391f0e",x"391f0d",x"412511",x"432612",x"462812",x"3e230f",x"462711",x"29160a",x"3c220f",x"402410",x"3b210e",x"3f230f",x"3f230f",x"3c210e",x"3c210f",x"3b200e",x"3f2410",x"3f2410",x"3c220f",x"3e230f",x"3e230f",x"000000",x"000000",x"000000",x"000000",x"3f2310",x"3f2310",x"513321",x"36271d",x"554b41",x"150e07",x"150e07",x"150e07",x"150e07",x"1e1208",x"150e07",x"150e07",x"150e07",x"1a1008",x"332419",x"32251c",x"40382f",x"40382f",x"000000",x"000000",x"524034",x"524034",x"4e2d16",x"3b2310",x"37200f",x"37200e",x"341d0d",x"351d0d",x"150e07",x"341d0c",x"321b0c",x"321b0b",x"321b0b",x"331c0c",x"331d0d",x"38200e",x"351d0d",x"321c0c",x"311b0c",x"331d0d",x"38200e",x"341e0d",x"351e0d",x"361e0e",x"331d0d",x"341d0d",x"2e190b",x"331c0c",x"321c0c",x"2a180a",x"2e1a0b",x"2d190b",x"2f1a0b",x"2f1b0c",x"2e1a0c",x"321c0d",x"301c0d",x"301c0d",x"2d1a0b",x"301b0c",x"2e1a0b",x"2c190b",x"2b180b",x"28170b",x"301c0d",x"26160a",x"2d1a0b",x"2d1a0c",x"2a180b",x"25150a",x"28170a",x"211309",x"241509",x"241509",x"26160a",x"201309",x"26160a",x"211409",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4c2b14",x"4c2b14",x"150e07",x"150e07",x"1d1209",x"55341c",x"55341c",x"362f26",x"462812",x"462812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"533016",x"533016",x"402411",x"3f230f",x"3f2310",x"432612",x"442712",x"3e2310",x"3a200f",x"3b200e",x"3b200d",x"311b0b",x"361e0d",x"42240e",x"393939",x"464646",x"4e4e4e",x"5c5c5c",x"575757",x"565656",x"464646",x"3f3f3f",x"000000",x"414141",x"565656",x"5b5b5b",x"424242",x"414141",x"4d4d4d",x"4b4b4b",x"363636",x"333333",x"363636",x"4c4c4c",x"5c5c5c",x"5b5b5b",x"4e4e4e",x"363636",x"373737",x"434343",x"4c4c4c",x"434343",x"3f3f3f",x"333333",x"343434",x"313131",x"333333",x"323232",x"494949",x"484848",x"464646",x"575757",x"494949",x"363636",x"383838",x"313131",x"353535",x"454545",x"515151",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"343434",x"434343",x"4f4f4f",x"000000",x"4b2a14",x"4b2a14",x"472712",x"2f1c0d",x"4b2c15",x"432713",x"39200f",x"472a14",x"452914",x"422713",x"3d2411",x"3e2310",x"3e2411",x"452711",x"3a210f",x"463226",x"3f210e",x"2e190b",x"311a0b",x"1b1008",x"2e1a0b",x"150e07",x"211309",x"1f1208",x"301b0b",x"371f0d",x"3d220f",x"3f2410",x"3e2310",x"402410",x"3f2310",x"3e230f",x"3e220f",x"3a200e",x"391f0d",x"381e0d",x"361e0d",x"381f0d",x"3b200e",x"3b210f",x"3a200e",x"3a200e",x"361d0d",x"361d0c",x"381e0d",x"381e0d",x"3a1f0d",x"371e0d",x"3b200e",x"3b200e",x"381e0d",x"391f0d",x"3a200d",x"371e0d",x"381e0d",x"3a200e",x"381f0d",x"3c210e",x"3d210e",x"391f0d",x"381e0d",x"3b210e",x"412410",x"3f2410",x"3c210f",x"3f230f",x"3f2310",x"3b210f",x"3e230f",x"3a200e",x"3d220f",x"391f0e",x"402310",x"422511",x"3f2410",x"3a210f",x"3a200e",x"381f0d",x"391f0d",x"301a0b",x"331c0b",x"201208",x"2e1a0b",x"150e07",x"1d1208",x"1e1208",x"29170a",x"170f07",x"181007",x"271609",x"2c180b",x"321c0c",x"321c0c",x"321c0c",x"2e190b",x"2a170a",x"180f07",x"472a14",x"4d3e33",x"4a2c16",x"432915",x"3f2613",x"3d2411",x"382010",x"412411",x"341e0e",x"361f0e",x"371f0d",x"301b0c",x"331c0d",x"301b0b",x"2d190b",x"301b0b",x"2e190b",x"2d1a0b",x"39200f",x"371f0d",x"2f1b0c",x"331c0c",x"371f0d",x"361e0d",x"361f0e",x"361e0e",x"361e0d",x"2f1b0c",x"321c0c",x"321c0c",x"2c190b",x"331d0d",x"361f0e",x"321c0d",x"361f0e",x"371f0d",x"341e0d",x"341d0d",x"341d0d",x"331c0c",x"2b180b",x"301a0b",x"2f1b0b",x"2d190b",x"321c0c",x"361e0d",x"2e190b",x"311b0b",x"311a0c",x"2c180a",x"321c0c",x"351d0d",x"2f1a0b",x"331c0c",x"2e1a0b",x"301a0b",x"301a0b",x"321c0c",x"331d0c",x"2f1b0c",x"351d0d",x"371e0d",x"301b0c",x"331c0c",x"341d0c",x"2e190b",x"341c0c",x"341c0c",x"351d0d",x"321b0c",x"351d0d",x"331c0c",x"2f1a0b",x"341d0c",x"39200e",x"321c0c",x"38200e",x"3c2210",x"301b0c",x"361e0d",x"472711",x"371f0d",x"3d220f",x"3c220f",x"3b200e",x"3d220f",x"39200e",x"3a200e",x"371f0d",x"3f230f",x"3e230f",x"2b180b",x"2b180b",x"26150a",x"221309",x"28170a",x"29170a",x"251509",x"27160a",x"231409",x"29170a",x"28160a",x"28170a",x"29170a",x"231409",x"28170a",x"25150a",x"2c190b",x"2b180a",x"28170a",x"2a170a",x"23150a",x"28170a",x"2c190b",x"2b190b",x"2c190b",x"2a180b",x"2a180a",x"23140a",x"27160a",x"27170a",x"29180b",x"25150a",x"27160a",x"231409",x"231409",x"241509",x"241509",x"211409",x"2c190b",x"27160a",x"28160a",x"221409",x"26160a",x"29170b",x"26160a",x"2d190b",x"2b190b",x"27160a",x"231409",x"28160b",x"2b190b",x"29180b",x"29170a",x"2b180b",x"29180b",x"2d190c",x"2a180b",x"2f1a0c",x"2a180a",x"27160a",x"28180b",x"271a0f",x"2d1c10",x"2c1c11",x"2c1b0f",x"402410",x"321c0c",x"341c0c",x"371e0d",x"371f0d",x"371e0d",x"3c220f",x"3c220f",x"402511",x"39200f",x"402410",x"3a210e",x"3c220f",x"402410",x"3b210e",x"3f230f",x"3f230f",x"3c210e",x"3c210f",x"3b200e",x"3f2410",x"3f2410",x"3c220f",x"3e230f",x"3e230f",x"000000",x"000000",x"000000",x"000000",x"3f230f",x"3f230f",x"543624",x"35281f",x"584e44",x"150e07",x"150e07",x"150e07",x"150e07",x"211309",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2017",x"2e221a",x"3b332b",x"3b332b",x"000000",x"000000",x"4a3e34",x"4a3e34",x"4e2e16",x"3a2210",x"37200f",x"3c2310",x"361f0e",x"331c0d",x"150e07",x"311b0b",x"321c0c",x"351d0d",x"321b0c",x"331c0c",x"311b0c",x"301a0b",x"311b0b",x"2e190b",x"2e190b",x"301b0b",x"2c180a",x"2b170a",x"2d180a",x"29160a",x"2a170a",x"2e190b",x"311b0b",x"2c190b",x"2c180a",x"28170a",x"2f1a0b",x"2f1a0b",x"311c0d",x"2f1b0c",x"301c0c",x"301b0c",x"2f1a0b",x"2e1a0b",x"2a170a",x"2a180a",x"261609",x"27160a",x"29170a",x"2b180b",x"2a180b",x"2a180b",x"2a170a",x"2a170a",x"28170a",x"27160a",x"261509",x"27160a",x"251509",x"221409",x"221409",x"231409",x"23150a",x"1a1008",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2a14",x"4a2a14",x"150e07",x"150e07",x"1f1309",x"5c381e",x"5c381e",x"423226",x"442611",x"442611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"563217",x"563217",x"3a200e",x"3b210e",x"412411",x"422511",x"3c210e",x"402410",x"341c0b",x"381f0c",x"391f0d",x"311b0b",x"361e0c",x"3f220d",x"333333",x"606060",x"343434",x"313131",x"363636",x"4a4a4a",x"424242",x"373737",x"474747",x"313131",x"414141",x"5b5b5b",x"353535",x"555555",x"505050",x"363636",x"404040",x"5d5d5d",x"474747",x"3c3c3c",x"353535",x"363636",x"343434",x"535353",x"5e5e5e",x"646464",x"424242",x"404040",x"3b3b3b",x"3d3d3d",x"343434",x"343434",x"565656",x"565656",x"4d4d4d",x"434343",x"424242",x"494949",x"424242",x"4a4a4a",x"4d4d4d",x"4f4f4f",x"555555",x"4f4f4f",x"595959",x"595959",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"323232",x"313131",x"323232",x"000000",x"4a2a13",x"4a2a13",x"492912",x"2f1b0c",x"4d2e16",x"412611",x"402511",x"432713",x"402612",x"422612",x"3e2310",x"3f2411",x"402511",x"442612",x"39210f",x"48382c",x"4a2a13",x"351d0d",x"331c0c",x"2e1a0b",x"311c0d",x"26160a",x"2a170a",x"201208",x"341d0d",x"371f0e",x"3a200f",x"3f2410",x"3f2410",x"422611",x"422611",x"442712",x"412411",x"3f2411",x"3f2410",x"3f2410",x"3b200f",x"3f2410",x"412511",x"3f2411",x"3f2410",x"442611",x"3c210f",x"371f0d",x"3e230f",x"3f2410",x"412411",x"402411",x"3e2310",x"3b210f",x"3f2310",x"3f230f",x"412510",x"412511",x"3b200e",x"391f0d",x"381f0d",x"3b200e",x"3c210f",x"3e220f",x"391f0e",x"3b200e",x"3b200e",x"3d220f",x"3f2310",x"3f240f",x"402410",x"3d220f",x"361c0c",x"3f2310",x"422511",x"412411",x"412511",x"3b200d",x"391f0c",x"361e0c",x"42250f",x"381f0d",x"3a200e",x"301a0b",x"2c1709",x"251509",x"261509",x"271509",x"261509",x"170f07",x"251509",x"251509",x"29170a",x"29170a",x"2e1a0b",x"311b0c",x"331c0d",x"321c0d",x"2d190b",x"2a180a",x"180f07",x"361f0f",x"41372d",x"3d2211",x"351e0f",x"382010",x"361d0e",x"3a200f",x"3c2210",x"3f2311",x"3c2110",x"3e2210",x"3a200e",x"3f230f",x"3e220f",x"3b200e",x"3e220f",x"3d220f",x"39200e",x"412511",x"422511",x"412511",x"412511",x"412410",x"3d210e",x"3c210f",x"422611",x"462812",x"381f0d",x"361d0c",x"38200e",x"3a210f",x"3c210f",x"3e2310",x"422611",x"412511",x"412511",x"3f2411",x"3e2310",x"422612",x"3b2210",x"3b210f",x"432612",x"3f2310",x"402410",x"3b220f",x"402411",x"3b210f",x"412410",x"3a200e",x"3b210f",x"422611",x"422611",x"412511",x"402411",x"3e230f",x"3f2410",x"402410",x"3d220f",x"3d220f",x"3e230f",x"361d0c",x"391e0d",x"3b200e",x"3c210e",x"3c210f",x"3d210e",x"381f0d",x"3a200e",x"3b200e",x"3e220f",x"402410",x"3f2410",x"452712",x"391f0d",x"3a200e",x"3f230f",x"432611",x"462812",x"442610",x"371e0c",x"3b200d",x"3c210e",x"412511",x"3d220f",x"3e220f",x"351c0b",x"391f0d",x"351c0c",x"331a0b",x"361d0c",x"3a1f0d",x"3b1f0d",x"3d210d",x"3b200d",x"3c200e",x"3a200d",x"391f0d",x"391f0d",x"3b200e",x"3f230f",x"3b200e",x"361c0c",x"381d0c",x"361c0c",x"331b0b",x"351c0b",x"361c0c",x"361d0c",x"351d0c",x"3b200e",x"381f0d",x"3a200e",x"381f0d",x"381f0e",x"3a200e",x"3e230f",x"3d220f",x"402410",x"402410",x"3f2310",x"3e2310",x"3d220f",x"3e2310",x"402410",x"412511",x"3a200e",x"361e0d",x"3a200e",x"422611",x"3e220f",x"391f0d",x"361e0d",x"3d220f",x"3c210f",x"39200f",x"422611",x"432611",x"402511",x"432712",x"3f2511",x"3e2310",x"432712",x"3f2410",x"422611",x"412410",x"452712",x"402511",x"442712",x"432611",x"402410",x"3f230f",x"3d220f",x"3f2310",x"402411",x"412510",x"3b210f",x"3f2410",x"381f0e",x"3f2410",x"3d220f",x"3e230f",x"3d220f",x"3b200e",x"3b200e",x"3b200e",x"3c210e",x"40240f",x"39200e",x"3a200e",x"3c210e",x"3d220f",x"402410",x"3f2310",x"422511",x"412410",x"3f2310",x"371c0c",x"3c210f",x"432612",x"4b2a14",x"4b2a14",x"000000",x"000000",x"000000",x"000000",x"3b200e",x"3b200e",x"523726",x"34271e",x"544a3f",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"2f2117",x"2f2219",x"342c25",x"342c25",x"000000",x"000000",x"40332a",x"40332a",x"4c2d15",x"37200f",x"38200f",x"39210f",x"38200e",x"39200f",x"150e07",x"321c0c",x"311b0c",x"341d0d",x"331d0d",x"361e0d",x"331c0c",x"321c0d",x"341d0d",x"341d0d",x"351e0d",x"351e0e",x"361f0e",x"351e0d",x"331d0d",x"2d190b",x"301b0b",x"341e0d",x"311c0c",x"2a180a",x"2c180a",x"331d0d",x"371f0e",x"301b0c",x"331d0d",x"2b190b",x"321d0d",x"301c0d",x"301c0d",x"311c0d",x"311c0d",x"2f1b0c",x"2e1b0c",x"311c0d",x"2f1b0c",x"301c0c",x"2e1a0c",x"2e1b0c",x"26160a",x"26160a",x"28170a",x"2a180b",x"2e1b0c",x"1a1008",x"1d1108",x"241509",x"231409",x"241509",x"211409",x"211409",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2b14",x"4a2b14",x"150e07",x"150e07",x"23150a",x"55331b",x"55331b",x"403227",x"452711",x"452711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"573117",x"573117",x"391f0d",x"3b200e",x"402410",x"412511",x"3f2411",x"3f2511",x"3d220e",x"3f230f",x"321b0b",x"2f1a0b",x"371e0d",x"323232",x"5d5d5d",x"3f3f3f",x"373737",x"323232",x"303030",x"3d3d3d",x"545454",x"3a3a3a",x"474747",x"333333",x"333333",x"323232",x"323232",x"3f3f3f",x"363636",x"323232",x"4d4d4d",x"424242",x"3a3a3a",x"363636",x"353535",x"363636",x"383838",x"333333",x"333333",x"636262",x"4e4e4e",x"323232",x"404040",x"585858",x"565656",x"4d4d4d",x"494949",x"494949",x"323232",x"454545",x"474747",x"3e3e3e",x"3f3f3f",x"444444",x"434343",x"474747",x"515151",x"5f5f5e",x"656565",x"656565",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"333333",x"323232",x"323232",x"000000",x"512f16",x"512f16",x"4e2c14",x"331e0e",x"4b2d16",x"442713",x"432712",x"442813",x"442813",x"3f2310",x"402511",x"3c2310",x"3d2310",x"462811",x"3c2210",x"564335",x"422410",x"341d0d",x"381f0e",x"2d190b",x"150e07",x"26160a",x"351e0e",x"1e1208",x"371f0e",x"3b220f",x"402512",x"3e2411",x"3d2310",x"3f2410",x"402410",x"3d220f",x"3c210f",x"381f0e",x"39200f",x"3d2310",x"3d2310",x"402411",x"3c220f",x"3c220f",x"3a210f",x"3d220f",x"422611",x"3f2410",x"3c210f",x"3a200e",x"3e2310",x"422611",x"381f0d",x"381e0d",x"381e0d",x"3b210e",x"3b200e",x"391f0e",x"402410",x"422511",x"432612",x"3f2411",x"3d2210",x"3c210f",x"3f2310",x"3c210f",x"3a200e",x"3c210f",x"3f230f",x"3f2410",x"422510",x"3b210f",x"442713",x"432612",x"442712",x"3c210e",x"3d210e",x"391f0c",x"361d0b",x"42250f",x"3c210d",x"422511",x"3c2210",x"321c0c",x"2d190a",x"2b170a",x"150e07",x"1e1108",x"261509",x"150e07",x"1c1108",x"1c1108",x"2b190b",x"2b190b",x"2f1a0c",x"321c0c",x"331c0c",x"321c0c",x"2d190b",x"2a180a",x"170f07",x"371f0e",x"523f32",x"472915",x"3d2312",x"402512",x"3e2412",x"3a2110",x"3c2110",x"3a2010",x"3b2110",x"3b2110",x"3a2110",x"39200e",x"391f0e",x"3c210f",x"3b210f",x"3c210f",x"371f0e",x"3c210f",x"3c210f",x"3c210f",x"3e220f",x"3c210f",x"3d220f",x"3b200e",x"3c210f",x"422511",x"422611",x"3a220f",x"3d2310",x"371f0d",x"3e2411",x"442713",x"442713",x"442611",x"402510",x"412411",x"3e220f",x"3d220f",x"3e2310",x"3a210f",x"432712",x"3f2410",x"3c220f",x"3f2410",x"3d2310",x"3d2210",x"3d220f",x"432611",x"3d210f",x"3a200e",x"3e220f",x"3f2511",x"3e220f",x"361d0d",x"391f0d",x"3b200e",x"3a200e",x"361d0c",x"412511",x"3d220f",x"37200e",x"412511",x"3f2411",x"3b210f",x"3a200e",x"3c220f",x"39200e",x"3b210f",x"3b210f",x"3e2310",x"3b210f",x"3d230f",x"422612",x"422611",x"432712",x"402410",x"351d0b",x"42240f",x"351d0b",x"3b200d",x"3a200c",x"422511",x"3f2410",x"3f230f",x"3b200e",x"371d0c",x"3a1f0d",x"391e0d",x"331a0b",x"361d0c",x"371c0c",x"361c0c",x"361d0c",x"3a1f0d",x"391f0d",x"361d0c",x"361d0c",x"341c0c",x"3a200e",x"3c210e",x"3b210e",x"3d220f",x"3c210f",x"3d220f",x"3d220f",x"3b210f",x"3a200e",x"361e0d",x"381f0d",x"3a200e",x"391f0d",x"371e0d",x"371f0d",x"3a200f",x"3a200e",x"3a200e",x"3c210f",x"3d220f",x"3a200e",x"3a200e",x"3d220f",x"39200e",x"361f0d",x"3b210e",x"3c210e",x"381f0e",x"3a200e",x"3e2310",x"3b210f",x"412511",x"3c2210",x"3d2210",x"412511",x"3f2511",x"3f2411",x"3d2310",x"3c220f",x"3c220f",x"3a200e",x"39200e",x"3b210f",x"402411",x"402511",x"422611",x"3c220f",x"3a210f",x"38200e",x"402410",x"3e220f",x"432712",x"3d220f",x"3d210f",x"3b210f",x"3d2310",x"3f2310",x"391f0e",x"321c0c",x"371e0d",x"391f0e",x"351d0c",x"3d220f",x"422511",x"442611",x"462813",x"462813",x"3f2410",x"3d220f",x"3f2410",x"3f2210",x"3e220f",x"3d220f",x"3f2310",x"422511",x"412410",x"3f2410",x"442712",x"442812",x"402411",x"472711",x"472711",x"000000",x"000000",x"000000",x"000000",x"391f0e",x"391f0e",x"513728",x"35281f",x"4b4238",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"281e16",x"2a1f17",x"332b24",x"332b24",x"000000",x"000000",x"453326",x"453326",x"4a2b15",x"3a2210",x"351f0e",x"351f0e",x"341d0d",x"361f0e",x"150e07",x"331c0c",x"331d0c",x"2f1b0c",x"2e1a0b",x"2e1a0b",x"341d0d",x"321c0d",x"2f1a0b",x"321c0c",x"331d0d",x"311c0c",x"311c0c",x"2b180b",x"331c0c",x"311c0c",x"331c0d",x"351e0d",x"321d0d",x"331d0d",x"341e0d",x"361f0e",x"311b0c",x"37200f",x"351f0e",x"331d0d",x"2e1b0c",x"321d0d",x"301b0c",x"2a180b",x"2d190b",x"301b0c",x"2a190b",x"311c0d",x"2e1a0c",x"2e1b0c",x"2f1b0c",x"2f1b0c",x"2a180b",x"2f1b0c",x"2e1a0b",x"2a180b",x"2a180b",x"241509",x"1f1209",x"251509",x"221409",x"251509",x"29180b",x"201309",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"492a13",x"492a13",x"150e07",x"150e07",x"22140a",x"54321b",x"54321b",x"463428",x"4b2a14",x"4b2a14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"522e15",x"522e15",x"3a1f0d",x"3f230f",x"3d220f",x"442712",x"422611",x"402511",x"3d210e",x"3d210e",x"371d0c",x"321c0b",x"3b200d",x"373737",x"5e5e5e",x"4f4b48",x"2e2e2e",x"2e2e2e",x"3b3b3b",x"444444",x"3f3f3f",x"323232",x"484848",x"585858",x"414141",x"404040",x"393939",x"3e3e3e",x"494949",x"3e3e3e",x"505050",x"3a3a3a",x"444444",x"000000",x"000000",x"3b3b3b",x"3b3b3b",x"333333",x"313131",x"383838",x"4d4d4d",x"333333",x"444444",x"505050",x"323232",x"323232",x"343434",x"323232",x"323232",x"323232",x"323232",x"3c3c3c",x"4e4e4e",x"4e4e4e",x"4f4f4f",x"505050",x"424242",x"5d5d5d",x"676767",x"676767",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"313131",x"313131",x"313131",x"313131",x"313131",x"000000",x"523016",x"523016",x"4b2913",x"301c0d",x"4d2e16",x"442813",x"412612",x"4a2b15",x"3e2411",x"3f230f",x"3f2410",x"39200f",x"3c220f",x"432410",x"3a210f",x"58483c",x"452712",x"331d0d",x"412410",x"331c0c",x"150e07",x"2a180b",x"341d0d",x"150e07",x"341d0d",x"351d0c",x"391f0e",x"381f0e",x"391f0e",x"3a200e",x"39200e",x"381f0e",x"381f0e",x"351d0d",x"341d0d",x"3b210f",x"3c230f",x"402511",x"402511",x"402511",x"381f0e",x"3a200e",x"3e2310",x"391f0d",x"3e230f",x"3f2310",x"422511",x"3f2410",x"412511",x"3d220f",x"3b200e",x"3a200e",x"3c220f",x"402410",x"402511",x"452813",x"422511",x"412612",x"432712",x"442813",x"3f2410",x"422511",x"452813",x"472914",x"432712",x"472914",x"472914",x"442712",x"452813",x"402410",x"3c200e",x"442610",x"40230e",x"42240f",x"3e220e",x"3f230e",x"42240f",x"412511",x"3e230f",x"321c0c",x"3d220f",x"341d0d",x"150e07",x"231409",x"2e1a0b",x"150e07",x"241509",x"241509",x"2b190b",x"2b190b",x"301b0c",x"321c0c",x"331c0d",x"301b0b",x"301a0b",x"2d190b",x"170f07",x"3c210f",x"4f3f33",x"432714",x"392111",x"3d2312",x"371f0f",x"3b2110",x"392010",x"3f2311",x"3b2111",x"3b2110",x"3a2110",x"3e2310",x"3f2310",x"3c220f",x"3e220f",x"3d220f",x"3c210f",x"3b210f",x"3b210f",x"432611",x"3d210f",x"3f2310",x"3e230f",x"3f2310",x"3e220f",x"3c210f",x"3c210f",x"3d220f",x"381f0e",x"3a210f",x"321c0c",x"3a200e",x"3b210e",x"381f0d",x"3b210e",x"3d220f",x"3b210f",x"371e0d",x"371e0d",x"3f2310",x"3f2410",x"412611",x"432712",x"3f2410",x"412511",x"381e0d",x"3e2310",x"3a200e",x"3f2410",x"3e220f",x"3f2410",x"442712",x"3e2310",x"3c220f",x"3c210f",x"3e220f",x"3f2310",x"402410",x"432611",x"4a2b15",x"412411",x"3f2411",x"402511",x"412511",x"412511",x"3d2210",x"3f2411",x"452913",x"402511",x"452813",x"422712",x"402511",x"402410",x"422511",x"3b200e",x"3a200c",x"311b0b",x"41240f",x"41240f",x"351d0b",x"381e0c",x"402411",x"402411",x"422511",x"3d220f",x"412410",x"412410",x"402310",x"3d220f",x"391f0d",x"3a1f0d",x"361c0c",x"251107",x"241106",x"241106",x"241106",x"251106",x"2a1408",x"331b0b",x"371e0c",x"361c0c",x"331b0b",x"381f0d",x"3a200e",x"381e0d",x"3a200e",x"341d0c",x"351d0c",x"381f0d",x"3a210f",x"3a210f",x"351d0d",x"371e0d",x"3b210e",x"3a200e",x"3e230f",x"3d220f",x"3d220f",x"3d220f",x"3d2310",x"3e230f",x"3d220f",x"3a200e",x"3d220f",x"3b210e",x"3c210f",x"361e0d",x"3c210f",x"3a200e",x"3e2310",x"371f0e",x"3e230f",x"351d0c",x"361e0d",x"371e0d",x"391f0e",x"381f0e",x"371e0d",x"371f0e",x"3a200e",x"2e1a0b",x"381f0e",x"3d2210",x"422611",x"402511",x"3c2310",x"3f2411",x"3b200f",x"3c210f",x"3f2310",x"3c210f",x"3b210f",x"3d2310",x"3f2410",x"402410",x"422611",x"3e220f",x"3c210f",x"3c210f",x"3e230f",x"422511",x"462913",x"452713",x"422611",x"432712",x"482914",x"432712",x"432611",x"402411",x"462814",x"442712",x"442712",x"482a14",x"462914",x"412511",x"3d220f",x"412410",x"41240f",x"472711",x"472711",x"000000",x"000000",x"000000",x"000000",x"361e0c",x"361e0c",x"553a27",x"32251c",x"4a4037",x"150e07",x"150e07",x"150e07",x"150e07",x"1b1008",x"150e07",x"150e07",x"150e07",x"1a1008",x"291d14",x"292018",x"352d26",x"352d26",x"000000",x"000000",x"433226",x"433226",x"4d2d16",x"37200f",x"361f0e",x"341e0e",x"331d0d",x"351e0e",x"150e07",x"341d0d",x"311b0c",x"2e1a0b",x"341d0d",x"301b0c",x"331d0d",x"351e0d",x"311c0c",x"351e0d",x"341d0d",x"351d0d",x"341d0d",x"331c0d",x"341d0d",x"311c0c",x"301b0c",x"351d0d",x"341d0d",x"351e0d",x"2e1a0b",x"341d0d",x"341d0d",x"2d190b",x"2f1a0b",x"2c190b",x"2d190b",x"2e1a0b",x"2d190b",x"2c190b",x"28160a",x"28160a",x"29180b",x"2e1b0c",x"301c0d",x"2f1c0d",x"311c0c",x"311c0d",x"2c180b",x"2d1a0b",x"2a170a",x"2c190b",x"2a180b",x"2c190b",x"28170a",x"28170a",x"211409",x"28170a",x"24150a",x"221409",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2c15",x"4b2c15",x"150e07",x"150e07",x"22140a",x"57341c",x"57341c",x"453226",x"492913",x"492913",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"543117",x"543117",x"3c200e",x"3f2310",x"3e220f",x"412511",x"442813",x"412511",x"3e220e",x"3d210e",x"3d220e",x"251509",x"3b200d",x"373737",x"5f5f5f",x"424141",x"3e3e3e",x"333333",x"2c2c2c",x"3b3b3b",x"333333",x"303030",x"323232",x"323232",x"414141",x"363636",x"3a3a3a",x"363636",x"303030",x"323232",x"333333",x"4f4f4f",x"595959",x"5a5a5a",x"323232",x"363636",x"3b3b3b",x"333333",x"313131",x"313131",x"3f3f3f",x"4d4d4d",x"4e4e4e",x"383838",x"3c3c3c",x"343434",x"343434",x"323333",x"333333",x"313131",x"323232",x"333333",x"333333",x"353535",x"3d3d3d",x"3f3f3f",x"424242",x"4b4b4b",x"656565",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313131",x"323232",x"313131",x"000000",x"512f16",x"512f16",x"4e2d15",x"37200f",x"482a14",x"442814",x"432713",x"442813",x"422612",x"3e2310",x"3d2310",x"3c2310",x"402411",x"442511",x"38200f",x"5c4d42",x"432611",x"2f1a0b",x"3d220f",x"3b210f",x"371f0e",x"311c0c",x"331c0c",x"150e07",x"301b0b",x"341c0c",x"361d0d",x"351c0c",x"331a0b",x"381e0d",x"39200e",x"39200e",x"381f0e",x"361f0e",x"361e0d",x"3a200e",x"3a200e",x"351e0d",x"391f0e",x"3a200e",x"39200e",x"371f0e",x"3a200f",x"341d0d",x"3d220f",x"3f2410",x"3f2411",x"3c2210",x"3f2410",x"402411",x"3f2310",x"3f2410",x"3c220f",x"402411",x"3e2411",x"402410",x"422511",x"402410",x"3f2310",x"3e2310",x"3c210f",x"3f2310",x"3e230f",x"452813",x"432712",x"422611",x"3b200e",x"3f2410",x"381f0d",x"371e0d",x"42250f",x"40240f",x"3b200d",x"381f0c",x"3d220e",x"40230f",x"412410",x"3a1f0e",x"3e2310",x"361f0e",x"3f2410",x"381f0e",x"351d0d",x"301a0b",x"2f190a",x"150e07",x"221309",x"221309",x"2c190b",x"2c190b",x"311c0d",x"331d0d",x"331d0d",x"311c0c",x"2d190b",x"2a180a",x"170f07",x"402410",x"544236",x"4a2c16",x"432814",x"422613",x"3e2312",x"392010",x"3e2311",x"402412",x"442714",x"432814",x"442713",x"452914",x"432813",x"432612",x"432612",x"432511",x"3f2310",x"3b210f",x"3a200e",x"402410",x"412510",x"422510",x"402410",x"402410",x"412410",x"3c210e",x"371e0d",x"361d0d",x"341c0c",x"3a200e",x"371e0c",x"381e0d",x"341b0b",x"341c0c",x"381f0d",x"3b200f",x"39200e",x"3d220f",x"3a210f",x"3c210f",x"3e230f",x"381f0d",x"412410",x"3e220f",x"3e220f",x"3b210f",x"3d220f",x"3f2310",x"3f220f",x"412411",x"402411",x"3c220f",x"3c220f",x"3c220f",x"39200f",x"3e2310",x"422612",x"432612",x"442712",x"462813",x"442712",x"3d220f",x"3a210f",x"3b210f",x"3c210f",x"381f0e",x"39200f",x"3e2411",x"3b2210",x"412611",x"38200e",x"422611",x"3e2310",x"3d220f",x"371d0c",x"3a1f0c",x"40230e",x"371e0c",x"41240f",x"3b200d",x"41240f",x"3f2310",x"402511",x"452812",x"422611",x"422511",x"3e220f",x"3c210e",x"391f0d",x"381d0c",x"381d0c",x"381d0c",x"381e0d",x"381d0c",x"361d0c",x"361d0c",x"371d0c",x"3a200e",x"39200e",x"412511",x"422511",x"3f230f",x"3d220f",x"402411",x"432612",x"412511",x"3b210f",x"3b200f",x"3d220f",x"3e230f",x"3d2310",x"422612",x"412612",x"3f2411",x"432712",x"412512",x"412511",x"432611",x"3e230f",x"3a200e",x"3d220f",x"3d220f",x"3f2310",x"3f2410",x"3d220f",x"3e230f",x"3c220f",x"3e220f",x"3a200e",x"371f0d",x"341c0c",x"371e0d",x"331c0c",x"341c0c",x"331b0b",x"321a0b",x"351d0c",x"361e0d",x"3a200e",x"412410",x"3a210f",x"3a200e",x"3c210f",x"3a200e",x"391f0e",x"3b210f",x"39200e",x"3b210e",x"3e230f",x"3e2310",x"3c210e",x"3e2310",x"402411",x"3c220f",x"3f2310",x"3e2310",x"3f2310",x"422611",x"3f2410",x"412411",x"432712",x"442712",x"442711",x"402411",x"3c210f",x"3f2410",x"3e2310",x"3d210f",x"402411",x"3c220f",x"462913",x"412511",x"3f2411",x"3b210e",x"3f2411",x"381f0d",x"3f220f",x"3f220e",x"452610",x"452610",x"000000",x"000000",x"000000",x"000000",x"3a200e",x"3a200e",x"553825",x"31271e",x"473e35",x"150e07",x"150e07",x"150e07",x"150e07",x"1a1008",x"150e07",x"150e07",x"150e07",x"150e07",x"2c1e15",x"251e18",x"352d25",x"352d25",x"000000",x"000000",x"3e3329",x"3e3329",x"4a2a14",x"3d2411",x"351f0e",x"351e0e",x"321d0d",x"321c0d",x"150e07",x"38200f",x"3b2310",x"3a210f",x"37200f",x"37200f",x"371f0f",x"38200e",x"331d0d",x"351d0d",x"311c0c",x"331c0d",x"321c0d",x"311c0c",x"2f1b0c",x"341d0d",x"321c0d",x"321c0c",x"311c0c",x"2d1a0b",x"2d190b",x"2e190b",x"321b0c",x"2e190b",x"2a170a",x"281609",x"29170a",x"2c190b",x"2d190b",x"2b180b",x"2e1a0c",x"2b180b",x"2a180b",x"2c190b",x"2b180a",x"26160a",x"2b180b",x"2c190b",x"2f1a0c",x"2f1a0c",x"2b190b",x"2e1a0b",x"2f1b0c",x"2a180b",x"28170a",x"241509",x"231509",x"241509",x"27170a",x"1a1008",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4e2d15",x"4e2d15",x"150e07",x"150e07",x"1f1309",x"4b2d18",x"4b2d18",x"413125",x"432611",x"432611",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"533016",x"533016",x"3c200e",x"412410",x"402410",x"432712",x"3a1f0d",x"422511",x"371e0c",x"371e0c",x"361d0c",x"29170a",x"422713",x"4d2c14",x"5b5b5b",x"636363",x"3b3b3b",x"3b3b3b",x"303030",x"333333",x"333333",x"3b3b3b",x"5b5b5b",x"444444",x"404040",x"454545",x"444444",x"454545",x"323232",x"323232",x"3b3b3b",x"505050",x"6b6966",x"6b6966",x"323232",x"323232",x"474747",x"515151",x"2d2e2e",x"494949",x"464646",x"323232",x"4d4d4d",x"5f5f5f",x"615f5e",x"615f5e",x"000000",x"000000",x"000000",x"000000",x"333333",x"313131",x"333333",x"353535",x"3d3d3d",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"313131",x"000000",x"000000",x"000000",x"502e15",x"502e15",x"512f16",x"351f0f",x"4c2d16",x"452813",x"402612",x"422712",x"412512",x"3c2310",x"3a210f",x"3f2511",x"3d220f",x"492812",x"3a210f",x"452812",x"553117",x"482a13",x"331d0d",x"3a210f",x"492913",x"311c0c",x"331d0d",x"3f2410",x"3e220f",x"3d1f0d",x"442510",x"351a0a",x"331909",x"3f210e",x"412410",x"41230f",x"432510",x"3e220f",x"452611",x"422510",x"472712",x"492912",x"482812",x"4c2b14",x"472811",x"462712",x"442611",x"462711",x"4a2b15",x"4c2d15",x"4e2d16",x"4e2d15",x"4f2e16",x"4e2e16",x"502f16",x"502f17",x"502f16",x"4a2a13",x"4e2d16",x"4d2c14",x"502e16",x"4f2d15",x"523017",x"523017",x"523017",x"502f16",x"523018",x"512f17",x"4f2d15",x"4a2a14",x"4c2c14",x"3a1e0c",x"452611",x"41240e",x"46270f",x"44250f",x"3f220d",x"4a2811",x"3f220d",x"4b2911",x"4d2c15",x"522f16",x"452712",x"452712",x"351f0e",x"3d2411",x"472a14",x"2b180b",x"381f0e",x"3f230f",x"522f16",x"522f16",x"2b180b",x"2b180b",x"311c0d",x"341d0d",x"341d0d",x"311b0b",x"2c180a",x"2c180b",x"170f07",x"3f2310",x"4c4036",x"452713",x"412513",x"3e2311",x"412613",x"462914",x"432712",x"442714",x"402513",x"442815",x"3f2411",x"422512",x"3f2311",x"3f2310",x"402410",x"402410",x"3f2410",x"3c2210",x"412411",x"422611",x"452813",x"452812",x"412511",x"452712",x"432611",x"402310",x"412410",x"3f240f",x"3e220f",x"361d0c",x"3b210e",x"361d0c",x"2f1709",x"321a0b",x"3b210e",x"3b200e",x"361d0d",x"321b0b",x"381f0e",x"371e0d",x"381f0e",x"3d220f",x"402410",x"412411",x"422511",x"3e220f",x"432611",x"3a200e",x"452712",x"402512",x"452813",x"412611",x"422612",x"402511",x"412511",x"442713",x"422612",x"412511",x"442712",x"412511",x"442713",x"402511",x"432712",x"452814",x"432713",x"3f2411",x"412612",x"422612",x"3b220f",x"3b210f",x"3e2310",x"361e0d",x"3d220f",x"43250f",x"3b210d",x"40230e",x"371e0c",x"341c0b",x"40230e",x"3e220e",x"412510",x"442712",x"472913",x"432712",x"442712",x"472914",x"452813",x"442611",x"422511",x"432510",x"452812",x"442712",x"432511",x"3f2310",x"3d220f",x"381e0d",x"381d0d",x"3c210f",x"402410",x"3c210e",x"3c210f",x"3e220f",x"3c210e",x"3b200e",x"3c210f",x"3b200e",x"381f0e",x"432612",x"3e2310",x"3d2310",x"402511",x"3e2411",x"402511",x"3d220f",x"3c210f",x"3e2310",x"3c220f",x"3d220f",x"402410",x"432612",x"452812",x"472913",x"462813",x"462813",x"432612",x"3c220f",x"3e2310",x"3b210f",x"3e220f",x"412510",x"3a200e",x"391f0d",x"351d0c",x"341d0c",x"2c1509",x"2b1508",x"331c0c",x"351d0c",x"361e0d",x"3e220f",x"381f0d",x"39200e",x"3d220f",x"3c210f",x"402410",x"3d220f",x"422611",x"3b200e",x"3e2410",x"3d210f",x"3d220f",x"452813",x"442713",x"432612",x"432612",x"412511",x"452813",x"432713",x"462914",x"432612",x"442711",x"472913",x"472813",x"462813",x"3e2410",x"432712",x"442813",x"422612",x"412612",x"452813",x"412612",x"412611",x"412511",x"3f2410",x"371e0d",x"3b210f",x"3c210e",x"381f0d",x"3f220e",x"3f220e",x"000000",x"000000",x"000000",x"000000",x"3d210e",x"3d210e",x"5a3b25",x"2e241c",x"483f36",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"2d1f15",x"261f18",x"3a322a",x"3a322a",x"000000",x"000000",x"3d3329",x"3d3329",x"492913",x"3a2110",x"38210f",x"38200f",x"37200f",x"311b0c",x"150e07",x"371f0f",x"3c2310",x"381f0e",x"351d0d",x"341d0d",x"371f0e",x"341d0d",x"351d0d",x"38200e",x"37200f",x"341e0d",x"39200e",x"351f0e",x"361f0e",x"341e0e",x"38200e",x"311c0c",x"311b0c",x"301b0c",x"2f1b0c",x"2f1a0b",x"28160a",x"301a0c",x"241308",x"201108",x"2a170a",x"29170a",x"261509",x"26160a",x"2c180a",x"2b180b",x"2b180b",x"2b180b",x"29170a",x"2b180b",x"311c0d",x"311c0d",x"2f1b0c",x"2e1a0c",x"2d190b",x"2f1b0c",x"311c0d",x"29170a",x"27170a",x"25150a",x"241509",x"251509",x"1f1309",x"29180b",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4f2d16",x"4f2d16",x"150e07",x"150e07",x"1c1108",x"492c17",x"492c17",x"412f22",x"3f230f",x"3f230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"533117",x"533117",x"391e0c",x"402410",x"3e220f",x"462813",x"412511",x"402410",x"41240f",x"341c0b",x"341c0b",x"2b1a0c",x"3f2411",x"523017",x"3b3b3b",x"353535",x"646464",x"646464",x"595959",x"616161",x"5c5c5c",x"484848",x"414141",x"424242",x"4b4b4b",x"494949",x"454545",x"434343",x"333333",x"313131",x"575757",x"494949",x"686867",x"6b6a68",x"323232",x"2c2c2c",x"3d3d3d",x"575757",x"565656",x"484848",x"464646",x"333333",x"3d3d3d",x"5b5b5b",x"616161",x"616161",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"533116",x"2e1b0c",x"452813",x"472a15",x"412613",x"3e2411",x"3f2411",x"3f2310",x"3d2310",x"3e2310",x"381f0e",x"4b2b13",x"3a210f",x"442812",x"4c2a13",x"4c2b13",x"492912",x"442711",x"492913",x"4a2a13",x"452712",x"482913",x"492913",x"472812",x"4c2b15",x"4d2c14",x"4c2c14",x"492913",x"4c2c14",x"502e16",x"4e2d15",x"462813",x"472812",x"472812",x"452611",x"472912",x"472812",x"412410",x"3e210e",x"3f230f",x"462812",x"472812",x"492a14",x"482913",x"492a14",x"472812",x"442712",x"452712",x"462812",x"442711",x"4c2c15",x"4c2c14",x"4d2c14",x"492913",x"472811",x"482812",x"492a13",x"4b2a13",x"4a2a13",x"4a2913",x"4b2a13",x"343434",x"404040",x"2f2f2f",x"2f2f2f",x"383838",x"3c3c3c",x"3d3d3d",x"482811",x"482812",x"482812",x"482812",x"323232",x"333333",x"323232",x"323232",x"313131",x"333333",x"262626",x"323232",x"312e2c",x"3e220f",x"432510",x"462611",x"343434",x"323232",x"333333",x"2b180b",x"301b0c",x"341d0d",x"321c0c",x"321b0b",x"2b170a",x"2a170a",x"170f07",x"3b200e",x"514034",x"4c2d17",x"442915",x"432714",x"3b2110",x"432712",x"381f0f",x"432613",x"402412",x"432613",x"402512",x"432613",x"412613",x"412511",x"432611",x"3f2410",x"3e2310",x"3f2411",x"3d2310",x"412612",x"3f2410",x"442813",x"3d2310",x"442712",x"3f2410",x"381f0e",x"3c220f",x"402410",x"412511",x"482913",x"3b1f0d",x"3d210e",x"402410",x"3f230f",x"381f0d",x"402410",x"3c220f",x"351d0d",x"381f0e",x"3e220f",x"3c210f",x"381f0d",x"381e0d",x"371d0c",x"351c0b",x"321b0c",x"3b1f0d",x"391e0d",x"3a200d",x"3b200e",x"3a200f",x"321c0c",x"391f0e",x"3d220f",x"3c220f",x"402310",x"381f0e",x"331c0c",x"3a200e",x"361d0d",x"341d0c",x"381f0d",x"3e2310",x"3b200e",x"381f0e",x"361d0c",x"341c0c",x"3b200e",x"3c210f",x"38200e",x"402411",x"3a1f0e",x"3c220f",x"3e220e",x"3d210e",x"3f230e",x"3c210d",x"43250f",x"42240f",x"432611",x"422611",x"391f0d",x"3f230f",x"3b200e",x"3b200e",x"3f2210",x"422410",x"40230f",x"3f220f",x"402310",x"402310",x"3f230f",x"3d220f",x"402310",x"3e220f",x"3e230f",x"39200e",x"412511",x"3e2410",x"3f2410",x"3e220f",x"402410",x"432611",x"452812",x"402411",x"3d220f",x"39200e",x"39200e",x"3d210f",x"381f0e",x"39200e",x"321c0d",x"39210f",x"3b210f",x"402410",x"432711",x"3f2411",x"3e2310",x"422611",x"462813",x"442712",x"3e2411",x"422612",x"422611",x"402411",x"3e2410",x"412511",x"381f0d",x"39200e",x"3d220f",x"3d220f",x"412511",x"351c0c",x"311b0b",x"3a200e",x"3e230f",x"361d0c",x"3d210f",x"402310",x"412410",x"3e220f",x"402410",x"3f230f",x"3a200e",x"381f0d",x"371e0d",x"381e0c",x"381e0c",x"381e0d",x"381e0d",x"371d0c",x"3a200e",x"3b200f",x"341d0c",x"39200e",x"3c210f",x"3b210f",x"3f230f",x"3d220f",x"3b210e",x"3e220f",x"3b200e",x"3a1f0d",x"391f0d",x"3c220f",x"381f0e",x"391f0e",x"371e0d",x"371e0d",x"381f0d",x"3a200e",x"3f2310",x"402310",x"3d2310",x"371e0d",x"381f0c",x"351e0c",x"41240f",x"3d220d",x"3d220d",x"000000",x"000000",x"000000",x"000000",x"3a1f0d",x"3a1f0d",x"5b3d2a",x"2e251d",x"483f36",x"150e07",x"150e07",x"150e07",x"150e07",x"1d1208",x"150e07",x"150e07",x"150e07",x"150e07",x"2b1e14",x"282019",x"3f372e",x"3f372e",x"000000",x"000000",x"41342b",x"41342b",x"452813",x"3a2210",x"38210f",x"392110",x"351f0e",x"331d0d",x"150e07",x"341d0d",x"3a2110",x"38200f",x"3a210f",x"2d1a0b",x"361f0e",x"341d0d",x"371f0e",x"3c2210",x"3a2210",x"341e0e",x"2f1c0c",x"311c0c",x"361f0e",x"341d0d",x"341e0d",x"331c0d",x"301b0b",x"301b0c",x"2f1b0b",x"311c0d",x"321c0d",x"2a170a",x"2a180b",x"2c190b",x"241509",x"221409",x"2a180b",x"2c190b",x"2b180b",x"2a180b",x"2b180b",x"2b180b",x"2a170a",x"2a180a",x"29160a",x"241409",x"2a170a",x"28160a",x"28160a",x"2b180b",x"2d190b",x"26160a",x"27160a",x"26160a",x"231409",x"271609",x"27170a",x"211309",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472913",x"472913",x"150e07",x"150e07",x"221409",x"4e2f1a",x"4e2f1a",x"483326",x"3f230f",x"3f230f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"553117",x"553117",x"381e0c",x"402410",x"412511",x"452813",x"3c210e",x"432712",x"3e2310",x"3d2310",x"3f2410",x"27170a",x"371f0e",x"472711",x"472711",x"474747",x"3e3c3b",x"3f3f3f",x"515151",x"484848",x"393939",x"363636",x"373737",x"424242",x"414141",x"494949",x"000000",x"000000",x"393939",x"393939",x"404040",x"4c4c4c",x"656565",x"646464",x"313131",x"313131",x"323232",x"323232",x"353535",x"353535",x"464646",x"343434",x"343434",x"464646",x"5b5b5b",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"43250f",x"492811",x"462611",x"482913",x"29180b",x"482a14",x"482b15",x"432813",x"3b210f",x"402511",x"3f2411",x"3e2310",x"3d220f",x"39200e",x"4c2c15",x"38200f",x"38200f",x"4c2a13",x"4c2b13",x"492912",x"442711",x"492913",x"4a2a13",x"452712",x"482913",x"492913",x"472812",x"4c2b15",x"4d2c14",x"4c2c14",x"492913",x"4c2c14",x"502e16",x"4e2d15",x"462813",x"472812",x"472812",x"452611",x"472912",x"472812",x"412410",x"3e210e",x"666666",x"626262",x"717171",x"5b5b5b",x"525252",x"492a14",x"472812",x"442712",x"452712",x"462812",x"442711",x"4c2c15",x"4c2c14",x"4d2c14",x"492913",x"472811",x"482812",x"492a13",x"4b2a13",x"323232",x"323232",x"333333",x"333333",x"2e2e2e",x"323232",x"323232",x"333333",x"313131",x"343434",x"3f3f3e",x"3f3f3f",x"303030",x"313131",x"2a2a2a",x"383838",x"4d4d4d",x"313131",x"303030",x"303030",x"2f2f2f",x"313131",x"333333",x"313131",x"313131",x"505050",x"505050",x"333333",x"333333",x"2b190b",x"301b0c",x"331d0d",x"321b0c",x"311b0c",x"2d190b",x"2a170a",x"160f07",x"371e0d",x"564538",x"412512",x"3b2211",x"442814",x"462914",x"422513",x"432712",x"3f2311",x"432712",x"442914",x"3e2411",x"452815",x"3d2210",x"3c210e",x"412511",x"3f2410",x"402410",x"3a210f",x"3c230f",x"3d2310",x"3e2410",x"3f2510",x"3e2310",x"432511",x"412410",x"402410",x"3f2310",x"3f2410",x"412510",x"402310",x"3c210f",x"3c210e",x"381e0d",x"412510",x"3f230f",x"381f0e",x"3c210f",x"371e0d",x"321b0b",x"341d0c",x"341c0c",x"331c0c",x"351d0c",x"351c0c",x"361d0c",x"361d0c",x"391f0d",x"3a1f0d",x"391e0d",x"3a200d",x"391f0e",x"3d220f",x"371e0d",x"361d0c",x"351c0c",x"371e0d",x"391f0d",x"331c0c",x"2d180a",x"321a0b",x"331c0c",x"331c0c",x"351d0c",x"3c210f",x"381f0e",x"3a200e",x"3b200e",x"341c0c",x"361d0c",x"3b200e",x"391f0d",x"3b200e",x"3c220f",x"42240f",x"3c210d",x"41240f",x"3c210d",x"3c210e",x"422511",x"412511",x"402410",x"391f0d",x"3a1f0d",x"3c210e",x"3d210e",x"3b200e",x"371d0c",x"371d0c",x"371c0c",x"371d0c",x"371c0c",x"361c0b",x"341b0b",x"371e0c",x"391f0d",x"391f0d",x"331c0c",x"341d0c",x"361e0d",x"3c210f",x"3a200e",x"3b200d",x"3e220e",x"3c210e",x"3c210e",x"361e0d",x"371d0d",x"422611",x"412410",x"3b200e",x"3e2410",x"3f2410",x"402410",x"422712",x"3c210f",x"492a14",x"412511",x"402410",x"412410",x"412411",x"402411",x"3d2310",x"402511",x"412611",x"422511",x"402410",x"3c210f",x"3d220f",x"3d220f",x"391f0d",x"3b210f",x"3f2310",x"3d220f",x"361d0d",x"361d0c",x"3a200e",x"3d220f",x"3d220f",x"3a200e",x"3d220e",x"391f0d",x"371d0c",x"3d220f",x"381f0d",x"391f0e",x"371d0c",x"361d0c",x"361d0c",x"321b0b",x"391e0d",x"311b0b",x"331c0c",x"39200e",x"381f0e",x"361d0d",x"331c0b",x"361d0c",x"371e0c",x"381f0d",x"381f0d",x"311a0b",x"311a0a",x"351c0c",x"381e0d",x"3a200d",x"3a200e",x"3b200e",x"3a200e",x"3b200e",x"371e0d",x"371d0c",x"381e0d",x"3b210e",x"3d220f",x"422510",x"3a200d",x"3d230c",x"44260f",x"472710",x"472710",x"000000",x"000000",x"000000",x"000000",x"3a1f0f",x"3a1f0f",x"563e2f",x"2a241d",x"4a4239",x"150e07",x"150e07",x"150e07",x"150e07",x"1f1208",x"150e07",x"150e07",x"150e07",x"150e07",x"2d2016",x"2a231c",x"473f35",x"473f35",x"000000",x"000000",x"3d3128",x"3d3128",x"4c2c16",x"36200f",x"3a2210",x"351e0e",x"311c0d",x"311c0c",x"150e07",x"361e0d",x"341e0d",x"371f0e",x"37200f",x"311c0d",x"321c0c",x"321d0d",x"351e0d",x"331d0d",x"311c0c",x"351e0d",x"301c0c",x"331d0d",x"361f0e",x"331d0d",x"331d0d",x"301b0c",x"311b0c",x"2e1a0b",x"2f1b0c",x"331d0d",x"2d190b",x"2a170a",x"2b180a",x"28160a",x"29170a",x"2a180b",x"2a180b",x"2d190b",x"2b180a",x"2b180a",x"2d190b",x"2c190b",x"241509",x"2c180a",x"29170a",x"271609",x"261509",x"29170a",x"2a170a",x"29170a",x"29170a",x"29170a",x"26160a",x"231409",x"211309",x"28160a",x"2b190b",x"27160a",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"150e07",x"150e07",x"221409",x"452a16",x"452a16",x"3f3025",x"42240f",x"42240f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d2b13",x"4d2b13",x"3a1f0d",x"3f230f",x"412411",x"452813",x"3b200e",x"371e0d",x"452712",x"432712",x"3f2410",x"2d1a0b",x"311a0b",x"4a2b14",x"442611",x"472812",x"371e0d",x"472913",x"432510",x"422611",x"462a14",x"452814",x"452813",x"442813",x"472a14",x"492c15",x"472b14",x"412612",x"432713",x"432713",x"452914",x"442813",x"462914",x"462914",x"472a15",x"422713",x"323232",x"323232",x"353535",x"402410",x"3d210e",x"371e0d",x"391f0e",x"3e2310",x"3f2310",x"422511",x"402410",x"432710",x"3f240f",x"3d220e",x"3f2410",x"3d220f",x"3d220f",x"452712",x"3d220f",x"402410",x"3f2410",x"3e2310",x"412411",x"412511",x"412511",x"402410",x"432611",x"3b200e",x"412410",x"3b200e",x"3a200e",x"3b200e",x"3d210f",x"3f2310",x"3f2410",x"432712",x"381f0c",x"492811",x"3b200c",x"492913",x"23150a",x"432713",x"3e2411",x"3a2210",x"3f2310",x"462814",x"432712",x"412511",x"3e230f",x"402410",x"543118",x"422711",x"422711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"6d6d6d",x"6e6d6d",x"666666",x"686159",x"4f4f4f",x"3f3f3f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"323232",x"323232",x"313130",x"383838",x"3f3f3f",x"323232",x"313131",x"323232",x"2f2f2f",x"333333",x"323232",x"3f3f3f",x"302f2e",x"353432",x"333333",x"323232",x"383838",x"000000",x"303030",x"2b2b2b",x"303030",x"2c2d2d",x"313131",x"323232",x"323232",x"626262",x"626262",x"323232",x"323232",x"2a180b",x"2e190b",x"341e0d",x"321c0c",x"311b0c",x"2d180a",x"2a170a",x"160f07",x"381f0d",x"5b483a",x"1a130c",x"19120b",x"19120b",x"17110a",x"2b190d",x"27180c",x"412410",x"442612",x"3b210f",x"422612",x"492a15",x"482a15",x"452712",x"391f0d",x"3f230f",x"3d210f",x"402410",x"412410",x"3d210f",x"3f230f",x"3f2410",x"3d220f",x"412410",x"3f230f",x"422511",x"422510",x"412410",x"412410",x"3f230f",x"3f230f",x"3e220f",x"3f230f",x"3f2410",x"3f230f",x"412410",x"412410",x"422410",x"3f230f",x"412510",x"3e230f",x"412410",x"412511",x"3d220f",x"381e0d",x"3a200e",x"482b15",x"482a14",x"452812",x"432611",x"422410",x"3e230f",x"3a200e",x"3e230f",x"3b200e",x"3d220f",x"361d0c",x"402410",x"3e2310",x"3f2310",x"462813",x"3b200e",x"3f2310",x"412511",x"452712",x"4a2b14",x"452813",x"452812",x"4a2b14",x"472914",x"432612",x"472a14",x"442610",x"442510",x"3c210d",x"3c210d",x"43250f",x"442711",x"422411",x"3e220f",x"452712",x"432510",x"442511",x"432510",x"432410",x"432510",x"432611",x"462711",x"40230f",x"3d200e",x"3e210e",x"3e220e",x"3d210f",x"40240f",x"3a1f0d",x"3a1f0d",x"371d0d",x"351b0b",x"381d0c",x"391d0c",x"3a1e0d",x"40220e",x"452611",x"472812",x"492a14",x"422511",x"472812",x"391f0c",x"42240f",x"3d220e",x"3f230e",x"41240f",x"3d210e",x"482a14",x"482813",x"4a2a14",x"3d220f",x"412410",x"3f230f",x"3d220f",x"3d220f",x"402410",x"432611",x"432611",x"442611",x"402410",x"3b210e",x"3f2410",x"3e230f",x"3f230f",x"3c210e",x"3d210e",x"402410",x"3e220f",x"381e0d",x"3f2310",x"3f230f",x"3f2410",x"3e230f",x"40230f",x"3e220f",x"432511",x"432611",x"442711",x"402410",x"432611",x"3a1e0d",x"3c200d",x"432812",x"462914",x"412612",x"3b210f",x"3c210f",x"3d220f",x"40230f",x"3e220f",x"3f230f",x"41230f",x"3e230f",x"402410",x"412510",x"402410",x"432611",x"3f220f",x"3e220f",x"432511",x"442711",x"482914",x"472913",x"462813",x"482914",x"4b2b15",x"472913",x"442712",x"492a11",x"42260e",x"47290f",x"40240d",x"4a2810",x"4a2810",x"000000",x"000000",x"000000",x"000000",x"3a1f0f",x"3a1f0f",x"5b4130",x"2a231c",x"4c433a",x"150e07",x"150e07",x"150e07",x"150e07",x"1c1108",x"150e07",x"150e07",x"150e07",x"1a1008",x"2d2219",x"332c25",x"4d433a",x"4d433a",x"000000",x"000000",x"3d3128",x"3d3128",x"4b2b14",x"3a2110",x"38200f",x"37200f",x"331d0d",x"2f1a0c",x"150e07",x"321c0b",x"321c0b",x"341d0c",x"321c0c",x"351e0e",x"361f0e",x"301b0b",x"2f1a0b",x"311b0c",x"321c0c",x"321c0d",x"361f0e",x"311c0c",x"361f0e",x"341e0d",x"341d0d",x"2f1a0b",x"2c180b",x"2f1a0b",x"2f1b0c",x"2f1a0b",x"2e1a0b",x"2a180a",x"2a170a",x"2c190b",x"2a180a",x"28160a",x"2a170a",x"2e1a0b",x"2e1a0b",x"2e190b",x"2a180a",x"2e1a0b",x"2f1b0c",x"29170a",x"28160a",x"29170a",x"2f1b0c",x"2f1b0c",x"341e0e",x"2f1b0c",x"2d190b",x"2d1a0c",x"27160a",x"231509",x"241509",x"231409",x"28170b",x"231509",x"1a1008",x"1a1008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2a14",x"4b2a14",x"150e07",x"150e07",x"201309",x"452916",x"452916",x"433024",x"4b2b13",x"4b2b13",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4c2a13",x"4c2a13",x"3e230f",x"402410",x"40230f",x"3c210e",x"402310",x"422511",x"412510",x"3f230f",x"412410",x"3a200e",x"422511",x"40230f",x"472912",x"3d200e",x"371e0d",x"472913",x"432510",x"422611",x"462a14",x"452814",x"452813",x"442813",x"472a14",x"492c15",x"472b14",x"412612",x"432713",x"432713",x"452914",x"442813",x"462914",x"462914",x"472a15",x"422713",x"432611",x"462a14",x"422511",x"402410",x"3d210e",x"371e0d",x"391f0e",x"3e2310",x"3f2310",x"422511",x"402410",x"432710",x"3f240f",x"3d220e",x"3f2410",x"3d220f",x"3d220f",x"452712",x"3d220f",x"402410",x"3f2410",x"3e2310",x"412411",x"412511",x"412511",x"402410",x"432611",x"3b200e",x"412410",x"3b200e",x"3a200e",x"3b200e",x"3d210f",x"3f2310",x"3f2410",x"432712",x"3f230f",x"3e220e",x"391f0d",x"3c210e",x"40230e",x"40230f",x"3e220e",x"3f230e",x"3e220e",x"432712",x"3e2410",x"3d2310",x"40240f",x"432711",x"4a2b13",x"432711",x"432711",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"6a6a6a",x"5d5d5d",x"6e6861",x"6f6963",x"6d6660",x"313131",x"323232",x"535353",x"605e5d",x"5f5d5d",x"575757",x"565656",x"5e5d5c",x"5e5d5c",x"565656",x"5b5a59",x"575757",x"545454",x"545454",x"525252",x"323232",x"3d3a38",x"333333",x"343434",x"3f3f3f",x"5b5a59",x"545454",x"2b2b2b",x"313131",x"2f2f2f",x"303030",x"2f2f2f",x"353432",x"353432",x"333333",x"333333",x"5a5a5a",x"4c4c4c",x"5f5e5d",x"505050",x"303030",x"313131",x"313131",x"313131",x"000000",x"606060",x"606060",x"323232",x"353434",x"29180b",x"2c190b",x"301b0c",x"311b0c",x"331c0c",x"281609",x"27160a",x"160e07",x"3d220f",x"432613",x"4a2c17",x"472a16",x"3d2311",x"3d2412",x"39200f",x"492a15",x"231409",x"150e07",x"150e07",x"150e07",x"3c210f",x"3e230f",x"38200f",x"442813",x"402612",x"422712",x"3c2310",x"412612",x"3f2411",x"39210f",x"3f2411",x"3f2311",x"301b0b",x"381f0e",x"3b2210",x"402511",x"38200f",x"3e2411",x"3c2310",x"392210",x"432713",x"442813",x"3a2110",x"402511",x"412612",x"422612",x"37200e",x"3d2210",x"3f2411",x"38200f",x"412511",x"3d2310",x"361e0d",x"39200e",x"381f0e",x"39200e",x"361f0e",x"3a210f",x"422612",x"3e2411",x"3c230f",x"402511",x"361f0e",x"412511",x"3b2210",x"422612",x"351f0e",x"3b220f",x"3f2410",x"351e0e",x"3e2410",x"3c230f",x"331c0d",x"3f2310",x"3b210f",x"39200e",x"2f1a0b",x"341c0c",x"371f0e",x"1f1208",x"472a14",x"442610",x"442510",x"3c210d",x"3c210d",x"43250f",x"442711",x"422411",x"3e220f",x"452712",x"432510",x"442511",x"432510",x"432410",x"432510",x"432611",x"462711",x"40230f",x"3d200e",x"3e210e",x"3e220e",x"3d210f",x"40240f",x"3a1f0d",x"3a1f0d",x"371d0d",x"351b0b",x"381d0c",x"391d0c",x"3a1e0d",x"40220e",x"452611",x"472812",x"492a14",x"422511",x"472812",x"391f0c",x"42240f",x"3d220e",x"3f230e",x"41240f",x"3d210e",x"482a14",x"482813",x"4a2a14",x"3d220f",x"412410",x"3f230f",x"3d220f",x"3d220f",x"402410",x"432611",x"432611",x"442611",x"402410",x"3b210e",x"3f2410",x"3e230f",x"3f230f",x"3c210e",x"3d210e",x"402410",x"3e220f",x"381e0d",x"3f2310",x"3f230f",x"3f2410",x"3e230f",x"40230f",x"3e220f",x"432511",x"432611",x"442711",x"402410",x"432611",x"3a1e0d",x"3c200d",x"432812",x"462914",x"412612",x"3b210f",x"3c210f",x"3d220f",x"40230f",x"3e220f",x"3f230f",x"41230f",x"3e230f",x"402410",x"412510",x"402410",x"432611",x"3f220f",x"3e220f",x"432511",x"442711",x"482914",x"472913",x"462813",x"482914",x"4b2b15",x"472913",x"442712",x"492a11",x"42260e",x"47290f",x"40240d",x"4a2810",x"4a2810",x"000000",x"000000",x"000000",x"000000",x"3a1f0f",x"3a1f0f",x"583f30",x"2c251e",x"4d443a",x"150e07",x"150e07",x"150e07",x"150e07",x"170f07",x"150e07",x"150e07",x"150e07",x"1c1108",x"382f27",x"473f36",x"51483f",x"51483f",x"000000",x"000000",x"3f332a",x"3f332a",x"4b2b14",x"351e0d",x"371f0e",x"2f1b0c",x"341e0e",x"2d190b",x"150e07",x"2d190b",x"351d0c",x"321c0b",x"2d190a",x"311c0c",x"331d0d",x"341e0d",x"331d0d",x"311c0d",x"321c0c",x"361e0d",x"331d0d",x"351e0d",x"361f0e",x"341d0d",x"331c0d",x"331d0d",x"2e1a0c",x"331d0d",x"331d0d",x"321d0d",x"2f1b0c",x"29170a",x"271509",x"2a170a",x"2d1a0b",x"2d1a0b",x"2e1a0b",x"2f1b0c",x"2f1a0c",x"2e1a0b",x"2d190b",x"2c190b",x"331d0d",x"331c0c",x"2c190b",x"241509",x"311b0c",x"321c0d",x"2d190b",x"2f1b0c",x"2a180a",x"331d0e",x"27170a",x"27170a",x"241409",x"241509",x"221409",x"1a1008",x"160e07",x"160e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d2c15",x"4d2c15",x"150e07",x"150e07",x"1f1309",x"4d2f1a",x"4d2f1a",x"3e3228",x"482812",x"482812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"532f16",x"532f16",x"462711",x"3d210e",x"422510",x"3f220f",x"442712",x"412611",x"3a200e",x"402310",x"422611",x"432711",x"422611",x"38220f",x"3e220f",x"412510",x"3c230f",x"3e210e",x"452813",x"38200f",x"462813",x"432713",x"452914",x"452914",x"452913",x"492b15",x"442914",x"442914",x"412914",x"422712",x"422612",x"412612",x"3f2411",x"402511",x"412712",x"422612",x"452914",x"412612",x"422814",x"381f0e",x"371f0e",x"3b210f",x"3a200e",x"3d2310",x"412612",x"422611",x"412610",x"442812",x"402610",x"402611",x"412512",x"3e2411",x"3f2511",x"402410",x"3b210f",x"3f2410",x"3d2310",x"3b210f",x"3c210f",x"3f2410",x"3e230f",x"3e220f",x"3a200e",x"3d220f",x"3c210f",x"361e0d",x"3a200e",x"321c0b",x"351e0d",x"3d220f",x"3d220f",x"39200e",x"3a200f",x"321c0b",x"311b0b",x"391f0d",x"331b0b",x"331c0b",x"381f0d",x"351d0b",x"3b210d",x"432712",x"402410",x"42250f",x"42270f",x"492b11",x"4e2d14",x"442811",x"442811",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"636362",x"676665",x"686767",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"636363",x"686868",x"6f6862",x"6a635c",x"5f5850",x"323232",x"4a4a4a",x"535353",x"605e5d",x"5f5d5d",x"575757",x"565656",x"5e5d5c",x"5e5d5c",x"565656",x"5b5a59",x"575757",x"545454",x"545454",x"525252",x"585756",x"464646",x"404040",x"3e3e3e",x"4d4c4c",x"5b5a59",x"545454",x"565656",x"444444",x"464646",x"535353",x"535353",x"525252",x"575757",x"5c5c5c",x"565656",x"5a5a5a",x"4c4c4c",x"5f5e5d",x"505050",x"494848",x"333333",x"313131",x"323232",x"000000",x"525252",x"525252",x"4c4742",x"45413e",x"26160a",x"27160a",x"2c190b",x"2a170a",x"301b0c",x"221308",x"1e1208",x"150e07",x"361e0d",x"341d0e",x"4f3019",x"462815",x"402513",x"402512",x"201309",x"201309",x"4d2c14",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"2b190d",x"2b190d",x"58473b",x"493e35",x"51463b",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"4a4138",x"4f453b",x"51483e",x"51483e",x"000000",x"000000",x"42352b",x"42352b",x"4a2a13",x"341d0d",x"38200e",x"361e0d",x"311d0d",x"2e1a0b",x"150e07",x"2a1709",x"341d0c",x"381f0d",x"351d0c",x"361d0c",x"351e0e",x"331d0d",x"2f1a0b",x"321c0d",x"331d0d",x"341e0d",x"341d0d",x"321d0d",x"321d0d",x"341d0d",x"361f0e",x"301b0c",x"2d190b",x"2f1a0b",x"2d190b",x"2a180a",x"2b180b",x"2e1a0b",x"301b0b",x"301b0c",x"341e0d",x"2e1a0c",x"2f1b0c",x"2f1a0b",x"311b0c",x"321c0c",x"311c0c",x"2f1b0c",x"321d0d",x"301b0c",x"311c0c",x"2f1b0c",x"311c0d",x"321e0d",x"2c1a0b",x"2c190b",x"2f1c0c",x"2d1a0c",x"29180b",x"27160a",x"251509",x"1f1208",x"1e1208",x"150e07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4b2b14",x"4b2b14",x"150e07",x"150e07",x"1f1309",x"452a18",x"452a18",x"463429",x"482812",x"482812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"402310",x"432612",x"472a14",x"462813",x"432611",x"472813",x"412511",x"3e220f",x"3e220f",x"3f2410",x"402510",x"412410",x"3e220f",x"462813",x"452813",x"442813",x"39200e",x"412511",x"462b14",x"442d16",x"452b15",x"412a15",x"412a15",x"422813",x"422612",x"422813",x"432813",x"402613",x"412713",x"402612",x"3b2310",x"3e2411",x"3a200f",x"3a210f",x"381f0e",x"3f2511",x"442813",x"402712",x"442913",x"38210f",x"371f0e",x"351e0d",x"422712",x"412711",x"3f2611",x"402610",x"3e250f",x"3d2410",x"3a220f",x"3d2411",x"3a2210",x"361e0e",x"341d0d",x"38200e",x"3c2310",x"3a210f",x"351d0d",x"301a0b",x"321c0c",x"331c0c",x"341d0d",x"39200e",x"3b210e",x"38200f",x"361e0e",x"3a210f",x"3b220f",x"3e2310",x"3d2411",x"351d0d",x"351d0d",x"361f0e",x"321b0b",x"301a0a",x"3c210d",x"3f230f",x"3e220e",x"2f1a0a",x"381f0d",x"3d210e",x"442912",x"492b12",x"4b2c11",x"4e2e12",x"502f12",x"452811",x"452811",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"626261",x"5c5c5c",x"676665",x"646464",x"616161",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5e5c5b",x"5e5c5b",x"746e67",x"675f58",x"635b54",x"605851",x"595148",x"6c655f",x"716b65",x"6b655e",x"706a64",x"706a64",x"746e68",x"756e68",x"726c66",x"736d67",x"6b6661",x"4a4a4a",x"4d4d4d",x"4b4b4b",x"545352",x"5e5851",x"424141",x"313131",x"494949",x"4c4b4b",x"5c5650",x"494541",x"333333",x"313131",x"333333",x"323232",x"323232",x"323232",x"373736",x"3e3d3b",x"43403d",x"4d4741",x"68625b",x"6c665f",x"5c5752",x"4a4948",x"313131",x"323232",x"323232",x"323232",x"5c5c5c",x"5c5c5c",x"333333",x"323232",x"211409",x"241509",x"26160a",x"27160a",x"29170a",x"201208",x"261509",x"150e07",x"3b220f",x"331d0d",x"3b2414",x"3b2414",x"462814",x"241509",x"211309",x"201309",x"2e1a0c",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"2a180b",x"2b190b",x"29180b",x"2d1a0c",x"28170a",x"251509",x"26160a",x"26160a",x"180f08",x"180f07",x"191008",x"170f07",x"190f08",x"191008",x"1c1108",x"1a1008",x"1b1108",x"190f08",x"180f08",x"160e07",x"160e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1c1108",x"1d1108",x"201309",x"1f1209",x"201309",x"211409",x"231409",x"221409",x"231409",x"241509",x"231409",x"211309",x"241409",x"231509",x"241509",x"231409",x"231409",x"231409",x"231409",x"231509",x"221308",x"221308",x"211309",x"221309",x"231409",x"231409",x"241409",x"231409",x"241509",x"241409",x"241509",x"241509",x"231409",x"221409",x"221409",x"241509",x"231409",x"231409",x"221409",x"211309",x"231409",x"221409",x"221409",x"211309",x"22140a",x"221409",x"221409",x"231409",x"221409",x"221409",x"211309",x"221409",x"211409",x"211309",x"201309",x"221409",x"24150a",x"24150a",x"211309",x"221409",x"221409",x"211409",x"221409",x"221409",x"211309",x"221409",x"231409",x"201308",x"221409",x"221409",x"24150a",x"241409",x"241409",x"24150a",x"24150a",x"221409",x"201309",x"231509",x"211309",x"1d1208",x"201309",x"211409",x"211309",x"201309",x"211409",x"211309",x"201409",x"201309",x"3f2411",x"55463a",x"4b4037",x"504539",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"160f08",x"150e07",x"150e07",x"150e07",x"554b41",x"51483e",x"50473d",x"50473d",x"3e220f",x"3c210e",x"44382f",x"44382f",x"472812",x"37200f",x"331d0d",x"331d0d",x"351f0e",x"2f1b0c",x"150e07",x"321c0b",x"361e0d",x"2e1a0a",x"331c0c",x"341d0c",x"38200f",x"351e0d",x"341d0d",x"301b0c",x"341d0d",x"351e0d",x"331d0d",x"321d0d",x"351e0d",x"361f0e",x"361f0e",x"331c0d",x"301b0c",x"29180a",x"321c0d",x"241509",x"2e1a0b",x"29170a",x"2f1a0b",x"361f0f",x"2f1c0d",x"331d0d",x"2c180b",x"301b0c",x"38200f",x"321d0d",x"351e0e",x"321c0d",x"351e0e",x"301b0c",x"2d190b",x"321c0c",x"331d0d",x"311c0c",x"2d1a0b",x"341d0c",x"331e0e",x"2d1a0c",x"29180b",x"27160a",x"231409",x"1f1208",x"27160a",x"27160a",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4a2a14",x"4a2a14",x"150e07",x"150e07",x"1c1108",x"412815",x"412815",x"473629",x"432510",x"432510",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2a13",x"4a2a13",x"3b200e",x"412510",x"492a14",x"452813",x"452812",x"422611",x"422611",x"402410",x"381f0d",x"3b200e",x"3b200e",x"3c210e",x"3b200e",x"3c210f",x"3d210f",x"381e0d",x"3c2310",x"462813",x"492b15",x"442813",x"412612",x"412713",x"432712",x"39200f",x"301a0b",x"2e1a0b",x"311a0b",x"361f0e",x"2e1a0b",x"27160a",x"150e07",x"150e07",x"311c0c",x"28170a",x"251509",x"2c170a",x"281408",x"221208",x"1d1108",x"170f07",x"251609",x"2e1b0c",x"3a220f",x"311d0b",x"311f0a",x"38230c",x"2c1b0a",x"3f240f",x"1e1308",x"37200e",x"181007",x"160e07",x"27170b",x"341e0d",x"361f0e",x"301b0c",x"311b0c",x"2f1b0c",x"231509",x"1d1208",x"29180b",x"39200f",x"38200f",x"351e0e",x"37200f",x"37200f",x"2e1b0c",x"341d0d",x"3c2310",x"38200e",x"3a210f",x"331c0d",x"39210f",x"3a200e",x"321b0b",x"40230e",x"3b210e",x"361e0c",x"41240f",x"462912",x"4c2e13",x"4a2c11",x"4e2e12",x"4b2c11",x"4b2b12",x"422610",x"422610",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"636262",x"616161",x"636261",x"77716b",x"676563",x"505050",x"404040",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"635f5c",x"635f5c",x"5a5147",x"6c645d",x"625951",x"6e6761",x"655e57",x"635c55",x"6d6760",x"6a645d",x"6a635c",x"68615b",x"675f58",x"666059",x"6f6861",x"6b645d",x"69635e",x"484848",x"343434",x"3b3a3a",x"34312e",x"5d554d",x"232222",x"333333",x"525252",x"3c3a37",x"615951",x"434240",x"323232",x"323232",x"393939",x"323232",x"363636",x"2f2f2f",x"31302f",x"44423f",x"504c48",x"59534d",x"605851",x"595149",x"4d4843",x"383736",x"323232",x"333333",x"323232",x"323232",x"686868",x"686868",x"333333",x"333333",x"1d1108",x"1f1208",x"211409",x"1f1208",x"1d1108",x"1b1008",x"160e07",x"150e07",x"3a210f",x"311b0c",x"2b180b",x"2e1a0c",x"372011",x"2e1b0c",x"2f1b0b",x"2e1a0b",x"2e1a0c",x"2d1a0b",x"301b0c",x"2d1a0b",x"2e1a0b",x"2d190b",x"2c190b",x"2c190b",x"2a180b",x"2d190b",x"2c190b",x"2a180b",x"2e1a0c",x"2b190b",x"2b180b",x"2b180b",x"2b170b",x"29170a",x"28160a",x"2b180a",x"28160a",x"28160a",x"29170a",x"27160a",x"27160a",x"27160a",x"28160a",x"28170a",x"28170a",x"28170a",x"28170a",x"2b180b",x"2a180b",x"2c190b",x"2b180b",x"29180b",x"2b180b",x"2a180b",x"2b180b",x"2b180b",x"2d1a0b",x"2b180b",x"29170a",x"2a170b",x"29180a",x"29170a",x"27160a",x"2c180a",x"29170a",x"29170a",x"2a180b",x"2a180a",x"2a180a",x"28170a",x"2b180b",x"29170a",x"2a170b",x"27160a",x"27160a",x"2d1a0b",x"2e1a0b",x"2d1a0b",x"2f1a0b",x"28160a",x"27170a",x"2a180b",x"2b190b",x"29180b",x"2d1a0c",x"28170a",x"251509",x"26160a",x"26160a",x"180f08",x"180f07",x"191008",x"170f07",x"190f08",x"191008",x"1c1108",x"1a1008",x"1b1108",x"190f08",x"180f08",x"160e07",x"160e07",x"160e07",x"170f07",x"180f07",x"1a1008",x"1c1108",x"1d1108",x"201309",x"1f1209",x"201309",x"211409",x"231409",x"221409",x"231409",x"241509",x"231409",x"211309",x"241409",x"231509",x"241509",x"231409",x"231409",x"231409",x"231409",x"231509",x"221308",x"221308",x"211309",x"221309",x"231409",x"231409",x"241409",x"231409",x"241509",x"241409",x"241509",x"241509",x"231409",x"221409",x"221409",x"241509",x"231409",x"231409",x"221409",x"211309",x"231409",x"221409",x"221409",x"211309",x"22140a",x"221409",x"221409",x"231409",x"221409",x"221409",x"211309",x"221409",x"211409",x"211309",x"201309",x"221409",x"24150a",x"24150a",x"211309",x"221409",x"221409",x"211409",x"221409",x"221409",x"211309",x"221409",x"231409",x"201308",x"221409",x"221409",x"24150a",x"241409",x"241409",x"24150a",x"24150a",x"221409",x"201309",x"231509",x"211309",x"1d1208",x"201309",x"211409",x"211309",x"201309",x"211409",x"211309",x"201409",x"201309",x"1f1309",x"201309",x"1f1309",x"28170a",x"2a180b",x"29180b",x"2c190b",x"2b180b",x"2a180b",x"28160a",x"2e1a0b",x"2b170b",x"28170a",x"2b190b",x"2a180b",x"27170a",x"29170a",x"3e220f",x"3c210e",x"42372d",x"42372d",x"462812",x"392110",x"351e0e",x"341d0d",x"331d0d",x"37200f",x"150e07",x"351d0c",x"341d0c",x"321c0b",x"311b0b",x"38210f",x"301b0c",x"351d0d",x"351e0d",x"2d190b",x"311c0c",x"331d0d",x"2c180a",x"2f1a0b",x"341d0d",x"2d190b",x"331c0c",x"301a0c",x"2d190b",x"2a180b",x"29190b",x"301b0c",x"2e1a0b",x"301b0c",x"2f1b0c",x"361f0e",x"2e1a0b",x"311c0d",x"2f1a0c",x"311b0c",x"331d0d",x"331d0d",x"37200f",x"311c0c",x"331d0d",x"311c0c",x"2c190b",x"2a170a",x"2d190b",x"2b180a",x"2c190b",x"2b180a",x"2c180b",x"2b190b",x"28170a",x"231509",x"29170a",x"231409",x"211409",x"1f1309",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482913",x"482913",x"150e07",x"150e07",x"191008",x"472b19",x"472b19",x"44372c",x"422410",x"422410",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"442510",x"442510",x"381f0d",x"3e220f",x"3f220f",x"402410",x"3c210e",x"3b210e",x"3d210f",x"3a200e",x"3b200e",x"40230f",x"3e2310",x"3f2410",x"3f2310",x"412410",x"3c210f",x"3f2310",x"412511",x"412511",x"432611",x"3d2310",x"3f240f",x"3c220f",x"28170b",x"150e07",x"150e07",x"26170a",x"311c0d",x"331d0d",x"38210f",x"1e1209",x"37200f",x"35200f",x"2f1b0c",x"3d2411",x"150e07",x"150e07",x"39200f",x"321d0d",x"150e07",x"150e07",x"301c0d",x"191007",x"35210d",x"412810",x"41260f",x"3b230d",x"3d240e",x"412710",x"251709",x"321d0c",x"1c1208",x"39210f",x"170f07",x"1f1309",x"150e07",x"311b0b",x"150e07",x"331d0d",x"150e07",x"150e07",x"351e0d",x"1d1208",x"150e07",x"39200e",x"3e2310",x"3f2410",x"150e07",x"1e1208",x"191008",x"301b0c",x"39200e",x"3e2310",x"3d2310",x"3b210f",x"39200e",x"442812",x"442811",x"442911",x"482a11",x"4d2e12",x"482a10",x"492b11",x"47290f",x"43270f",x"482911",x"3c210d",x"3c210d",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"616161",x"616161",x"6c655f",x"6d665f",x"645d55",x"383838",x"363636",x"676462",x"605f5e",x"61605f",x"6a6865",x"686663",x"61605e",x"5c5b5a",x"676461",x"666564",x"6d6660",x"5d564e",x"68615a",x"574f46",x"574f45",x"595149",x"574f46",x"5a5249",x"5a5148",x"5c534b",x"5c544c",x"5d544c",x"625a52",x"635b54",x"5a5550",x"333333",x"323232",x"373635",x"46423e",x"5e564d",x"323232",x"2f2f2f",x"323232",x"4a4540",x"5a534b",x"363534",x"323232",x"323232",x"393939",x"313131",x"373737",x"343434",x"484747",x"3e3a36",x"56504b",x"5d564f",x"6e6660",x"544e47",x"47433f",x"333332",x"323232",x"333333",x"323232",x"323232",x"555555",x"555555",x"333333",x"323232",x"221409",x"1f1209",x"180f07",x"160e07",x"311c0d",x"180f07",x"1a1008",x"231509",x"2a180b",x"341d0d",x"221409",x"29170b",x"2e1b0c",x"201309",x"1f1209",x"2c190b",x"2a180b",x"211409",x"24150a",x"29170a",x"2f1c0d",x"221409",x"26160a",x"2a180b",x"29170a",x"2a180a",x"29170a",x"28170a",x"2a180a",x"27160a",x"211308",x"221309",x"28170a",x"2b180a",x"2a180b",x"28160a",x"28160a",x"231509",x"27160a",x"241509",x"231409",x"221409",x"211309",x"221409",x"201308",x"241509",x"251509",x"26160a",x"28170a",x"261509",x"221409",x"251509",x"241509",x"28170a",x"28170a",x"28170a",x"2b190b",x"2a180b",x"27160a",x"28170a",x"231509",x"29180b",x"25160a",x"28170a",x"25150a",x"27170a",x"25150a",x"24150a",x"231509",x"24150a",x"211409",x"1f1309",x"201309",x"231509",x"201309",x"23160a",x"211409",x"26160a",x"221409",x"201309",x"351e0e",x"381f0e",x"3d2310",x"452913",x"422612",x"402511",x"3a2310",x"402611",x"38220f",x"391f0e",x"361e0d",x"3b210f",x"3e2411",x"3f2411",x"442713",x"3e2310",x"412612",x"422611",x"351e0d",x"29170a",x"170f07",x"180f07",x"180f07",x"180f07",x"191008",x"1a1008",x"1c1108",x"1c1108",x"1d1208",x"1e1208",x"1f1209",x"201309",x"211409",x"221409",x"231409",x"25160a",x"25160a",x"25150a",x"25150a",x"25160a",x"25160a",x"25160a",x"25150a",x"25160a",x"26160a",x"241509",x"241509",x"231409",x"241509",x"241509",x"251509",x"251509",x"241509",x"231409",x"231409",x"241509",x"241509",x"231409",x"211409",x"211409",x"221409",x"211309",x"1f1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1c1108",x"1b1008",x"1b1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"1a1008",x"191008",x"191008",x"1a1008",x"1a1008",x"191008",x"191008",x"191008",x"191008",x"191008",x"191008",x"191008",x"1a1008",x"1c1108",x"1d1208",x"1f1309",x"201309",x"23150a",x"25160a",x"25160a",x"28170b",x"28180b",x"29180b",x"28170a",x"29180b",x"2b1a0c",x"2a190b",x"29180b",x"29180b",x"26180b",x"25160a",x"25150a",x"241509",x"241509",x"26160a",x"24160a",x"26160a",x"25160a",x"26160a",x"25160a",x"231509",x"211309",x"201208",x"201309",x"211309",x"201309",x"201309",x"1e1208",x"1c1108",x"1b1108",x"1f1209",x"3d230f",x"3f2410",x"43372d",x"43372d",x"4e2d14",x"38200f",x"311c0d",x"311c0c",x"321c0c",x"38200f",x"150e07",x"37200f",x"38200f",x"341d0d",x"3b220f",x"2e1a0b",x"301a0b",x"351d0d",x"28170a",x"2c190b",x"2d190b",x"2d190b",x"2f1a0b",x"2c180b",x"2b180a",x"2b180a",x"2f1a0b",x"301b0b",x"2c190b",x"27160a",x"2b180a",x"2c190b",x"2d190b",x"2a170a",x"29170a",x"2d190b",x"29170a",x"2c180a",x"2d190b",x"2b180a",x"2e1a0b",x"311c0c",x"2e1a0b",x"2e1a0b",x"2f1a0b",x"2e1a0b",x"2f1a0b",x"2d190b",x"231409",x"311c0c",x"2e1a0c",x"2e1a0c",x"2e1a0b",x"29180b",x"2a180b",x"24150a",x"28170a",x"25150a",x"25160a",x"170f07",x"150e07",x"150e07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"472812",x"472812",x"150e07",x"150e07",x"27160a",x"462a17",x"462a17",x"4b3d32",x"472812",x"472812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4d2c14",x"4d2c14",x"3f2410",x"3c210e",x"3c210e",x"40230f",x"3e220f",x"3e230f",x"412511",x"3c210f",x"3f230f",x"412410",x"3e2310",x"432611",x"412411",x"462813",x"3e220f",x"442712",x"412510",x"452813",x"442713",x"3c2310",x"3d230f",x"402410",x"3f2410",x"452813",x"412611",x"432712",x"150e07",x"150e07",x"3e2511",x"1f1208",x"150e07",x"170f07",x"2b190b",x"150e07",x"402511",x"391f0e",x"361d0d",x"27160a",x"2d1a0b",x"311e0e",x"150e07",x"231509",x"3f2611",x"2c1c09",x"442a11",x"442910",x"4e3013",x"3b240d",x"2a1b09",x"341f0c",x"1d1308",x"311d0c",x"37210f",x"27170b",x"3d230f",x"39200f",x"3e2310",x"150e07",x"29180b",x"201309",x"2a190b",x"150e07",x"38200f",x"150e07",x"150e07",x"3b220f",x"3c210f",x"3e2310",x"3d220f",x"26160a",x"341d0d",x"361f0e",x"3d2310",x"3d2310",x"40240f",x"432611",x"482c12",x"4a2c11",x"4c2d12",x"462810",x"47290f",x"44270e",x"46290f",x"43260f",x"43260f",x"3d220e",x"3d220e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5a5a",x"636261",x"615951",x"716b65",x"5e5750",x"726d68",x"4a4a4a",x"676462",x"605f5e",x"61605f",x"6a6865",x"686663",x"61605e",x"5c5b5a",x"676461",x"706a64",x"5f5f5f",x"4f4f4f",x"545454",x"565656",x"595755",x"4d4d4c",x"3c3c3c",x"434343",x"4a4a4a",x"636262",x"5d5c5b",x"4f4f4f",x"494949",x"434343",x"545454",x"545454",x"565656",x"4e4e4e",x"5a5a5a",x"595959",x"5d5d5c",x"545353",x"585857",x"555453",x"4c4b4b",x"343434",x"333333",x"333333",x"343434",x"333333",x"323232",x"333232",x"484746",x"3f3b36",x"58524d",x"635c55",x"676059",x"5b554e",x"43403c",x"343433",x"333333",x"333333",x"333333",x"000000",x"3f3f3f",x"3f3f3f",x"313131",x"323232",x"27170a",x"221509",x"1a1008",x"160f07",x"2a180b",x"1a1008",x"1c1108",x"1e1208",x"201309",x"231509",x"2b180b",x"231409",x"221409",x"231509",x"24150a",x"26170a",x"231509",x"231409",x"25160a",x"231409",x"231509",x"241509",x"231409",x"231409",x"231409",x"251509",x"241509",x"241409",x"251509",x"27160a",x"27160a",x"27160a",x"27160a",x"27170a",x"27160a",x"26160a",x"26160a",x"26160a",x"26160a",x"251509",x"231409",x"25150a",x"25160a",x"241509",x"27170a",x"25150a",x"241509",x"241409",x"26160a",x"241509",x"27160a",x"26160a",x"26160a",x"27160a",x"27160a",x"28170a",x"28170b",x"26160a",x"26160a",x"241509",x"25160a",x"231509",x"25160a",x"24160a",x"231509",x"231509",x"23150a",x"231509",x"24150a",x"23150a",x"24150a",x"22150a",x"23150a",x"211409",x"1d1108",x"1c1108",x"1a1008",x"191008",x"180f08",x"27170a",x"2b180b",x"2a170a",x"2d190b",x"2d1a0c",x"392311",x"2f1e0e",x"311d0d",x"38200f",x"301d0d",x"2c1a0c",x"311d0d",x"2f1d0d",x"331e0d",x"2e1a0b",x"361e0e",x"351e0e",x"37200e",x"361f0f",x"24150a",x"1d1108",x"1d1108",x"1d1208",x"1d1208",x"1e1209",x"201309",x"211409",x"23150a",x"23150a",x"241509",x"25150a",x"25160a",x"251509",x"27160a",x"28170a",x"28170a",x"2a180b",x"2d1a0c",x"2c1a0c",x"29180b",x"271609",x"29180b",x"28170b",x"29170a",x"29180b",x"251509",x"251509",x"241509",x"27160a",x"261509",x"261509",x"261509",x"28170a",x"29170a",x"29170a",x"29170a",x"29170a",x"28170a",x"26160a",x"26160a",x"25150a",x"241509",x"231409",x"211309",x"211309",x"211309",x"211309",x"201309",x"211409",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1e1208",x"1d1108",x"1d1108",x"1d1108",x"1c1108",x"1d1208",x"1c1108",x"1d1208",x"1c1108",x"1d1208",x"1c1108",x"1d1208",x"1d1209",x"1c1208",x"1c1108",x"1c1108",x"1c1108",x"1d1208",x"1d1208",x"1f1309",x"211409",x"23150a",x"24160a",x"231509",x"231409",x"26160a",x"27160a",x"27170a",x"2d1a0c",x"2b180b",x"29170a",x"29170a",x"29180b",x"2c1b0c",x"2f1e0e",x"301c0d",x"2f1c0d",x"2e1c0d",x"2d1b0c",x"2c1b0c",x"2c1b0c",x"2b190b",x"2a180a",x"2b190b",x"2c190b",x"2b190b",x"2d1a0c",x"2d1a0c",x"2a180b",x"2a190b",x"2a180b",x"29180b",x"28170a",x"27170a",x"25160a",x"231509",x"201309",x"1d1208",x"26160a",x"26160a",x"413328",x"413328",x"4a2a13",x"3a210f",x"361f0e",x"3b220f",x"3a210f",x"3e2411",x"341d0d",x"381f0e",x"35200f",x"301a0b",x"2f1a0b",x"331d0c",x"2f1a0b",x"2d190a",x"2d190b",x"2f1a0b",x"2d190b",x"2e1a0b",x"2c190b",x"2f1b0c",x"2d1a0b",x"321c0c",x"29170a",x"301b0c",x"2f1a0b",x"2f1a0b",x"2d190b",x"2b180b",x"2e1a0b",x"29170a",x"2a170a",x"2b180b",x"2e1a0b",x"2c190b",x"311c0c",x"2d190b",x"2c190b",x"2c180a",x"301b0c",x"2a170a",x"2e1a0c",x"2f1a0c",x"301b0c",x"311c0d",x"321c0c",x"2f1b0c",x"2f1b0c",x"301b0c",x"2f1b0c",x"2b180b",x"2e1b0c",x"2b190b",x"331e0e",x"2f1c0d",x"2b190b",x"201309",x"180f08",x"180f08",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"482812",x"482812",x"150e07",x"150e07",x"29180b",x"432917",x"432917",x"46392e",x"452610",x"452610",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4a2a13",x"4a2a13",x"3e220f",x"3b200e",x"412410",x"40230f",x"3e220f",x"412410",x"3e220f",x"3c210e",x"3e220f",x"422511",x"3f2410",x"442712",x"422611",x"452712",x"402410",x"38200e",x"402410",x"3f230f",x"412410",x"3f230f",x"391f0e",x"39200e",x"321c0d",x"191008",x"331c0c",x"3a1f0d",x"3d220f",x"150e07",x"1c1108",x"2e1a0b",x"3e2411",x"150e07",x"150e07",x"3c230f",x"150e07",x"3d2310",x"150e07",x"25160a",x"3c2411",x"150e07",x"2a190c",x"191007",x"442a13",x"4f3216",x"4b2e13",x"4a2d13",x"4e3013",x"4e3014",x"2f1e0a",x"271909",x"221608",x"201508",x"261709",x"331d0d",x"351f0e",x"191008",x"39210f",x"3e2411",x"321d0d",x"3c2411",x"412612",x"191008",x"38200f",x"331e0e",x"38200f",x"311d0d",x"2b190b",x"1b1108",x"2b190b",x"341e0d",x"351e0e",x"3a210f",x"3f2411",x"3f2410",x"3d230f",x"472913",x"462a11",x"442811",x"4a2c12",x"4d2e14",x"4b2d13",x"4d2e13",x"4d2d13",x"4a2c13",x"502f15",x"452812",x"452812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"4d4d4d",x"4d4d4d",x"5a524a",x"615a54",x"5a534c",x"5c544d",x"615952",x"625b54",x"665f59",x"69635c",x"6b645e",x"6d6660",x"6a635c",x"6a645e",x"6e6861",x"6b645e",x"40403f",x"313131",x"363636",x"363534",x"514a44",x"47423e",x"2c2c2c",x"1b1b1b",x"3b3b3a",x"59544e",x"4e4943",x"333333",x"313131",x"323232",x"333333",x"323232",x"323232",x"333333",x"393736",x"433f3b",x"524c46",x"5c554d",x"595149",x"564f49",x"3d3b39",x"303030",x"323232",x"313131",x"343434",x"333333",x"323232",x"333232",x"484746",x"3f3b36",x"58524d",x"635c55",x"676059",x"5b554e",x"43403c",x"343433",x"333333",x"333333",x"333333",x"000000",x"323232",x"323232",x"323232",x"323232",x"2a190b",x"26170a",x"1c1108",x"2d1a0c",x"2a190b",x"301c0d",x"27170b",x"321d0d",x"331d0d",x"311c0d",x"311c0d",x"39200f",x"2f1b0c",x"2c1a0c",x"29180b",x"28180b",x"28170a",x"27170b",x"2b190b",x"311c0d",x"331d0d",x"2f1c0d",x"321e0e",x"2f1b0d",x"2b190b",x"2a190b",x"2c190b",x"2c1a0c",x"2f1c0d",x"2b190b",x"2c190b",x"2d1a0c",x"2d1a0c",x"2d1a0c",x"2d1a0c",x"29180a",x"2c190b",x"2b190b",x"29170a",x"28160a",x"2c1a0c",x"2c1a0c",x"2c190b",x"29170a",x"29170a",x"2f1a0b",x"2f1a0b",x"361e0d",x"341d0c",x"351d0c",x"381f0d",x"331c0c",x"331c0c",x"361e0d",x"38200e",x"37200e",x"3a220f",x"361f0e",x"361f0e",x"351e0e",x"331d0d",x"341d0d",x"341d0d",x"331d0d",x"311b0c",x"2f1a0b",x"341d0d",x"341e0d",x"311c0d",x"2c180a",x"301b0c",x"321c0c",x"321d0d",x"301b0c",x"2d1a0c",x"36200f",x"311d0e",x"2f1b0c",x"2f1b0c",x"301c0c",x"2f1b0c",x"34200f",x"331e0d",x"3b2311",x"372110",x"372110",x"35200f",x"352210",x"392311",x"35200f",x"331f0e",x"38210f",x"392210",x"38210f",x"3b2210",x"3c2310",x"3c2310",x"3a210f",x"23150a",x"23150a",x"23150a",x"23150a",x"24160a",x"26160a",x"28180b",x"29180b",x"2a190b",x"2b190b",x"2d1a0c",x"2d1a0c",x"2d1a0c",x"2e1b0c",x"2e1b0c",x"2f1c0c",x"2f1b0c",x"2f1b0c",x"311d0d",x"311c0d",x"2f1b0c",x"2f1b0c",x"301c0d",x"2d1a0c",x"2d1a0c",x"2e1a0c",x"2f1c0d",x"2f1c0d",x"2e1b0c",x"2d1a0c",x"2d1a0b",x"2f1c0d",x"2f1b0c",x"2e1a0c",x"2e1a0c",x"2f1b0c",x"2f1b0c",x"2e1b0c",x"2c1a0b",x"2b190b",x"2b190b",x"2b190b",x"28170a",x"26160a",x"28180b",x"28180b",x"27170b",x"25150a",x"231409",x"211309",x"221409",x"231509",x"221409",x"221409",x"221409",x"211409",x"1f1208",x"211309",x"211409",x"211409",x"211409",x"221409",x"211409",x"211409",x"211409",x"201309",x"201209",x"201309",x"201309",x"1f1208",x"1f1208",x"201309",x"221409",x"201309",x"201309",x"231409",x"27160a",x"26160a",x"28170a",x"2b190c",x"2e1b0c",x"2d1a0c",x"2d1a0b",x"2f1b0c",x"2f1b0c",x"301b0c",x"311e0e",x"331e0e",x"37210f",x"36200f",x"33200f",x"34200f",x"342110",x"37200f",x"321d0e",x"331f0e",x"351f0f",x"341f0e",x"331d0d",x"331d0e",x"321d0d",x"311d0d",x"311c0d",x"321d0e",x"311d0d",x"301c0d",x"311c0d",x"2f1c0d",x"2e1b0c",x"2c1a0c",x"29180b",x"26160a",x"23150a",x"2a190b",x"28180b",x"41352b",x"41352b",x"4d2d15",x"3d2310",x"3a200f",x"3b2210",x"3b220f",x"3a2110",x"39200f",x"3a210f",x"3b2210",x"371f0e",x"331d0d",x"39210f",x"382210",x"39210f",x"361f0e",x"351e0e",x"351f0e",x"331d0d",x"321d0d",x"2b190b",x"331d0d",x"351e0e",x"361f0e",x"321c0d",x"341f0e",x"321d0d",x"311c0d",x"301c0c",x"2e1a0b",x"29180a",x"2e1b0c",x"2e1b0c",x"2f1b0c",x"2f1a0b",x"231409",x"331d0d",x"2f1a0b",x"301b0c",x"321c0c",x"2f1a0b",x"301b0c",x"2a170a",x"2f1a0b",x"301b0c",x"341d0d",x"2b190b",x"2e1b0c",x"2c190b",x"311c0d",x"301c0c",x"2d1a0b",x"251509",x"301b0c",x"2a180b",x"2b180b",x"211409",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3e210e",x"3e210e",x"150e07",x"150e07",x"28160a",x"442918",x"442918",x"322a22",x"492912",x"492912",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"482711",x"482711",x"3f230f",x"3d210f",x"3e230f",x"3b200e",x"351d0c",x"391f0d",x"3b210e",x"412410",x"3b200e",x"3c210e",x"3b200e",x"412410",x"3c2310",x"452812",x"422611",x"442813",x"422612",x"452914",x"492b15",x"432611",x"412411",x"3f2410",x"3b2210",x"3d2310",x"361e0d",x"331d0d",x"371f0e",x"3b2310",x"3d2310",x"3b2210",x"2f1b0c",x"29180b",x"29180b",x"2e1b0c",x"38200f",x"341d0d",x"2f1b0c",x"331d0d",x"371f0e",x"1b1108",x"22150a",x"3c2311",x"3e2410",x"321e0c",x"38230c",x"422910",x"40280e",x"4f3014",x"2d1c0a",x"3e2410",x"341e0d",x"2f1b0b",x"2d1a0c",x"3a2210",x"3a2210",x"341d0d",x"311b0c",x"2b190b",x"351d0d",x"241509",x"1e1209",x"301c0d",x"301c0d",x"38200f",x"361f0e",x"38200e",x"3a210f",x"381f0e",x"331c0c",x"341d0d",x"371f0e",x"371f0e",x"3e2310",x"3d2410",x"3f2511",x"402611",x"452811",x"412610",x"442811",x"472a11",x"452910",x"482a11",x"45280f",x"3f230f",x"44260f",x"3d230e",x"3d230e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"606060",x"606060",x"6b655f",x"6f6863",x"726c67",x"6f6a65",x"76716c",x"736e69",x"75706a",x"6f6963",x"6e6862",x"766f6a",x"746e68",x"746e68",x"756f6a",x"756e69",x"414141",x"323232",x"323232",x"3c3a38",x"564f47",x"3e3c39",x"292929",x"575757",x"373533",x"5c554e",x"615f5d",x"545454",x"373737",x"333333",x"313131",x"2d2d2d",x"343434",x"333332",x"3d3b38",x"45403b",x"554e47",x"5d554d",x"575048",x"4c4742",x"373634",x"313131",x"323232",x"333333",x"333333",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"383838",x"383838",x"323232",x"323232",x"29170b",x"25150a",x"25160a",x"27160a",x"2c190c",x"2e1b0c",x"341e0e",x"321c0d",x"301b0c",x"311b0c",x"331c0d",x"2f1a0c",x"331d0d",x"351e0e",x"2d1a0c",x"37200f",x"311c0d",x"38200f",x"37200e",x"311c0d",x"321d0d",x"351e0d",x"331d0d",x"321c0c",x"2d190b",x"2c180b",x"2e190b",x"2d190b",x"271609",x"27160a",x"2d190b",x"2c180a",x"2c190b",x"2f1a0b",x"301b0c",x"2d190b",x"29170a",x"28160a",x"27160a",x"28170a",x"261509",x"27160a",x"2c180b",x"28160a",x"2d190b",x"321c0c",x"331c0c",x"361e0d",x"321c0c",x"331c0c",x"331c0c",x"381f0e",x"371f0d",x"321b0b",x"341c0c",x"361d0d",x"3a200f",x"3b2210",x"3a210f",x"3a210f",x"3a210f",x"37200f",x"3a2210",x"38210f",x"351e0e",x"351e0d",x"39200e",x"392110",x"341e0e",x"331c0c",x"311c0c",x"321d0d",x"38210f",x"331e0e",x"321d0d",x"2b180b",x"321c0d",x"2d1a0b",x"301c0d",x"351e0e",x"2e1a0c",x"341e0d",x"351e0e",x"321d0d",x"331e0e",x"392210",x"382110",x"321d0d",x"361f0e",x"35200f",x"372110",x"392210",x"3b2310",x"37200f",x"3b2210",x"381f0e",x"3a210f",x"3c2310",x"3d2411",x"3a2210",x"331d0d",x"351e0d",x"311c0c",x"361e0d",x"2a180b",x"2c190b",x"2e1b0c",x"2f1b0c",x"301c0d",x"331c0d",x"321c0c",x"331d0d",x"311c0c",x"361d0d",x"361e0d",x"361f0d",x"381f0e",x"38200f",x"38210f",x"37200f",x"37200e",x"351f0e",x"331d0d",x"331d0d",x"331d0d",x"301b0c",x"2f1a0b",x"2e190b",x"2d190b",x"2d190b",x"2d190b",x"2d190a",x"2c180a",x"2d190b",x"2d190b",x"2e1a0b",x"301b0c",x"2f1a0b",x"2e190b",x"2e190b",x"2d190b",x"2d190b",x"2c180a",x"2b180a",x"2d190b",x"2d180a",x"2b180a",x"301b0c",x"2e190b",x"2f1b0c",x"2f1a0b",x"2a170a",x"2b170a",x"2e190b",x"301b0c",x"2b180b",x"2c180b",x"2c190b",x"2d190b",x"311d0d",x"311d0d",x"321d0d",x"321d0d",x"351f0e",x"321d0d",x"301c0d",x"2f1b0c",x"2c190b",x"2f1b0c",x"311c0d",x"311c0d",x"2c190b",x"321c0c",x"2d1a0c",x"37200f",x"392110",x"341e0e",x"361f0e",x"351e0e",x"36200e",x"37200f",x"351f0e",x"39200f",x"39200e",x"3a210f",x"3b210f",x"3d2310",x"412612",x"402612",x"3e2411",x"3c2210",x"412612",x"412612",x"422813",x"442813",x"3e2411",x"3e2411",x"321c0d",x"331d0d",x"331d0d",x"36200f",x"3a2210",x"331d0d",x"341d0d",x"361e0d",x"371e0d",x"351e0d",x"38200f",x"361f0e",x"39210f",x"37200e",x"211409",x"221409",x"45382e",x"45382e",x"462711",x"381f0e",x"371f0e",x"39200f",x"3a210f",x"36200e",x"39210f",x"3a2210",x"39200f",x"351f0e",x"361f0e",x"361f0e",x"331d0d",x"301b0c",x"2d190b",x"2d190b",x"2e190b",x"2e190b",x"2b180a",x"2c180a",x"311b0c",x"251509",x"2e190b",x"2b180b",x"2d190b",x"2c190b",x"2c180b",x"221409",x"28160a",x"2b180a",x"29170a",x"27160a",x"27160a",x"2a170a",x"27160a",x"2c190b",x"301b0c",x"2f1b0c",x"2c180a",x"2d190b",x"28160a",x"321c0c",x"2e1a0b",x"2b180a",x"2a170a",x"2a180a",x"2c1a0b",x"321d0d",x"311c0d",x"2c1a0c",x"311c0d",x"2f1b0d",x"311d0d",x"311d0d",x"29180b",x"1e1208",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3c200e",x"3c200e",x"150e07",x"150e07",x"24160a",x"402717",x"402717",x"3c2e24",x"482812",x"482812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"4e2c15",x"4e2c15",x"412511",x"462913",x"472913",x"432611",x"432611",x"442712",x"3a210f",x"361f0e",x"391f0e",x"391f0d",x"442712",x"472914",x"462914",x"462914",x"472a14",x"462813",x"422611",x"3b220f",x"3d220f",x"3e2310",x"402410",x"422611",x"3e2310",x"3e2310",x"3a210f",x"3d230f",x"412511",x"402511",x"3a210f",x"3e2410",x"371f0e",x"321b0c",x"271408",x"321c0c",x"3a200f",x"3d2310",x"3b210f",x"3b220f",x"3a200e",x"38200e",x"3a2210",x"3f2512",x"3d2310",x"412610",x"462a12",x"452910",x"482c12",x"452a11",x"402510",x"432711",x"412611",x"3a210e",x"3e2410",x"422712",x"422611",x"38210f",x"351d0d",x"3c220f",x"3d230f",x"38200e",x"361f0d",x"39200e",x"37200f",x"39200f",x"38200f",x"3c2310",x"3e2410",x"3a210f",x"3d2310",x"38200e",x"38200f",x"38200e",x"321c0c",x"3d220f",x"3e230f",x"432611",x"3f250f",x"3a210e",x"3e230f",x"41260f",x"452810",x"422710",x"472911",x"44270f",x"4b2b12",x"40240f",x"40240f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"5a5856",x"5a5856",x"6d6660",x"615951",x"615a53",x"69635c",x"756f69",x"746e69",x"726b65",x"746e69",x"716b65",x"706a63",x"746e69",x"76706b",x"726c66",x"6e6964",x"5d5d5d",x"373737",x"363635",x"474441",x"605851",x"383735",x"333333",x"393939",x"3e3b37",x"5b544c",x"555452",x"535352",x"4d4d4d",x"323232",x"333333",x"323232",x"333333",x"363535",x"3f3c39",x"4e4943",x"5a544c",x"5d564e",x"5a534c",x"484440",x"373636",x"333333",x"323232",x"323232",x"323232",x"3c3c3c",x"3a3a3a",x"323232",x"323232",x"323232",x"323232",x"414141",x"313131",x"323232",x"363636",x"363636",x"343434",x"2f2f2f",x"2f2f2f",x"2e2e2e",x"383838",x"383838",x"313131",x"333232",x"2a190b",x"25150a",x"211409",x"2a180b",x"2f1c0d",x"321d0d",x"351e0e",x"341e0e",x"361f0e",x"37200e",x"341e0e",x"321d0d",x"321c0d",x"39200f",x"351e0d",x"361f0e",x"361e0e",x"39210f",x"341e0d",x"301c0c",x"2f1a0b",x"331c0c",x"351d0d",x"321c0d",x"311b0c",x"2f1a0b",x"301a0b",x"2d190b",x"29170a",x"29170a",x"321c0c",x"331c0c",x"351e0d",x"331c0d",x"341d0d",x"301c0c",x"2e1a0c",x"2d190b",x"2d1a0c",x"2a180b",x"29170a",x"29170a",x"2c190b",x"2d1a0b",x"321d0d",x"361f0e",x"3d2311",x"3c2210",x"3c2210",x"3c2210",x"3f2411",x"3b210f",x"3d220f",x"351d0d",x"371e0d",x"3d2310",x"3d2311",x"3c2311",x"3e2411",x"3d2411",x"39200f",x"371f0e",x"351e0e",x"331d0d",x"331d0d",x"361e0d",x"3a2110",x"38200e",x"38200e",x"351e0d",x"2f1b0c",x"36200f",x"361f0e",x"321c0d",x"351e0e",x"311c0c",x"291609",x"241308",x"2b180b",x"2c190b",x"341e0d",x"351e0e",x"331d0d",x"2e1a0b",x"29180b",x"36200f",x"35200f",x"351e0e",x"361f0e",x"37200f",x"351e0d",x"36200f",x"38200f",x"361f0e",x"3b2210",x"39200f",x"351d0d",x"3a210f",x"3d2310",x"3f2511",x"39200f",x"361e0d",x"311c0c",x"2f1b0c",x"2c190b",x"2d1a0b",x"301c0c",x"321c0d",x"341e0e",x"351f0e",x"38200f",x"3a210f",x"39210f",x"37200e",x"39200f",x"3a210f",x"371f0d",x"371f0e",x"361f0e",x"361e0e",x"351e0e",x"361f0e",x"331c0d",x"301b0c",x"2f1a0c",x"311c0c",x"301b0c",x"2f1a0c",x"2d190b",x"2e190b",x"2f1a0b",x"2f1a0b",x"311b0c",x"311b0c",x"331d0d",x"321c0c",x"321c0c",x"321c0d",x"341e0d",x"341e0e",x"341e0e",x"331d0d",x"311b0c",x"311b0c",x"2f1a0b",x"311b0c",x"321c0d",x"351e0e",x"351f0e",x"351f0e",x"331d0d",x"311c0d",x"321d0d",x"341e0d",x"351e0d",x"301b0c",x"2b170a",x"311c0c",x"321c0d",x"321e0e",x"341e0e",x"361f0e",x"37200f",x"311c0d",x"321d0d",x"2c180b",x"2d1a0c",x"2d190b",x"2c190b",x"351f0e",x"311c0d",x"331d0d",x"311c0c",x"301c0d",x"351f0e",x"351f0e",x"37200f",x"301b0c",x"341d0d",x"271408",x"331c0c",x"331d0d",x"3b210f",x"39200f",x"3a210f",x"38200e",x"371f0e",x"3e2411",x"3e2411",x"3d2310",x"3c2210",x"3e2411",x"3d2310",x"402612",x"3e2411",x"39210f",x"3e2411",x"361f0f",x"2f1a0b",x"351f0e",x"351f0e",x"341e0e",x"39210f",x"361e0d",x"381f0e",x"361e0e",x"371f0e",x"361e0e",x"371f0e",x"3b220f",x"361f0e",x"23150a",x"23150a",x"4b3c31",x"4b3c31",x"492a13",x"3b2210",x"38200f",x"351e0d",x"2f1b0b",x"321d0d",x"3b220f",x"38200f",x"361f0e",x"331d0d",x"321c0c",x"2f1a0b",x"351d0d",x"351e0d",x"331c0c",x"2e1a0b",x"28170a",x"2b180a",x"2d190b",x"311b0c",x"2f1a0b",x"2d190b",x"2a190b",x"2f1b0c",x"2e1a0b",x"2e1a0b",x"2d1a0b",x"331d0d",x"2e1a0c",x"241509",x"301a0b",x"2a170a",x"2c190b",x"2f1b0c",x"2d1a0b",x"2e1a0c",x"321d0d",x"2f1b0c",x"351e0e",x"301c0d",x"311d0d",x"2f1b0c",x"321d0d",x"271609",x"2e1a0b",x"2f1b0c",x"2e1b0c",x"321d0d",x"341e0e",x"311d0d",x"2c1a0b",x"29180b",x"28170a",x"2e1b0c",x"2b180b",x"29180b",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"341a0b",x"341a0b",x"150e07",x"150e07",x"28170a",x"4f3e32",x"4f3e32",x"473224",x"482812",x"482812",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"492913",x"492913",x"422611",x"452712",x"422611",x"3f2410",x"3a200e",x"381e0d",x"3c210e",x"341d0d",x"3e230f",x"3a200e",x"3b200e",x"432511",x"3a200d",x"3d220f",x"3d220f",x"402411",x"442712",x"3e2310",x"3c210f",x"3d220f",x"3f2310",x"3b210f",x"3c220f",x"39200e",x"3a200e",x"371e0d",x"381f0d",x"341d0c",x"38200e",x"3b210f",x"3e2310",x"3e2411",x"3b2210",x"381f0e",x"331c0d",x"3a210f",x"3f2410",x"3f2411",x"402511",x"412512",x"412612",x"3c220f",x"39200e",x"3b210f",x"3f250f",x"422711",x"402511",x"412611",x"402410",x"462912",x"422711",x"412610",x"40250f",x"452911",x"482a13",x"442812",x"3c230f",x"39200e",x"3c220f",x"381f0e",x"3a210d",x"39200e",x"38210e",x"3a220f",x"351e0e",x"3c220f",x"402511",x"442813",x"3b2210",x"39200f",x"3a2210",x"3b2210",x"361e0d",x"391f0d",x"3e230f",x"432711",x"3e240f",x"40260f",x"412610",x"40250f",x"40260e",x"44280f",x"43280e",x"3d220d",x"41230e",x"3c220e",x"3c220e",x"331d0e",x"37200f",x"2e1b0c",x"2f1b0c",x"341e0d",x"341d0d",x"2e1a0c",x"2d1a0b",x"311c0d",x"5a5856",x"5a5856",x"6d6660",x"615951",x"615a53",x"69635c",x"756f69",x"746e69",x"726b65",x"746e69",x"716b65",x"706a63",x"746e69",x"76706b",x"726c66",x"6e6964",x"5d5d5d",x"373737",x"363635",x"474441",x"605851",x"383735",x"333333",x"393939",x"3e3b37",x"5b544c",x"555452",x"2f2f2f",x"313131",x"323232",x"606060",x"595958",x"5b5a5a",x"545454",x"626262",x"686665",x"686562",x"625f5d",x"353535",x"454545",x"3a3a3a",x"353535",x"3b3b3b",x"3b3b3b",x"363636",x"3c3c3c",x"3a3a3a",x"323232",x"323232",x"323232",x"323232",x"414141",x"313131",x"323232",x"363636",x"363636",x"343434",x"2f2f2f",x"2f2f2f",x"2e2e2e",x"333333",x"333333",x"323232",x"343434",x"29180b",x"241509",x"1e1208",x"25160a",x"301c0c",x"341f0e",x"331d0e",x"311c0d",x"331d0d",x"37200f",x"36200e",x"331e0e",x"2e1b0c",x"39210f",x"2c180b",x"301b0b",x"301a0b",x"3a210f",x"361f0e",x"2e1a0c",x"2c1a0b",x"341d0d",x"311b0c",x"2b180a",x"2a180a",x"2d190b",x"2a160a",x"2c180a",x"2b180b",x"2a180b",x"331d0d",x"341d0d",x"311b0c",x"2f1a0b",x"2e190b",x"29170a",x"271609",x"271609",x"27160a",x"28160a",x"29170a",x"29170a",x"301b0c",x"2d190b",x"321d0d",x"351e0d",x"39210f",x"39200e",x"391f0e",x"361d0d",x"331c0c",x"361f0d",x"3b210f",x"3b200e",x"351d0d",x"341d0d",x"38200e",x"351d0d",x"381f0e",x"38200e",x"371f0e",x"371f0e",x"361e0d",x"361f0d",x"351e0d",x"361f0e",x"361e0e",x"351e0d",x"351e0d",x"331d0d",x"301b0b",x"2e190b",x"2e190b",x"311c0c",x"321c0d",x"331d0d",x"38200f",x"331d0d",x"2e1a0b",x"301b0c",x"2d1a0c",x"361f0e",x"361f0e",x"3c2210",x"341e0e",x"331e0e",x"301b0c",x"331d0d",x"321c0d",x"351e0e",x"331d0e",x"361f0f",x"38210f",x"3a210f",x"38200f",x"39200f",x"39200f",x"3c220f",x"3c2210",x"3d2311",x"3d2310",x"3a210f",x"3a210e",x"321c0c",x"2c190b",x"2d1a0b",x"301c0c",x"331e0e",x"39210f",x"361f0e",x"39200f",x"3a220f",x"3c2310",x"3a220f",x"38200f",x"3a2210",x"371f0e",x"321c0c",x"321b0c",x"351e0e",x"371f0e",x"361f0e",x"361f0e",x"331d0d",x"301a0c",x"2d190b",x"2e190b",x"2d180b",x"2b170a",x"2b170a",x"2d190b",x"311b0c",x"331d0d",x"331d0d",x"321c0c",x"2f1a0b",x"2f1a0b",x"2c180a",x"2c180a",x"2d190b",x"2e190b",x"2e190b",x"2f1a0b",x"301b0b",x"321c0c",x"331d0d",x"341e0d",x"341e0d",x"361f0e",x"361f0e",x"321c0c",x"2e190b",x"2d190b",x"2c180b",x"311c0c",x"321c0d",x"2f1b0b",x"2c190b",x"2c190b",x"29170a",x"2d1a0b",x"311c0c",x"321c0d",x"37200e",x"2f1a0c",x"2f1a0c",x"311c0c",x"311c0c",x"311c0c",x"321c0c",x"301b0c",x"2f1b0c",x"2d190b",x"2d190a",x"2c180a",x"301b0c",x"301b0c",x"351e0e",x"361f0e",x"351f0e",x"321c0d",x"301b0c",x"351e0d",x"38200f",x"3a210f",x"3b2210",x"3e2411",x"3d2411",x"3b210f",x"381f0e",x"3a200f",x"3c220f",x"3d2310",x"412512",x"3e2410",x"402511",x"3f2411",x"341e0e",x"331d0d",x"321d0d",x"341e0d",x"361f0e",x"351f0e",x"39210f",x"38200e",x"38200e",x"351d0d",x"381f0d",x"361e0d",x"39200f",x"37200f",x"23150a",x"23150a",x"48392e",x"48392e",x"4c2d16",x"3b2210",x"3b2310",x"3a210f",x"301a0b",x"2e1a0b",x"311c0c",x"361f0e",x"311c0c",x"361f0e",x"3a210f",x"2f1a0c",x"321c0c",x"301a0b",x"311b0c",x"2d190a",x"28150a",x"311a0b",x"311b0c",x"321c0d",x"331d0d",x"2e1a0b",x"2b180b",x"27160a",x"29170a",x"28160a",x"261509",x"261509",x"2a170a",x"2a180a",x"2c190b",x"29170a",x"29180b",x"2d1a0b",x"2e1b0c",x"311c0c",x"2f1b0c",x"2e1a0c",x"2e1a0b",x"29170a",x"2a170a",x"2d1a0b",x"311b0c",x"2b180b",x"2a170a",x"29170a",x"2b180b",x"29170a",x"2c180b",x"2c190b",x"2b190b",x"2b190b",x"29170a",x"2b190b",x"29170a",x"1f1309",x"170f07",x"170f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"371e0c",x"371e0c",x"150e07",x"150e07",x"221409",x"43352b",x"43352b",x"30271e",x"4d2b14",x"4d2b14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"412411",x"412411",x"543218",x"5a351a",x"573318",x"553119",x"512f16",x"4d2b14",x"4d2b14",x"4e2b14",x"533016",x"4a2a12",x"502d15",x"542f16",x"522e16",x"482812",x"512e15",x"4f2b15",x"4e2c14",x"4c2a14",x"462711",x"4c2b14",x"512d15",x"553117",x"533017",x"513018",x"563219",x"543118",x"522f16",x"4e2c14",x"4f2c14",x"4a2912",x"4c2a13",x"492912",x"4c2a13",x"482711",x"442511",x"462711",x"4c2b14",x"4a2912",x"462611",x"3f200e",x"41220e",x"462711",x"462711",x"4d2b14",x"502e16",x"4f2d15",x"4d2b14",x"4b2b13",x"4a2a13",x"44260f",x"492911",x"502e14",x"502e15",x"4d2c14",x"513015",x"4b2b13",x"502d14",x"472811",x"472711",x"40230f",x"442610",x"4a2911",x"4a2912",x"4a2a12",x"452712",x"4a2b13",x"4f2d15",x"4f2d14",x"4d2b14",x"472711",x"482811",x"492812",x"472711",x"4d2c14",x"482913",x"4e2e15",x"513016",x"492b13",x"4b2c13",x"4e2e14",x"4a2b12",x"502e13",x"4b2b11",x"4d2b12",x"4c2a11",x"492811",x"311c0d",x"331d0e",x"37200f",x"2e1b0c",x"2f1b0c",x"341e0d",x"341d0d",x"2e1a0c",x"2d1a0b",x"311c0d",x"321d0d",x"2c190b",x"2d1a0c",x"331d0d",x"2b180b",x"2c190b",x"2d1a0c",x"321d0d",x"2f1c0d",x"2f1c0d",x"2f1b0c",x"412612",x"361f0e",x"2c190b",x"301b0c",x"341d0d",x"341d0d",x"311b0b",x"321c0c",x"371f0e",x"311c0c",x"29160a",x"150e07",x"26160a",x"482913",x"482913",x"323232",x"323232",x"2d2d2d",x"323232",x"393939",x"515151",x"505050",x"454545",x"353535",x"353535",x"343434",x"3a3a3a",x"3a3a3a",x"3c3c3c",x"404040",x"3f3f3f",x"3e3e3e",x"3f3f3f",x"414141",x"424242",x"454545",x"383838",x"323232",x"343434",x"323232",x"3b3b3b",x"404040",x"414141",x"414141",x"323232",x"424242",x"434343",x"444444",x"353535",x"32302f",x"343434",x"323232",x"323232",x"28170a",x"221409",x"190f07",x"241509",x"2c190b",x"321c0c",x"29180b",x"2c190b",x"2d190b",x"321d0d",x"351e0e",x"2c190b",x"2f1b0c",x"2f1a0b",x"2c180b",x"2f1b0c",x"2f1b0c",x"2c1a0c",x"2a190b",x"321d0d",x"301c0c",x"341d0d",x"301b0c",x"311c0d",x"2e1a0b",x"2a170a",x"2d190b",x"261509",x"2c190b",x"2d190b",x"2e1a0b",x"2b180a",x"2a170a",x"2b170a",x"2d190b",x"2c190b",x"27160a",x"261509",x"26150a",x"28170a",x"28160a",x"29170a",x"311b0c",x"2c190b",x"341e0e",x"3b2210",x"3e2511",x"412612",x"3d2310",x"3d2310",x"3c220f",x"381f0e",x"3a200f",x"3d2310",x"3a200e",x"3c2210",x"3c220f",x"39200e",x"3a210f",x"39200f",x"361e0d",x"381f0e",x"361e0d",x"331c0d",x"341d0d",x"361f0e",x"38200f",x"38200f",x"3d2311",x"38200f",x"39210f",x"37200e",x"311c0c",x"321c0c",x"2e1a0b",x"2f1a0b",x"321c0c",x"2b180b",x"2d190b",x"2e190b",x"2f1a0c",x"321c0c",x"2e1a0b",x"2c180a",x"2a160a",x"2d180a",x"2d190b",x"301b0c",x"321d0d",x"351e0e",x"351e0e",x"331c0d",x"361e0e",x"351e0d",x"331c0c",x"321c0c",x"39200e",x"3b220f",x"371f0e",x"3b220f",x"381f0e",x"38200e",x"371f0d",x"351e0d",x"2a170a",x"29170a",x"2d190b",x"301b0c",x"341e0d",x"331d0d",x"351e0d",x"38200e",x"38200e",x"371f0e",x"331c0d",x"361e0d",x"361e0d",x"371e0d",x"37200e",x"39200f",x"3a220f",x"38210f",x"37200f",x"351e0e",x"351e0d",x"341d0d",x"331c0d",x"2e1a0b",x"301b0b",x"2e190b",x"2e1a0b",x"301b0c",x"321c0c",x"301b0c",x"2b170a",x"2c180a",x"2d190a",x"311b0c",x"311b0c",x"2f1a0b",x"2e190b",x"2f1a0b",x"2e190b",x"311b0c",x"331d0d",x"311b0c",x"351e0d",x"3a220f",x"37200f",x"3b2310",x"36200f",x"37200e",x"361f0e",x"331c0c",x"301b0c",x"311c0d",x"341d0d",x"361e0e",x"341d0d",x"311c0c",x"2e1a0c",x"341e0d",x"331d0d",x"351e0d",x"321c0c",x"311b0c",x"321c0c",x"311c0c",x"311c0d",x"39210f",x"321d0d",x"351e0e",x"361f0f",x"301b0c",x"301c0c",x"2f1b0c",x"29170a",x"2e1a0b",x"301b0c",x"311b0c",x"2e190b",x"2d190b",x"321c0c",x"371f0e",x"361e0d",x"341d0d",x"2d180a",x"2e180b",x"311b0c",x"311b0c",x"371f0e",x"3b2210",x"3d2310",x"3a210f",x"38200e",x"381f0e",x"381f0e",x"2b180a",x"2c180b",x"301c0c",x"301b0c",x"341e0d",x"321c0d",x"361f0e",x"341d0d",x"331d0d",x"311b0c",x"321b0b",x"341d0c",x"351d0d",x"361e0e",x"26160a",x"25160a",x"47362b",x"47362b",x"452712",x"371f0d",x"361e0d",x"371e0d",x"331c0c",x"361e0d",x"38200f",x"37200e",x"361f0f",x"37200e",x"3b220f",x"341e0d",x"361f0e",x"351e0e",x"2e1a0b",x"2e1a0b",x"2c180a",x"2d1a0b",x"2c190b",x"29180a",x"311b0c",x"2b180a",x"2b170a",x"241409",x"28170a",x"28170a",x"29170a",x"29170a",x"2c190b",x"28170a",x"301b0b",x"29170a",x"2e1a0b",x"2c190b",x"321d0e",x"351f0f",x"341f0e",x"321d0d",x"311c0d",x"2f1b0c",x"2e1a0c",x"2c190b",x"2d1a0b",x"2d1a0b",x"2b180b",x"2d1a0c",x"2f1b0c",x"2d1a0b",x"2c190b",x"29170b",x"2b180b",x"29180b",x"2c190b",x"27170a",x"28170a",x"25160a",x"180f07",x"180f07",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"3d210f",x"3d210f",x"150e07",x"150e07",x"29170a",x"41342a",x"41342a",x"3e3229",x"4b2a14",x"4b2a14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"492a14",x"492a14",x"533117",x"583319",x"553218",x"533017",x"4f2d15",x"4d2c14",x"4d2b14",x"4e2c14",x"522f16",x"4b2912",x"502d15",x"532f16",x"522e15",x"482912",x"4f2d15",x"4f2b14",x"4d2c14",x"4c2a14",x"452711",x"4c2b13",x"512d15",x"553118",x"543117",x"523118",x"563318",x"533018",x"533016",x"4e2c14",x"4e2c14",x"4c2a13",x"4d2a13",x"482914",x"1f1308",x"160e07",x"251708",x"1b1108",x"1b1108",x"211508",x"181007",x"201408",x"1b1108",x"1d1208",x"281909",x"271809",x"211508",x"1a1107",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"211409",x"1c1108",x"1d1108",x"191008",x"180f08",x"180f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"27160a",x"472913",x"472913",x"313131",x"313131",x"313131",x"252525",x"313131",x"575756",x"4e4e4e",x"414141",x"282828",x"373737",x"343434",x"343434",x"343434",x"363636",x"363636",x"3a3a3a",x"3b3b3b",x"414141",x"474747",x"4c4c4c",x"595959",x"4c4c4c",x"323232",x"313131",x"333333",x"333333",x"313131",x"383838",x"3e3e3e",x"454545",x"494949",x"4c4c4c",x"565656",x"404040",x"343434",x"323232",x"323232",x"323232",x"29180b",x"24150a",x"191008",x"1c1108",x"2a180a",x"1a1008",x"1c1108",x"201309",x"201309",x"28170a",x"2a180a",x"2e190b",x"201309",x"201309",x"241509",x"231409",x"27160a",x"201308",x"211309",x"29170a",x"1f1208",x"201208",x"231309",x"29170a",x"251509",x"27160a",x"241409",x"231509",x"2f1b0c",x"25160a",x"26160a",x"29180b",x"2c190b",x"2d1a0b",x"2b190b",x"28170a",x"27170a",x"28170b",x"28170b",x"26160a",x"27160a",x"29170b",x"2e1a0c",x"2d190b",x"321d0d",x"38200f",x"39200f",x"3d2310",x"3c2210",x"3d2411",x"3d2310",x"3c220f",x"402511",x"3f2411",x"3d2310",x"3d2310",x"3c2310",x"3e2410",x"3b2210",x"3b2210",x"3c2310",x"38200e",x"3a220f",x"3b2210",x"3a2210",x"3c2311",x"331d0d",x"351e0e",x"39210f",x"38200e",x"37200e",x"39210f",x"37200f",x"361f0e",x"351e0e",x"351e0e",x"341e0e",x"36200f",x"361f0e",x"321d0e",x"301c0d",x"2c190b",x"2f1b0d",x"341e0e",x"311c0d",x"2d190b",x"331d0d",x"331e0e",x"38210f",x"37200f",x"38210f",x"351e0e",x"37200f",x"3a210f",x"39200f",x"3d2310",x"3b2210",x"3a210f",x"27170a",x"25150a",x"2c1a0b",x"2b190b",x"29170a",x"2b190b",x"2d1a0c",x"2e1a0b",x"2d190b",x"2e1a0b",x"2f1a0c",x"301b0c",x"301b0c",x"301b0c",x"2f1b0c",x"2d190b",x"2e190b",x"2d190b",x"2e1a0b",x"2b180a",x"2d190b",x"2a180a",x"2b180a",x"29170a",x"271609",x"261509",x"241409",x"271609",x"29170a",x"28160a",x"28160a",x"29170a",x"2a180a",x"2b190b",x"2b180b",x"2c1a0b",x"2c190b",x"2c190b",x"2d1a0c",x"2c1a0c",x"2b190b",x"2c190b",x"2c190b",x"2b190b",x"28170a",x"2a180b",x"2a180b",x"2a180b",x"2a180b",x"2c1a0c",x"2a180b",x"2b190b",x"2b190b",x"2a180b",x"2b190c",x"29170b",x"2a190b",x"2a190b",x"29180b",x"29180b",x"29180b",x"2a180b",x"2a180b",x"2b190b",x"2b190c",x"2a190b",x"29180b",x"2b190c",x"2a190b",x"2c1a0c",x"29180b",x"27160a",x"29180b",x"2a180b",x"28170b",x"29180b",x"29180b",x"28170b",x"28170b",x"27170b",x"26170a",x"27170b",x"27170b",x"28170b",x"28170b",x"29180b",x"27170a",x"2b190b",x"2b190b",x"28170a",x"26160a",x"2b190c",x"2d1a0c",x"2d1b0c",x"2d1a0c",x"2c1a0b",x"2c190b",x"2d1a0c",x"2e1b0c",x"2b190b",x"2f1c0d",x"2e1b0c",x"2e1b0c",x"2a180b",x"2f1b0c",x"2e1b0c",x"2d190b",x"2e1a0c",x"2d1b0c",x"2b190b",x"28170a",x"251509",x"231409",x"351e0d",x"351d0d",x"463a2f",x"463a2f",x"432510",x"391f0e",x"331c0c",x"331c0c",x"301b0b",x"27160a",x"2c180b",x"2c180a",x"2f1a0b",x"2d190a",x"29160a",x"2d170a",x"2c180a",x"311b0c",x"2e1a0b",x"2f1a0b",x"2f1a0b",x"2f1a0b",x"341d0d",x"311c0c",x"321c0d",x"311c0c",x"311c0d",x"321d0d",x"341e0d",x"2f1b0c",x"301c0d",x"301c0d",x"2f1b0c",x"27160a",x"2f1b0c",x"2e1b0c",x"2c190b",x"2f1b0c",x"321d0d",x"351e0e",x"2c1a0c",x"311c0d",x"301c0d",x"311c0d",x"2c190b",x"2f1b0c",x"2c1a0c",x"2e1b0c",x"2e1a0c",x"2b190b",x"2a180b",x"2b190b",x"2c1a0c",x"24150a",x"311c0d",x"2c190b",x"2b190c",x"2e1b0c",x"2c1a0c",x"2c1a0c",x"191008",x"191008",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"150e07",x"150e07",x"150e07",x"150e07",x"351d0d",x"513f33",x"513f33",x"534438",x"4d2c14",x"4d2c14",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"492a14",x"533117",x"583319",x"553218",x"533017",x"4f2d15",x"4d2c14",x"4d2b14",x"4e2c14",x"522f16",x"4b2912",x"502d15",x"532f16",x"522e15",x"482912",x"4f2d15",x"4f2b14",x"4d2c14",x"4c2a14",x"452711",x"4c2b13",x"512d15",x"553118",x"543117",x"523118",x"563318",x"533018",x"533016",x"4e2c14",x"4e2c14",x"4c2a13",x"3d2411",x"3d2411",x"180f07",x"160e07",x"211508",x"191107",x"191007",x"1e1308",x"170f07",x"1d1308",x"1a1107",x"1b1108",x"241708",x"231608",x"1f1408",x"191007",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e2310",x"3e2310",x"242424",x"242424",x"313131",x"303030",x"303030",x"4c4c4c",x"4a4a4a",x"414141",x"363636",x"353535",x"323232",x"313131",x"323232",x"323232",x"323232",x"313131",x"383838",x"3a3a3a",x"464646",x"505050",x"5e5e5e",x"494442",x"313131",x"313131",x"323232",x"333333",x"303030",x"383838",x"383838",x"414141",x"3d3d3d",x"4e4e4e",x"565656",x"424242",x"303030",x"333333",x"323232",x"323232",x"241509",x"1f1208",x"1e1208",x"201309",x"26160a",x"1a1008",x"231409",x"28170a",x"2c190b",x"26160a",x"1d1108",x"1d1108",x"1e1208",x"26160a",x"1e1208",x"25150a",x"28170a",x"2a180b",x"1c1108",x"1d1108",x"251509",x"26160a",x"1c1108",x"1e1108",x"231409",x"29170a",x"271609",x"1c1108",x"1c1008",x"190f07",x"1c0f07",x"251509",x"261609",x"1f1208",x"201308",x"231409",x"241509",x"201309",x"211309",x"231509",x"221409",x"221409",x"231409",x"241509",x"241409",x"251509",x"29170a",x"2b180b",x"2d1a0b",x"2f1b0c",x"2e1a0b",x"2f1b0c",x"2f1b0c",x"2f1b0c",x"2e1b0c",x"2c190b",x"2b180b",x"2a180b",x"28170a",x"29170a",x"26160a",x"26160a",x"24150a",x"25150a",x"25160a",x"26160a",x"27170a",x"26160a",x"25160a",x"24160a",x"24150a",x"25150a",x"26160a",x"201309",x"1f1309",x"1d1108",x"1b1108",x"191008",x"180f08",x"2c190b",x"2e1a0b",x"321c0d",x"301b0c",x"301b0c",x"351e0e",x"331d0d",x"311c0d",x"341d0d",x"2a180b",x"351e0e",x"37200f",x"36200e",x"351e0d",x"39200e",x"39200e",x"39210f",x"3a210f",x"371f0f",x"341e0e",x"28180a",x"2a190b",x"28180a",x"241509",x"231409",x"241509",x"28170a",x"2b190b",x"2a180a",x"28160a",x"2b180b",x"2d1a0b",x"2c190b",x"2b190b",x"2a180a",x"2b190b",x"2c190b",x"2c190b",x"2c190b",x"2c190b",x"2b180b",x"28170a",x"27160a",x"29170a",x"26160a",x"251509",x"231409",x"241509",x"241509",x"241409",x"221309",x"201208",x"1c1007",x"1a0f07",x"1f1108",x"241409",x"241509",x"251509",x"26160a",x"26160a",x"251509",x"251509",x"26150a",x"26160a",x"251509",x"251509",x"241509",x"241409",x"221409",x"231409",x"251509",x"27160a",x"26160a",x"26160a",x"26160a",x"27170a",x"26160a",x"27160a",x"26160a",x"26160a",x"26160a",x"27160a",x"26160a",x"26160a",x"27170a",x"25150a",x"26160a",x"26160a",x"27170b",x"28170b",x"27170a",x"28170b",x"27170a",x"26160a",x"25160a",x"25160a",x"24150a",x"211409",x"201309",x"1f1209",x"1f1209",x"1e1208",x"1f1209",x"1f1309",x"201309",x"211309",x"211409",x"211409",x"221409",x"221409",x"231409",x"23150a",x"24150a",x"25160a",x"26160a",x"24150a",x"241509",x"26160a",x"25150a",x"27170a",x"26160a",x"28180b",x"28180b",x"28180b",x"29180b",x"27160a",x"241509",x"231409",x"241509",x"24150a",x"221409",x"1e1208",x"2f1b0b",x"331d0d",x"311b0b",x"311b0b",x"4b2a12",x"442511",x"442611",x"472812",x"412510",x"3e2310",x"402410",x"3d220f",x"371e0d",x"3d220f",x"40230f",x"3a200d",x"381e0d",x"361d0c",x"361e0c",x"331c0c",x"361d0c",x"331b0b",x"2e180a",x"211006",x"231106",x"361d0c",x"351d0c",x"371e0d",x"3b200f",x"3c210f",x"361f0d",x"351d0d",x"39200e",x"3d2210",x"361e0d",x"331c0d",x"311b0c",x"321b0b",x"321b0b",x"321b0b",x"361e0d",x"371f0e",x"341d0d",x"38200e",x"39200e",x"39200f",x"3a210f",x"3a210f",x"38200e",x"371f0e",x"371f0e",x"3a210f",x"331d0d",x"39200f",x"37200e",x"38200f",x"351e0d",x"331d0d",x"351e0e",x"331d0e",x"211409",x"211409",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1108",x"1d1108",x"442610",x"40240f",x"402310",x"351e0f",x"351e0f",x"4e301c",x"513520",x"513520",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"38200f",x"38200f",x"170f07",x"150e07",x"1d1308",x"181007",x"180f07",x"1b1108",x"160f07",x"1b1108",x"181007",x"191007",x"201408",x"1f1408",x"1c1208",x"170f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"3e220f",x"3e220f",x"313131",x"313131",x"343434",x"303030",x"333333",x"323232",x"333333",x"373737",x"404040",x"343434",x"313131",x"313131",x"323232",x"333333",x"323232",x"343434",x"333333",x"393939",x"474747",x"515151",x"5c5c5c",x"4d4d4d",x"333333",x"333333",x"303030",x"333333",x"313131",x"333333",x"313131",x"3a3a3a",x"464646",x"565656",x"5d5d5d",x"404040",x"333333",x"313131",x"2a2a2a",x"2a2a2a",x"1d1208",x"38200f",x"3e2310",x"412611",x"412511",x"3e220f",x"402310",x"432511",x"3f220f",x"432510",x"422511",x"3e230f",x"452711",x"452812",x"432611",x"432511",x"422410",x"3c210e",x"40220f",x"3e220e",x"3d210f",x"3d220f",x"3d220e",x"371c0c",x"3c210e",x"452611",x"412410",x"381f0d",x"3f230f",x"3f230f",x"3e230f",x"3f230f",x"3f230f",x"3a200e",x"3c210e",x"3d220f",x"3d220f",x"3b200e",x"3a200f",x"472a15",x"432813",x"432713",x"442813",x"402612",x"3f2411",x"3a200e",x"381f0d",x"371e0d",x"3a200e",x"3a200e",x"402410",x"452813",x"422612",x"412511",x"442813",x"3f2410",x"3e220f",x"3e220f",x"371d0d",x"371e0d",x"3a200e",x"3d2310",x"3e2411",x"402511",x"402511",x"412512",x"381f0e",x"371f0e",x"3b210f",x"3c220f",x"3e2410",x"3e2310",x"402511",x"3f2410",x"3d2310",x"3c2210",x"3f2411",x"3d2310",x"3b2210",x"3c220f",x"452812",x"3f2411",x"3f2411",x"3e2411",x"432712",x"3d2310",x"3f2411",x"412511",x"3d220f",x"3d210e",x"3e220f",x"3f2310",x"3f2410",x"432511",x"432611",x"422511",x"442611",x"462813",x"442812",x"442712",x"2d1b0b",x"361f0e",x"351f0e",x"331d0d",x"341d0d",x"37200e",x"3a210f",x"361e0d",x"391f0e",x"361e0d",x"371e0d",x"391f0e",x"3b210e",x"3b210e",x"3b210f",x"39210f",x"38200e",x"331c0c",x"341c0d",x"321c0c",x"321c0c",x"321b0c",x"321c0c",x"351e0d",x"311b0c",x"2e190a",x"2d180a",x"361e0d",x"331c0c",x"351d0d",x"331c0c",x"351e0d",x"351e0d",x"361e0d",x"351e0d",x"361e0d",x"361e0d",x"381f0e",x"381f0e",x"381f0e",x"3a200e",x"3d220f",x"3f2612",x"3c2411",x"422712",x"3e2411",x"3e2411",x"3a200e",x"331c0c",x"361d0d",x"341d0d",x"381e0d",x"3b210f",x"3e2411",x"3f2511",x"38200f",x"3c2310",x"3b220f",x"381f0e",x"351d0d",x"351d0c",x"341c0c",x"341d0c",x"39200f",x"39210f",x"37200e",x"37200e",x"3b220f",x"351e0d",x"351d0d",x"371f0e",x"38200e",x"39210f",x"38200e",x"371f0e",x"361f0e",x"3b220f",x"341e0e",x"361f0e",x"38200f",x"341e0e",x"37200e",x"2d1a0c",x"2b190b",x"29180b",x"2c190b",x"29180b",x"29180b",x"2e1b0c",x"2e1a0c",x"2b190b",x"2b190b",x"2a170a",x"29170a",x"221409",x"231509",x"29170a",x"321c0c",x"3a200e",x"3c2210",x"3b220f",x"3c2310",x"3d2310",x"3c2310",x"3e2411",x"3b220f",x"39200f",x"3e2410",x"412511",x"3a200e",x"3c210e",x"402310",x"432611",x"432611",x"432610",x"4a2913",x"3f230f",x"381f0e",x"3b210e",x"381f0e",x"331c0c",x"2e1a0b",x"341d0c",x"311b0c",x"39200f",x"341d0d",x"331d0d",x"321c0c",x"301b0c",x"361e0d",x"2e1a0b",x"2e190b",x"351d0d",x"301b0b",x"311b0c",x"341d0c",x"261308",x"241308",x"321c0c",x"38200e",x"311b0a",x"371e0c",x"371e0d",x"331b0c",x"361d0d",x"2d190b",x"361e0d",x"38200f",x"38200f",x"311b0c",x"301c0c",x"351e0d",x"331c0c",x"331c0d",x"311b0c",x"331c0c",x"311b0b",x"231409",x"2d190b",x"351d0d",x"321c0c",x"2c190b",x"311b0c",x"321c0d",x"2f1b0b",x"311c0c",x"2d190b",x"301a0b",x"301b0b",x"311b0b",x"3d220f",x"331d0e",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"1d1108",x"442610",x"40240f",x"402310",x"000000",x"351e0f",x"4e301c",x"513520",x"513520",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000"),
(x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"311c0c",x"311c0c",x"160e07",x"150e07",x"191007",x"160f07",x"160f07",x"180f07",x"160e07",x"170f07",x"160f07",x"170f07",x"1a1107",x"191007",x"180f07",x"160f07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"150e07",x"442711",x"442711",x"323232",x"323232",x"303030",x"2e2e2e",x"323232",x"323232",x"333333",x"373737",x"363636",x"343434",x"2d2d2d",x"333333",x"313131",x"5b5957",x"605d5a",x"6a6765",x"656361",x"646362",x"565554",x"515150",x"4f4e4e",x"676767",x"313131",x"333333",x"2c2c2c",x"323232",x"44413d",x"63605d",x"656360",x"595857",x"51504f",x"555554",x"51504f",x"616161",x"323232",x"313131",x"303030",x"303030",x"150e07",x"2d1c0f",x"412513",x"3f2512",x"442713",x"452712",x"442712",x"452712",x"442611",x"432510",x"41240f",x"41240f",x"452711",x"472912",x"492a13",x"482913",x"4b2b14",x"432611",x"462711",x"442510",x"422410",x"3e220e",x"422410",x"40220f",x"3d200d",x"452611",x"4a2a14",x"462711",x"462811",x"432611",x"41240f",x"3c210e",x"3c210e",x"3e220f",x"412410",x"452611",x"452711",x"452711",x"462812",x"4a2a14",x"492b14",x"4a2c14",x"482914",x"462812",x"422511",x"452812",x"452812",x"412511",x"432511",x"412410",x"40230f",x"402310",x"442611",x"432712",x"452712",x"452712",x"442611",x"432611",x"422510",x"432611",x"442712",x"412511",x"412410",x"412510",x"452712",x"462812",x"432611",x"412410",x"422410",x"402410",x"3f210e",x"3f230f",x"3f220f",x"3d210e",x"3b200e",x"402310",x"442611",x"452712",x"442611",x"452712",x"482912",x"472812",x"462812",x"422511",x"402410",x"3f230f",x"3f230f",x"402410",x"402310",x"3c220e",x"3a200e",x"351d0c",x"321c0c",x"381f0e",x"39200e",x"3e230f",x"3b210f",x"3b210f",x"3d2310",x"412511",x"29190a",x"311c0c",x"331d0d",x"361f0e",x"39200e",x"3c220e",x"3e240f",x"412510",x"432711",x"432711",x"432711",x"452711",x"442711",x"402510",x"40240f",x"432611",x"3f2510",x"3f2410",x"3b220f",x"3d2310",x"381f0e",x"371e0d",x"341d0c",x"361d0d",x"371e0d",x"381f0e",x"351e0d",x"351d0d",x"361e0d",x"3a200f",x"3a210e",x"3b210e",x"381f0d",x"371e0d",x"38200e",x"3a210f",x"3b210f",x"3e2310",x"402411",x"3a200e",x"3c220f",x"3f2410",x"422612",x"3d2310",x"39200e",x"381e0e",x"381e0d",x"3f2410",x"432612",x"3e230f",x"3e220f",x"3d220f",x"3f230f",x"3d210e",x"3f230f",x"412511",x"3f2310",x"432611",x"432611",x"442712",x"432611",x"432611",x"442612",x"432712",x"432612",x"422611",x"412511",x"422611",x"412511",x"3d220f",x"3e220f",x"3c210f",x"402410",x"3f230f",x"3f2310",x"432511",x"3f2410",x"402410",x"3f2410",x"3e230f",x"3f2310",x"432612",x"402410",x"3f2310",x"3e2310",x"412511",x"3f2410",x"402510",x"402410",x"3c220f",x"3e220f",x"371e0d",x"351d0d",x"371e0d",x"321b0b",x"331c0b",x"381e0d",x"3e220f",x"412511",x"432611",x"442712",x"462913",x"432611",x"432610",x"412510",x"412510",x"40240f",x"432711",x"472812",x"442710",x"4d2d13",x"4e2e13",x"4e2e13",x"000000",x"000000",x"4a2913",x"3f230f",x"381f0e",x"3b210e",x"381f0e",x"331c0c",x"2e1a0b",x"341d0c",x"311b0c",x"39200f",x"341d0d",x"331d0d",x"321c0c",x"301b0c",x"361e0d",x"2e1a0b",x"2e190b",x"351d0d",x"301b0b",x"311b0c",x"341d0c",x"261308",x"241308",x"321c0c",x"38200e",x"311b0a",x"371e0c",x"371e0d",x"331b0c",x"361d0d",x"2d190b",x"361e0d",x"38200f",x"38200f",x"311b0c",x"301c0c",x"351e0d",x"331c0c",x"331c0d",x"311b0c",x"331c0c",x"311b0b",x"231409",x"2d190b",x"351d0d",x"321c0c",x"2c190b",x"311b0c",x"321c0d",x"2f1b0b",x"311c0c",x"2d190b",x"301a0b",x"301b0b",x"311b0b",x"3d220f",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000",x"000000")
);

end texture;

package body texture is


end texture;
